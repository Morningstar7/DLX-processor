library IEEE;
use IEEE.std_logic_1164.all;

entity FETCH is 
	generic (	N:		integer);
	port (		JUMP_ADDR:	in 	std_logic_vector(N-1 downto 0);		--ADDRESS FOR BRANCHING AND JUMPING
			BPU_ADDR:	in	std_logic_vector(N-1 downto 0);
			NPC_IN:		in	std_logic_vector(N-1 downto 0);
			BRANCH_SEL:	in	std_logic;
			BRANCH_SEL_BPU:	in	std_logic;
			SEL_N_TAKEN:	in	std_logic;
			EN:		in	std_logic;
			RST:		in	std_logic;
			CLK:		in	std_logic;
			DATA_IN_INSTR:	in	std_logic_vector(7 downto 0);
			H_M_CACHE:	out	std_logic;
			ADDR_IRAM:	out	std_logic_vector(N-1 downto 0);
			PC_OUT:		out	std_logic_vector(N-1 downto 0);
			NPC: 		out	std_logic_vector(N-1 downto 0);		--NEW PROGRAM COUNTER
			INSTRUCTION:	out	std_logic_vector(n-1 downto 0));	--INSTRUCTION OUT
end FETCH;

architecture STRUCTURAL of FETCH is

	component REG
		generic (	N:	integer);
		port (		D: 	in 	std_logic_vector(N-1 downto 0);
				Q: 	out	std_logic_vector(N-1 downto 0);
				EN:	in	std_logic;
				RST:	in 	std_logic;
				CLK: 	in	std_logic);
	end component;
	
	component CACHE
		generic (	N:		integer;
				TAG_BIT:	integer;
				SET_BIT:	integer;
				N_DATA:		integer);
		port (		ADDR:		in	std_logic_vector(N-1 downto 0);
				ADDR_OUT:	out	std_logic_vector(N-1 downto 0);
				DATA_IN:	in	std_logic_vector(7 downto 0);
				DATA_OUT:	out	std_logic_vector(N-1 downto 0);
				RST:		in	std_logic;
				LOAD:		in	std_logic;
				CLK:		in	std_logic;
				HIT_MISS:	out	std_logic);
	end component;
	
	component RCA_GEN_NO_C
		generic (	N:	integer);
		Port (		A:	in	std_logic_vector(N-1 downto 0);
				B:	in	std_logic_vector(N-1 downto 0);
				S:	out	std_logic_vector(N-1 downto 0);
				Co:	out	std_logic);
	end component;
	
	component MUX21_GEN
		generic (	N: 	integer);
		port (		A:	in	std_logic_vector(N-1 downto 0);
				B:	in	std_logic_vector(N-1 downto 0);
				SEL:	in	std_logic;
				Y:	out	std_logic_vector(N-1 downto 0));
	end component;
	
	--PC SIGNALS:
	--####################
	signal OUT_PC:	std_logic_vector(N-1 downto 0);
	--####################
	
	--CACHE SIGNALS:
	--####################
	signal OUT_CACHE:	std_logic_vector(N-1 downto 0);
	signal CACHE_LOAD:	std_logic;
	signal HIT_MISS:	std_logic;
	--####################
	
	--ADDER SIGNALS:
	--####################
	signal A_ADDER:		std_logic_vector(N-3 downto 0);
	signal B_ADDER:		std_logic_vector(N-3 downto 0);
	signal OUT_ADDER:	std_logic_vector(N-3 downto 0);
	signal Co_ADDER:	std_logic;
	--####################
	
	--MUX SIGNALS:
	--####################
	signal B_MUX:	std_logic_vector(N-1 downto 0);
	signal OUT_MUX:	std_logic_vector(N-1 downto 0);
	signal OUT_MUX_1:	std_logic_vector(N-1 downto 0);
	signal OUT_MUX_2:	std_logic_vector(N-1 downto 0);
	--####################
	
	begin
	
		PC: REG	generic map (	N => N)
			port map (	D => OUT_MUX_2,
					Q => OUT_PC,
					EN => EN,
					RST => RST,
					CLK => CLK);
		
		INSTRUCTION_CACHE: CACHE	generic map (	N => N,
								TAG_BIT => 23,
								SET_BIT => 4,
								N_DATA => 5)
						port map (	ADDR => OUT_PC,
								ADDR_OUT => ADDR_IRAM,
								DATA_IN => DATA_IN_INSTR,
								DATA_OUT => OUT_CACHE,
								RST => RST,
								LOAD => CACHE_LOAD,
								CLK => CLK,
								HIT_MISS => HIT_MISS);
		
		--CACHE SIGNAL ASSOCIATION:
		--####################
		CACHE_LOAD <= not HIT_MISS and not RST;
		H_M_CACHE <= HIT_MISS;
		--####################
		
		PC_ADDER: RCA_GEN_NO_C	generic map (	N => N-2)
					port map (	A => A_ADDER,
							B => B_ADDER,
							S => OUT_ADDER,
							Co => Co_ADDER);
		
		--ADDER SIGNAL ASSOCIATION:
		--####################
		A_ADDER <= OUT_PC(N-1 downto 2);
		B_ADDER <= (0 => '1', others => '0');
		--####################
		
		MUX_PC: MUX21_GEN	generic map (	N => N)
					port map (	A => JUMP_ADDR,
							B => B_MUX,
							SEL => BRANCH_SEL,
							Y => OUT_MUX);

		MUX_BPU: MUX21_GEN	generic map (	N => N)
					port map (	A => BPU_ADDR,
							B => OUT_MUX,
							SEL => BRANCH_SEL_BPU,
							Y => OUT_MUX_1);

		MUX_N_TAKEN: MUX21_GEN	generic map (	N => N)
					port map (	A => NPC_IN,
							B => OUT_MUX_1,
							SEL => SEL_N_TAKEN,
							Y => OUT_MUX_2);
		
		--MUX SIGNAL ASSOCIATION:
		--####################
		B_MUX <= OUT_ADDER & OUT_PC(1 downto 0);
		--####################
		
		--FETCH SIGNAL ASSOCIATION:
		--####################
		NPC <= OUT_ADDER & OUT_PC(1 downto 0);
		INSTRUCTION <= OUT_CACHE;
		PC_OUT <= OUT_PC;
		--####################

end STRUCTURAL;

configuration CFG_FETCH_STRUCTURAL of FETCH is
	for STRUCTURAL
		for all: REG
			use configuration WORK.CFG_REG_SYN_STRUCTURAL;
		end for;
		for all: CACHE
			use configuration WORK.CFG_CACHE_STRUCTURAL;
		end for;
		for all: RCA_GEN_NO_C
			use configuration WORK.CFG_RCA_GEN_NO_C_STRUCTURAL;
		end for;
		for all: MUX21_GEN
			use configuration WORK.CFG_MUX21_GEN_STRUCTURAL;
		end for;
	end for;
end CFG_FETCH_STRUCTURAL;