
module FSM_DIVISOR_DW01_inc_0 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   \carry[31] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ,
         \carry[11] , \carry[10] , \carry[9] , \carry[8] , \carry[7] ,
         \carry[6] , \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA_X1 U1_1_30 ( .A(A[30]), .B(\carry[30] ), .CO(\carry[31] ), .S(SUM[30]) );
  HA_X1 U1_1_29 ( .A(A[29]), .B(\carry[29] ), .CO(\carry[30] ), .S(SUM[29]) );
  HA_X1 U1_1_28 ( .A(A[28]), .B(\carry[28] ), .CO(\carry[29] ), .S(SUM[28]) );
  HA_X1 U1_1_27 ( .A(A[27]), .B(\carry[27] ), .CO(\carry[28] ), .S(SUM[27]) );
  HA_X1 U1_1_26 ( .A(A[26]), .B(\carry[26] ), .CO(\carry[27] ), .S(SUM[26]) );
  HA_X1 U1_1_25 ( .A(A[25]), .B(\carry[25] ), .CO(\carry[26] ), .S(SUM[25]) );
  HA_X1 U1_1_24 ( .A(A[24]), .B(\carry[24] ), .CO(\carry[25] ), .S(SUM[24]) );
  HA_X1 U1_1_23 ( .A(A[23]), .B(\carry[23] ), .CO(\carry[24] ), .S(SUM[23]) );
  HA_X1 U1_1_22 ( .A(A[22]), .B(\carry[22] ), .CO(\carry[23] ), .S(SUM[22]) );
  HA_X1 U1_1_21 ( .A(A[21]), .B(\carry[21] ), .CO(\carry[22] ), .S(SUM[21]) );
  HA_X1 U1_1_20 ( .A(A[20]), .B(\carry[20] ), .CO(\carry[21] ), .S(SUM[20]) );
  HA_X1 U1_1_19 ( .A(A[19]), .B(\carry[19] ), .CO(\carry[20] ), .S(SUM[19]) );
  HA_X1 U1_1_18 ( .A(A[18]), .B(\carry[18] ), .CO(\carry[19] ), .S(SUM[18]) );
  HA_X1 U1_1_17 ( .A(A[17]), .B(\carry[17] ), .CO(\carry[18] ), .S(SUM[17]) );
  HA_X1 U1_1_16 ( .A(A[16]), .B(\carry[16] ), .CO(\carry[17] ), .S(SUM[16]) );
  HA_X1 U1_1_15 ( .A(A[15]), .B(\carry[15] ), .CO(\carry[16] ), .S(SUM[15]) );
  HA_X1 U1_1_14 ( .A(A[14]), .B(\carry[14] ), .CO(\carry[15] ), .S(SUM[14]) );
  HA_X1 U1_1_13 ( .A(A[13]), .B(\carry[13] ), .CO(\carry[14] ), .S(SUM[13]) );
  HA_X1 U1_1_12 ( .A(A[12]), .B(\carry[12] ), .CO(\carry[13] ), .S(SUM[12]) );
  HA_X1 U1_1_11 ( .A(A[11]), .B(\carry[11] ), .CO(\carry[12] ), .S(SUM[11]) );
  HA_X1 U1_1_10 ( .A(A[10]), .B(\carry[10] ), .CO(\carry[11] ), .S(SUM[10]) );
  HA_X1 U1_1_9 ( .A(A[9]), .B(\carry[9] ), .CO(\carry[10] ), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(\carry[8] ), .CO(\carry[9] ), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(\carry[7] ), .CO(\carry[8] ), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(\carry[6] ), .CO(\carry[7] ), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(\carry[5] ), .CO(\carry[6] ), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(\carry[31] ), .B(A[31]), .Z(SUM[31]) );
  INV_X1 U2 ( .A(A[0]), .ZN(SUM[0]) );
endmodule


module FORW_FSM_OPCODE_SIZE6_N_ADDR5_DW01_inc_1 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   \carry[31] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ,
         \carry[11] , \carry[10] , \carry[9] , \carry[8] , \carry[7] ,
         \carry[6] , \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA_X1 U1_1_30 ( .A(A[30]), .B(\carry[30] ), .CO(\carry[31] ), .S(SUM[30]) );
  HA_X1 U1_1_29 ( .A(A[29]), .B(\carry[29] ), .CO(\carry[30] ), .S(SUM[29]) );
  HA_X1 U1_1_28 ( .A(A[28]), .B(\carry[28] ), .CO(\carry[29] ), .S(SUM[28]) );
  HA_X1 U1_1_27 ( .A(A[27]), .B(\carry[27] ), .CO(\carry[28] ), .S(SUM[27]) );
  HA_X1 U1_1_26 ( .A(A[26]), .B(\carry[26] ), .CO(\carry[27] ), .S(SUM[26]) );
  HA_X1 U1_1_25 ( .A(A[25]), .B(\carry[25] ), .CO(\carry[26] ), .S(SUM[25]) );
  HA_X1 U1_1_24 ( .A(A[24]), .B(\carry[24] ), .CO(\carry[25] ), .S(SUM[24]) );
  HA_X1 U1_1_23 ( .A(A[23]), .B(\carry[23] ), .CO(\carry[24] ), .S(SUM[23]) );
  HA_X1 U1_1_22 ( .A(A[22]), .B(\carry[22] ), .CO(\carry[23] ), .S(SUM[22]) );
  HA_X1 U1_1_21 ( .A(A[21]), .B(\carry[21] ), .CO(\carry[22] ), .S(SUM[21]) );
  HA_X1 U1_1_20 ( .A(A[20]), .B(\carry[20] ), .CO(\carry[21] ), .S(SUM[20]) );
  HA_X1 U1_1_19 ( .A(A[19]), .B(\carry[19] ), .CO(\carry[20] ), .S(SUM[19]) );
  HA_X1 U1_1_18 ( .A(A[18]), .B(\carry[18] ), .CO(\carry[19] ), .S(SUM[18]) );
  HA_X1 U1_1_17 ( .A(A[17]), .B(\carry[17] ), .CO(\carry[18] ), .S(SUM[17]) );
  HA_X1 U1_1_16 ( .A(A[16]), .B(\carry[16] ), .CO(\carry[17] ), .S(SUM[16]) );
  HA_X1 U1_1_15 ( .A(A[15]), .B(\carry[15] ), .CO(\carry[16] ), .S(SUM[15]) );
  HA_X1 U1_1_14 ( .A(A[14]), .B(\carry[14] ), .CO(\carry[15] ), .S(SUM[14]) );
  HA_X1 U1_1_13 ( .A(A[13]), .B(\carry[13] ), .CO(\carry[14] ), .S(SUM[13]) );
  HA_X1 U1_1_12 ( .A(A[12]), .B(\carry[12] ), .CO(\carry[13] ), .S(SUM[12]) );
  HA_X1 U1_1_11 ( .A(A[11]), .B(\carry[11] ), .CO(\carry[12] ), .S(SUM[11]) );
  HA_X1 U1_1_10 ( .A(A[10]), .B(\carry[10] ), .CO(\carry[11] ), .S(SUM[10]) );
  HA_X1 U1_1_9 ( .A(A[9]), .B(\carry[9] ), .CO(\carry[10] ), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(\carry[8] ), .CO(\carry[9] ), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(\carry[7] ), .CO(\carry[8] ), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(\carry[6] ), .CO(\carry[7] ), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(\carry[5] ), .CO(\carry[6] ), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(\carry[31] ), .B(A[31]), .Z(SUM[31]) );
  INV_X1 U2 ( .A(A[0]), .ZN(SUM[0]) );
endmodule


module FORW_FSM_OPCODE_SIZE6_N_ADDR5_DW01_inc_0 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   \carry[31] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ,
         \carry[11] , \carry[10] , \carry[9] , \carry[8] , \carry[7] ,
         \carry[6] , \carry[5] , \carry[4] , \carry[3] , \carry[2] ;

  HA_X1 U1_1_30 ( .A(A[30]), .B(\carry[30] ), .CO(\carry[31] ), .S(SUM[30]) );
  HA_X1 U1_1_29 ( .A(A[29]), .B(\carry[29] ), .CO(\carry[30] ), .S(SUM[29]) );
  HA_X1 U1_1_28 ( .A(A[28]), .B(\carry[28] ), .CO(\carry[29] ), .S(SUM[28]) );
  HA_X1 U1_1_27 ( .A(A[27]), .B(\carry[27] ), .CO(\carry[28] ), .S(SUM[27]) );
  HA_X1 U1_1_26 ( .A(A[26]), .B(\carry[26] ), .CO(\carry[27] ), .S(SUM[26]) );
  HA_X1 U1_1_25 ( .A(A[25]), .B(\carry[25] ), .CO(\carry[26] ), .S(SUM[25]) );
  HA_X1 U1_1_24 ( .A(A[24]), .B(\carry[24] ), .CO(\carry[25] ), .S(SUM[24]) );
  HA_X1 U1_1_23 ( .A(A[23]), .B(\carry[23] ), .CO(\carry[24] ), .S(SUM[23]) );
  HA_X1 U1_1_22 ( .A(A[22]), .B(\carry[22] ), .CO(\carry[23] ), .S(SUM[22]) );
  HA_X1 U1_1_21 ( .A(A[21]), .B(\carry[21] ), .CO(\carry[22] ), .S(SUM[21]) );
  HA_X1 U1_1_20 ( .A(A[20]), .B(\carry[20] ), .CO(\carry[21] ), .S(SUM[20]) );
  HA_X1 U1_1_19 ( .A(A[19]), .B(\carry[19] ), .CO(\carry[20] ), .S(SUM[19]) );
  HA_X1 U1_1_18 ( .A(A[18]), .B(\carry[18] ), .CO(\carry[19] ), .S(SUM[18]) );
  HA_X1 U1_1_17 ( .A(A[17]), .B(\carry[17] ), .CO(\carry[18] ), .S(SUM[17]) );
  HA_X1 U1_1_16 ( .A(A[16]), .B(\carry[16] ), .CO(\carry[17] ), .S(SUM[16]) );
  HA_X1 U1_1_15 ( .A(A[15]), .B(\carry[15] ), .CO(\carry[16] ), .S(SUM[15]) );
  HA_X1 U1_1_14 ( .A(A[14]), .B(\carry[14] ), .CO(\carry[15] ), .S(SUM[14]) );
  HA_X1 U1_1_13 ( .A(A[13]), .B(\carry[13] ), .CO(\carry[14] ), .S(SUM[13]) );
  HA_X1 U1_1_12 ( .A(A[12]), .B(\carry[12] ), .CO(\carry[13] ), .S(SUM[12]) );
  HA_X1 U1_1_11 ( .A(A[11]), .B(\carry[11] ), .CO(\carry[12] ), .S(SUM[11]) );
  HA_X1 U1_1_10 ( .A(A[10]), .B(\carry[10] ), .CO(\carry[11] ), .S(SUM[10]) );
  HA_X1 U1_1_9 ( .A(A[9]), .B(\carry[9] ), .CO(\carry[10] ), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(\carry[8] ), .CO(\carry[9] ), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(\carry[7] ), .CO(\carry[8] ), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(\carry[6] ), .CO(\carry[7] ), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(\carry[5] ), .CO(\carry[6] ), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(\carry[31] ), .B(A[31]), .Z(SUM[31]) );
  INV_X1 U2 ( .A(A[0]), .ZN(SUM[0]) );
endmodule


module GENERAL_PROPAGATE_26 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_438 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_25 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_436 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_24 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_434 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_23 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_432 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_22 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_430 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_21 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_428 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_20 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_426 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_19 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_424 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_18 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_422 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_17 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_420 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_16 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_418 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_15 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_416 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_14 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_414 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_13 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_412 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_12 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_410 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_11 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_408 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_10 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_406 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_9 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_404 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_8 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_402 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_7 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_400 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_6 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_398 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_5 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_396 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_4 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_394 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_3 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_392 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_2 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_390 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module GENERAL_PROPAGATE_1 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_388 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module MUX41_GEN_N16_1 ( A, B, C, D, SEL, Y );
  input [15:0] A;
  input [15:0] B;
  input [15:0] C;
  input [15:0] D;
  input [1:0] SEL;
  output [15:0] Y;
  wire   n1, n2, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74;

  NAND2_X1 U38 ( .A1(n74), .A2(n73), .ZN(Y[9]) );
  NAND2_X1 U39 ( .A1(n68), .A2(n67), .ZN(Y[8]) );
  NAND2_X1 U40 ( .A1(n66), .A2(n65), .ZN(Y[7]) );
  NAND2_X1 U41 ( .A1(n64), .A2(n63), .ZN(Y[6]) );
  NAND2_X1 U42 ( .A1(n62), .A2(n61), .ZN(Y[5]) );
  NAND2_X1 U43 ( .A1(n60), .A2(n59), .ZN(Y[4]) );
  NAND2_X1 U44 ( .A1(n58), .A2(n57), .ZN(Y[3]) );
  NAND2_X1 U45 ( .A1(n56), .A2(n55), .ZN(Y[2]) );
  NAND2_X1 U46 ( .A1(n54), .A2(n53), .ZN(Y[1]) );
  NAND2_X1 U47 ( .A1(n52), .A2(n51), .ZN(Y[15]) );
  NAND2_X1 U48 ( .A1(n50), .A2(n49), .ZN(Y[14]) );
  NAND2_X1 U49 ( .A1(n48), .A2(n47), .ZN(Y[13]) );
  NAND2_X1 U50 ( .A1(n46), .A2(n45), .ZN(Y[12]) );
  NAND2_X1 U51 ( .A1(n44), .A2(n43), .ZN(Y[11]) );
  NAND2_X1 U52 ( .A1(n42), .A2(n41), .ZN(Y[10]) );
  NAND2_X1 U53 ( .A1(n40), .A2(n39), .ZN(Y[0]) );
  BUF_X1 U1 ( .A(n71), .Z(n1) );
  NOR3_X4 U2 ( .A1(n1), .A2(n69), .A3(n72), .ZN(n70) );
  INV_X1 U3 ( .A(SEL[0]), .ZN(n2) );
  AND2_X1 U4 ( .A1(SEL[1]), .A2(n2), .ZN(n72) );
  AND2_X1 U5 ( .A1(SEL[0]), .A2(SEL[1]), .ZN(n69) );
  NOR2_X1 U6 ( .A1(n2), .A2(SEL[1]), .ZN(n71) );
  AOI22_X1 U7 ( .A1(B[3]), .A2(n72), .B1(C[3]), .B2(n1), .ZN(n57) );
  AOI22_X1 U8 ( .A1(B[0]), .A2(n72), .B1(C[0]), .B2(n1), .ZN(n39) );
  AOI22_X1 U9 ( .A1(B[1]), .A2(n72), .B1(C[1]), .B2(n1), .ZN(n53) );
  AOI22_X1 U10 ( .A1(B[2]), .A2(n72), .B1(C[2]), .B2(n1), .ZN(n55) );
  AOI22_X1 U11 ( .A1(B[4]), .A2(n72), .B1(C[4]), .B2(n1), .ZN(n59) );
  AOI22_X1 U12 ( .A1(B[5]), .A2(n72), .B1(C[5]), .B2(n1), .ZN(n61) );
  AOI22_X1 U13 ( .A1(B[6]), .A2(n72), .B1(C[6]), .B2(n1), .ZN(n63) );
  AOI22_X1 U14 ( .A1(B[7]), .A2(n72), .B1(C[7]), .B2(n1), .ZN(n65) );
  AOI22_X1 U15 ( .A1(B[8]), .A2(n72), .B1(C[8]), .B2(n1), .ZN(n67) );
  AOI22_X1 U16 ( .A1(B[9]), .A2(n72), .B1(C[9]), .B2(n1), .ZN(n73) );
  AOI22_X1 U17 ( .A1(B[10]), .A2(n72), .B1(C[10]), .B2(n1), .ZN(n41) );
  AOI22_X1 U18 ( .A1(B[11]), .A2(n72), .B1(C[11]), .B2(n1), .ZN(n43) );
  AOI22_X1 U19 ( .A1(B[12]), .A2(n72), .B1(C[12]), .B2(n1), .ZN(n45) );
  AOI22_X1 U20 ( .A1(B[13]), .A2(n72), .B1(C[13]), .B2(n1), .ZN(n47) );
  AOI22_X1 U21 ( .A1(B[14]), .A2(n72), .B1(C[14]), .B2(n1), .ZN(n49) );
  AOI22_X1 U22 ( .A1(B[15]), .A2(n72), .B1(C[15]), .B2(n1), .ZN(n51) );
  AOI22_X1 U23 ( .A1(D[14]), .A2(n70), .B1(A[14]), .B2(n69), .ZN(n50) );
  AOI22_X1 U24 ( .A1(D[15]), .A2(n70), .B1(A[15]), .B2(n69), .ZN(n52) );
  AOI22_X1 U25 ( .A1(D[12]), .A2(n70), .B1(A[12]), .B2(n69), .ZN(n46) );
  AOI22_X1 U26 ( .A1(D[10]), .A2(n70), .B1(A[10]), .B2(n69), .ZN(n42) );
  AOI22_X1 U27 ( .A1(D[8]), .A2(n70), .B1(A[8]), .B2(n69), .ZN(n68) );
  AOI22_X1 U28 ( .A1(D[6]), .A2(n70), .B1(A[6]), .B2(n69), .ZN(n64) );
  AOI22_X1 U29 ( .A1(D[13]), .A2(n70), .B1(A[13]), .B2(n69), .ZN(n48) );
  AOI22_X1 U30 ( .A1(D[4]), .A2(n70), .B1(A[4]), .B2(n69), .ZN(n60) );
  AOI22_X1 U31 ( .A1(D[11]), .A2(n70), .B1(A[11]), .B2(n69), .ZN(n44) );
  AOI22_X1 U32 ( .A1(D[7]), .A2(n70), .B1(A[7]), .B2(n69), .ZN(n66) );
  AOI22_X1 U33 ( .A1(D[9]), .A2(n70), .B1(A[9]), .B2(n69), .ZN(n74) );
  AOI22_X1 U34 ( .A1(D[2]), .A2(n70), .B1(A[2]), .B2(n69), .ZN(n56) );
  AOI22_X1 U35 ( .A1(D[5]), .A2(n70), .B1(A[5]), .B2(n69), .ZN(n62) );
  AOI22_X1 U36 ( .A1(D[3]), .A2(n70), .B1(A[3]), .B2(n69), .ZN(n58) );
  AOI22_X1 U37 ( .A1(D[1]), .A2(n70), .B1(A[1]), .B2(n69), .ZN(n54) );
  AOI22_X1 U54 ( .A1(D[0]), .A2(n70), .B1(A[0]), .B2(n69), .ZN(n40) );
endmodule


module REG_N16_1_3 ( D, Q, EN, RST, CLK );
  input [15:0] D;
  output [15:0] Q;
  input EN, RST, CLK;
  wire   n1, n2, n3, n4;

  FD_1_48 FF_0 ( .D(D[0]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[0]) );
  FD_1_47 FF_1 ( .D(D[1]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[1]) );
  FD_1_46 FF_2 ( .D(D[2]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[2]) );
  FD_1_45 FF_3 ( .D(D[3]), .CLK(CLK), .EN(n1), .RST(n3), .Q(Q[3]) );
  FD_1_44 FF_4 ( .D(D[4]), .CLK(CLK), .EN(n1), .RST(n3), .Q(Q[4]) );
  FD_1_43 FF_5 ( .D(D[5]), .CLK(CLK), .EN(n1), .RST(n3), .Q(Q[5]) );
  FD_1_42 FF_6 ( .D(D[6]), .CLK(CLK), .EN(n1), .RST(n3), .Q(Q[6]) );
  FD_1_41 FF_7 ( .D(D[7]), .CLK(CLK), .EN(n1), .RST(n3), .Q(Q[7]) );
  FD_1_40 FF_8 ( .D(D[8]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[8]) );
  FD_1_39 FF_9 ( .D(D[9]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[9]) );
  FD_1_38 FF_10 ( .D(D[10]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[10]) );
  FD_1_37 FF_11 ( .D(D[11]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[11]) );
  FD_1_36 FF_12 ( .D(D[12]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[12]) );
  FD_1_35 FF_13 ( .D(D[13]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[13]) );
  FD_1_34 FF_14 ( .D(D[14]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[14]) );
  FD_1_33 FF_15 ( .D(D[15]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[15]) );
  BUF_X1 U1 ( .A(RST), .Z(n3) );
  BUF_X1 U2 ( .A(RST), .Z(n4) );
  CLKBUF_X1 U3 ( .A(EN), .Z(n1) );
  CLKBUF_X1 U4 ( .A(EN), .Z(n2) );
endmodule


module REG_N16_1_2 ( D, Q, EN, RST, CLK );
  input [15:0] D;
  output [15:0] Q;
  input EN, RST, CLK;
  wire   n1, n2;

  FD_1_32 FF_0 ( .D(D[0]), .CLK(CLK), .EN(n1), .RST(RST), .Q(Q[0]) );
  FD_1_31 FF_1 ( .D(D[1]), .CLK(CLK), .EN(n1), .RST(RST), .Q(Q[1]) );
  FD_1_30 FF_2 ( .D(D[2]), .CLK(CLK), .EN(n1), .RST(RST), .Q(Q[2]) );
  FD_1_29 FF_3 ( .D(D[3]), .CLK(CLK), .EN(n1), .RST(RST), .Q(Q[3]) );
  FD_1_28 FF_4 ( .D(D[4]), .CLK(CLK), .EN(n1), .RST(RST), .Q(Q[4]) );
  FD_1_27 FF_5 ( .D(D[5]), .CLK(CLK), .EN(n1), .RST(RST), .Q(Q[5]) );
  FD_1_26 FF_6 ( .D(D[6]), .CLK(CLK), .EN(n1), .RST(RST), .Q(Q[6]) );
  FD_1_25 FF_7 ( .D(D[7]), .CLK(CLK), .EN(n1), .RST(RST), .Q(Q[7]) );
  FD_1_24 FF_8 ( .D(D[8]), .CLK(CLK), .EN(n2), .RST(RST), .Q(Q[8]) );
  FD_1_23 FF_9 ( .D(D[9]), .CLK(CLK), .EN(n2), .RST(RST), .Q(Q[9]) );
  FD_1_22 FF_10 ( .D(D[10]), .CLK(CLK), .EN(n2), .RST(RST), .Q(Q[10]) );
  FD_1_21 FF_11 ( .D(D[11]), .CLK(CLK), .EN(n2), .RST(RST), .Q(Q[11]) );
  FD_1_20 FF_12 ( .D(D[12]), .CLK(CLK), .EN(n2), .RST(RST), .Q(Q[12]) );
  FD_1_19 FF_13 ( .D(D[13]), .CLK(CLK), .EN(n2), .RST(RST), .Q(Q[13]) );
  FD_1_18 FF_14 ( .D(D[14]), .CLK(CLK), .EN(n2), .RST(RST), .Q(Q[14]) );
  FD_1_17 FF_15 ( .D(D[15]), .CLK(CLK), .EN(n2), .RST(RST), .Q(Q[15]) );
  CLKBUF_X1 U1 ( .A(EN), .Z(n1) );
  CLKBUF_X1 U2 ( .A(EN), .Z(n2) );
endmodule


module REG_N16_1_1 ( D, Q, EN, RST, CLK );
  input [15:0] D;
  output [15:0] Q;
  input EN, RST, CLK;
  wire   n1, n2, n3, n4;

  FD_1_16 FF_0 ( .D(D[0]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[0]) );
  FD_1_15 FF_1 ( .D(D[1]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[1]) );
  FD_1_14 FF_2 ( .D(D[2]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[2]) );
  FD_1_13 FF_3 ( .D(D[3]), .CLK(CLK), .EN(n1), .RST(n3), .Q(Q[3]) );
  FD_1_12 FF_4 ( .D(D[4]), .CLK(CLK), .EN(n1), .RST(n3), .Q(Q[4]) );
  FD_1_11 FF_5 ( .D(D[5]), .CLK(CLK), .EN(n1), .RST(n3), .Q(Q[5]) );
  FD_1_10 FF_6 ( .D(D[6]), .CLK(CLK), .EN(n1), .RST(n3), .Q(Q[6]) );
  FD_1_9 FF_7 ( .D(D[7]), .CLK(CLK), .EN(n1), .RST(n3), .Q(Q[7]) );
  FD_1_8 FF_8 ( .D(D[8]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[8]) );
  FD_1_7 FF_9 ( .D(D[9]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[9]) );
  FD_1_6 FF_10 ( .D(D[10]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[10]) );
  FD_1_5 FF_11 ( .D(D[11]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[11]) );
  FD_1_4 FF_12 ( .D(D[12]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[12]) );
  FD_1_3 FF_13 ( .D(D[13]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[13]) );
  FD_1_2 FF_14 ( .D(D[14]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[14]) );
  FD_1_1 FF_15 ( .D(D[15]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[15]) );
  BUF_X1 U1 ( .A(RST), .Z(n3) );
  BUF_X1 U2 ( .A(RST), .Z(n4) );
  CLKBUF_X1 U3 ( .A(EN), .Z(n1) );
  CLKBUF_X1 U4 ( .A(EN), .Z(n2) );
endmodule


module MUX21_GEN_N16_2 ( A, B, SEL, Y );
  input [15:0] A;
  input [15:0] B;
  output [15:0] Y;
  input SEL;
  wire   SB;
  wire   [15:0] Y1;
  wire   [15:0] Y2;

  INV_1_10 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_192 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_191 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_190 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_189 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_188 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_187 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_186 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_185 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_184 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_183 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_182 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_181 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_180 UND1_4 ( .A(A[4]), .B(SEL), .Y(Y1[4]) );
  NAND_GATE_179 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  NAND_GATE_178 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_177 UND1_5 ( .A(A[5]), .B(SEL), .Y(Y1[5]) );
  NAND_GATE_176 UND2_5 ( .A(B[5]), .B(SB), .Y(Y2[5]) );
  NAND_GATE_175 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_174 UND1_6 ( .A(A[6]), .B(SEL), .Y(Y1[6]) );
  NAND_GATE_173 UND2_6 ( .A(B[6]), .B(SB), .Y(Y2[6]) );
  NAND_GATE_172 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_171 UND1_7 ( .A(A[7]), .B(SEL), .Y(Y1[7]) );
  NAND_GATE_170 UND2_7 ( .A(B[7]), .B(SB), .Y(Y2[7]) );
  NAND_GATE_169 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  NAND_GATE_168 UND1_8 ( .A(A[8]), .B(SEL), .Y(Y1[8]) );
  NAND_GATE_167 UND2_8 ( .A(B[8]), .B(SB), .Y(Y2[8]) );
  NAND_GATE_166 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  NAND_GATE_165 UND1_9 ( .A(A[9]), .B(SEL), .Y(Y1[9]) );
  NAND_GATE_164 UND2_9 ( .A(B[9]), .B(SB), .Y(Y2[9]) );
  NAND_GATE_163 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  NAND_GATE_162 UND1_10 ( .A(A[10]), .B(SEL), .Y(Y1[10]) );
  NAND_GATE_161 UND2_10 ( .A(B[10]), .B(SB), .Y(Y2[10]) );
  NAND_GATE_160 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  NAND_GATE_159 UND1_11 ( .A(A[11]), .B(SEL), .Y(Y1[11]) );
  NAND_GATE_158 UND2_11 ( .A(B[11]), .B(SB), .Y(Y2[11]) );
  NAND_GATE_157 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  NAND_GATE_156 UND1_12 ( .A(A[12]), .B(SEL), .Y(Y1[12]) );
  NAND_GATE_155 UND2_12 ( .A(B[12]), .B(SB), .Y(Y2[12]) );
  NAND_GATE_154 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  NAND_GATE_153 UND1_13 ( .A(A[13]), .B(SEL), .Y(Y1[13]) );
  NAND_GATE_152 UND2_13 ( .A(B[13]), .B(SB), .Y(Y2[13]) );
  NAND_GATE_151 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  NAND_GATE_150 UND1_14 ( .A(A[14]), .B(SEL), .Y(Y1[14]) );
  NAND_GATE_149 UND2_14 ( .A(B[14]), .B(SB), .Y(Y2[14]) );
  NAND_GATE_148 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  NAND_GATE_147 UND1_15 ( .A(A[15]), .B(SEL), .Y(Y1[15]) );
  NAND_GATE_146 UND2_15 ( .A(B[15]), .B(SB), .Y(Y2[15]) );
  NAND_GATE_145 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
endmodule


module MUX21_GEN_N16_1 ( A, B, SEL, Y );
  input [15:0] A;
  input [15:0] B;
  output [15:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4;
  wire   [15:0] Y1;
  wire   [15:0] Y2;

  INV_1_9 UIV ( .A(n1), .Y(SB) );
  NAND_GATE_144 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  NAND_GATE_143 UND2_0 ( .A(B[0]), .B(n4), .Y(Y2[0]) );
  NAND_GATE_142 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_141 UND1_1 ( .A(A[1]), .B(n1), .Y(Y1[1]) );
  NAND_GATE_140 UND2_1 ( .A(B[1]), .B(n4), .Y(Y2[1]) );
  NAND_GATE_139 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_138 UND1_2 ( .A(A[2]), .B(n1), .Y(Y1[2]) );
  NAND_GATE_137 UND2_2 ( .A(B[2]), .B(n4), .Y(Y2[2]) );
  NAND_GATE_136 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_135 UND1_3 ( .A(A[3]), .B(n1), .Y(Y1[3]) );
  NAND_GATE_134 UND2_3 ( .A(B[3]), .B(n3), .Y(Y2[3]) );
  NAND_GATE_133 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_132 UND1_4 ( .A(A[4]), .B(n1), .Y(Y1[4]) );
  NAND_GATE_131 UND2_4 ( .A(B[4]), .B(n3), .Y(Y2[4]) );
  NAND_GATE_130 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_129 UND1_5 ( .A(A[5]), .B(n1), .Y(Y1[5]) );
  NAND_GATE_128 UND2_5 ( .A(B[5]), .B(n3), .Y(Y2[5]) );
  NAND_GATE_127 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_126 UND1_6 ( .A(A[6]), .B(n1), .Y(Y1[6]) );
  NAND_GATE_125 UND2_6 ( .A(B[6]), .B(n3), .Y(Y2[6]) );
  NAND_GATE_124 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_123 UND1_7 ( .A(A[7]), .B(n1), .Y(Y1[7]) );
  NAND_GATE_122 UND2_7 ( .A(B[7]), .B(n3), .Y(Y2[7]) );
  NAND_GATE_121 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  NAND_GATE_120 UND1_8 ( .A(A[8]), .B(n1), .Y(Y1[8]) );
  NAND_GATE_119 UND2_8 ( .A(B[8]), .B(n3), .Y(Y2[8]) );
  NAND_GATE_118 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  NAND_GATE_117 UND1_9 ( .A(A[9]), .B(n1), .Y(Y1[9]) );
  NAND_GATE_116 UND2_9 ( .A(B[9]), .B(n3), .Y(Y2[9]) );
  NAND_GATE_115 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  NAND_GATE_114 UND1_10 ( .A(A[10]), .B(n1), .Y(Y1[10]) );
  NAND_GATE_113 UND2_10 ( .A(B[10]), .B(n3), .Y(Y2[10]) );
  NAND_GATE_112 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  NAND_GATE_111 UND1_11 ( .A(A[11]), .B(n1), .Y(Y1[11]) );
  NAND_GATE_110 UND2_11 ( .A(B[11]), .B(n3), .Y(Y2[11]) );
  NAND_GATE_109 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  NAND_GATE_108 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  NAND_GATE_107 UND2_12 ( .A(B[12]), .B(n3), .Y(Y2[12]) );
  NAND_GATE_106 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  NAND_GATE_105 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  NAND_GATE_104 UND2_13 ( .A(B[13]), .B(n3), .Y(Y2[13]) );
  NAND_GATE_103 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  NAND_GATE_102 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  NAND_GATE_101 UND2_14 ( .A(B[14]), .B(n3), .Y(Y2[14]) );
  NAND_GATE_100 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  NAND_GATE_99 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  NAND_GATE_98 UND2_15 ( .A(B[15]), .B(n3), .Y(Y2[15]) );
  NAND_GATE_97 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  BUF_X1 U1 ( .A(SB), .Z(n3) );
  BUF_X1 U2 ( .A(SB), .Z(n4) );
  BUF_X1 U3 ( .A(SEL), .Z(n1) );
  BUF_X1 U4 ( .A(SEL), .Z(n2) );
endmodule


module BOOTH_ENCODER_7 ( TO_ENC, ENC );
  input [2:0] TO_ENC;
  output [2:0] ENC;
  wire   n1, n2, n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(TO_ENC[2]), .ZN(n4) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(n2) );
  NAND2_X1 U3 ( .A1(n1), .A2(TO_ENC[2]), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n2), .A2(n3), .ZN(ENC[1]) );
  INV_X1 U5 ( .A(n5), .ZN(n1) );
  NAND2_X2 U6 ( .A1(TO_ENC[0]), .A2(TO_ENC[1]), .ZN(n5) );
  INV_X1 U7 ( .A(TO_ENC[1]), .ZN(n6) );
  OAI21_X1 U8 ( .B1(TO_ENC[0]), .B2(TO_ENC[1]), .A(n4), .ZN(ENC[0]) );
  INV_X1 U9 ( .A(TO_ENC[0]), .ZN(n7) );
  NAND3_X1 U10 ( .A1(TO_ENC[2]), .A2(n7), .A3(n6), .ZN(ENC[2]) );
endmodule


module BOOTH_ENCODER_6 ( TO_ENC, ENC );
  input [2:0] TO_ENC;
  output [2:0] ENC;
  wire   n3, n4;

  NAND2_X1 U3 ( .A1(TO_ENC[2]), .A2(n4), .ZN(ENC[2]) );
  XOR2_X1 U4 ( .A(n3), .B(TO_ENC[2]), .Z(ENC[1]) );
  NAND2_X1 U5 ( .A1(TO_ENC[0]), .A2(TO_ENC[1]), .ZN(n3) );
  NOR2_X1 U1 ( .A1(TO_ENC[0]), .A2(TO_ENC[1]), .ZN(n4) );
  OR2_X1 U2 ( .A1(n4), .A2(TO_ENC[2]), .ZN(ENC[0]) );
endmodule


module BOOTH_ENCODER_5 ( TO_ENC, ENC );
  input [2:0] TO_ENC;
  output [2:0] ENC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;

  NAND2_X2 U1 ( .A1(TO_ENC[1]), .A2(TO_ENC[0]), .ZN(n6) );
  INV_X2 U2 ( .A(TO_ENC[2]), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n6), .A2(n5), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n1), .A2(n2), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n3), .A2(n4), .ZN(ENC[1]) );
  INV_X1 U6 ( .A(n6), .ZN(n1) );
  INV_X1 U7 ( .A(n5), .ZN(n2) );
  OAI21_X1 U8 ( .B1(TO_ENC[0]), .B2(TO_ENC[1]), .A(n5), .ZN(ENC[0]) );
  INV_X1 U9 ( .A(TO_ENC[0]), .ZN(n8) );
  INV_X1 U10 ( .A(TO_ENC[1]), .ZN(n7) );
  NAND3_X1 U11 ( .A1(TO_ENC[2]), .A2(n8), .A3(n7), .ZN(ENC[2]) );
endmodule


module BOOTH_ENCODER_4 ( TO_ENC, ENC );
  input [2:0] TO_ENC;
  output [2:0] ENC;
  wire   n3, n4;

  NAND2_X1 U3 ( .A1(TO_ENC[2]), .A2(n4), .ZN(ENC[2]) );
  XOR2_X1 U4 ( .A(n3), .B(TO_ENC[2]), .Z(ENC[1]) );
  NAND2_X1 U5 ( .A1(TO_ENC[0]), .A2(TO_ENC[1]), .ZN(n3) );
  OR2_X1 U1 ( .A1(n4), .A2(TO_ENC[2]), .ZN(ENC[0]) );
  NOR2_X1 U2 ( .A1(TO_ENC[0]), .A2(TO_ENC[1]), .ZN(n4) );
endmodule


module BOOTH_ENCODER_3 ( TO_ENC, ENC );
  input [2:0] TO_ENC;
  output [2:0] ENC;
  wire   n3, n4;

  NAND2_X1 U3 ( .A1(TO_ENC[2]), .A2(n4), .ZN(ENC[2]) );
  XOR2_X1 U4 ( .A(n3), .B(TO_ENC[2]), .Z(ENC[1]) );
  NAND2_X1 U5 ( .A1(TO_ENC[0]), .A2(TO_ENC[1]), .ZN(n3) );
  OR2_X1 U1 ( .A1(n4), .A2(TO_ENC[2]), .ZN(ENC[0]) );
  NOR2_X1 U2 ( .A1(TO_ENC[0]), .A2(TO_ENC[1]), .ZN(n4) );
endmodule


module BOOTH_ENCODER_2 ( TO_ENC, ENC );
  input [2:0] TO_ENC;
  output [2:0] ENC;
  wire   n2, n3;

  OR2_X2 U1 ( .A1(n3), .A2(TO_ENC[2]), .ZN(ENC[0]) );
  NAND2_X1 U2 ( .A1(TO_ENC[2]), .A2(n3), .ZN(ENC[2]) );
  AND2_X2 U3 ( .A1(TO_ENC[0]), .A2(TO_ENC[1]), .ZN(n2) );
  XNOR2_X2 U4 ( .A(n2), .B(TO_ENC[2]), .ZN(ENC[1]) );
  NOR2_X1 U5 ( .A1(TO_ENC[0]), .A2(TO_ENC[1]), .ZN(n3) );
endmodule


module BOOTH_ENCODER_1 ( TO_ENC, ENC );
  input [2:0] TO_ENC;
  output [2:0] ENC;
  wire   n3, n4;

  NAND2_X1 U3 ( .A1(TO_ENC[2]), .A2(n4), .ZN(ENC[2]) );
  XOR2_X1 U4 ( .A(n3), .B(TO_ENC[2]), .Z(ENC[1]) );
  NAND2_X1 U5 ( .A1(TO_ENC[0]), .A2(TO_ENC[1]), .ZN(n3) );
  OR2_X1 U1 ( .A1(n4), .A2(TO_ENC[2]), .ZN(ENC[0]) );
  NOR2_X1 U2 ( .A1(TO_ENC[0]), .A2(TO_ENC[1]), .ZN(n4) );
endmodule


module RCA_GEN_NO_C_N19_6 ( A, B, S, Co );
  input [18:0] A;
  input [18:0] B;
  output [18:0] S;
  output Co;

  wire   [17:0] CTMP;

  HA_6 HA_INST ( .A(A[0]), .B(B[0]), .S(S[0]), .Co(CTMP[0]) );
  FA_172 FAI_0 ( .A(A[1]), .B(B[1]), .Ci(CTMP[0]), .S(S[1]), .Co(CTMP[1]) );
  FA_171 FAI_1 ( .A(A[2]), .B(B[2]), .Ci(CTMP[1]), .S(S[2]), .Co(CTMP[2]) );
  FA_170 FAI_2 ( .A(A[3]), .B(B[3]), .Ci(CTMP[2]), .S(S[3]), .Co(CTMP[3]) );
  FA_169 FAI_3 ( .A(A[4]), .B(B[4]), .Ci(CTMP[3]), .S(S[4]), .Co(CTMP[4]) );
  FA_168 FAI_4 ( .A(A[5]), .B(B[5]), .Ci(CTMP[4]), .S(S[5]), .Co(CTMP[5]) );
  FA_167 FAI_5 ( .A(A[6]), .B(B[6]), .Ci(CTMP[5]), .S(S[6]), .Co(CTMP[6]) );
  FA_166 FAI_6 ( .A(A[7]), .B(B[7]), .Ci(CTMP[6]), .S(S[7]), .Co(CTMP[7]) );
  FA_165 FAI_7 ( .A(A[8]), .B(B[8]), .Ci(CTMP[7]), .S(S[8]), .Co(CTMP[8]) );
  FA_164 FAI_8 ( .A(A[9]), .B(B[9]), .Ci(CTMP[8]), .S(S[9]), .Co(CTMP[9]) );
  FA_163 FAI_9 ( .A(A[10]), .B(B[10]), .Ci(CTMP[9]), .S(S[10]), .Co(CTMP[10])
         );
  FA_162 FAI_10 ( .A(A[11]), .B(B[11]), .Ci(CTMP[10]), .S(S[11]), .Co(CTMP[11]) );
  FA_161 FAI_11 ( .A(A[12]), .B(B[12]), .Ci(CTMP[11]), .S(S[12]), .Co(CTMP[12]) );
  FA_160 FAI_12 ( .A(A[13]), .B(B[13]), .Ci(CTMP[12]), .S(S[13]), .Co(CTMP[13]) );
  FA_159 FAI_13 ( .A(A[14]), .B(B[14]), .Ci(CTMP[13]), .S(S[14]), .Co(CTMP[14]) );
  FA_158 FAI_14 ( .A(A[15]), .B(B[15]), .Ci(CTMP[14]), .S(S[15]), .Co(CTMP[15]) );
  FA_157 FAI_15 ( .A(A[16]), .B(B[16]), .Ci(CTMP[15]), .S(S[16]), .Co(CTMP[16]) );
  FA_156 FAI_16 ( .A(A[17]), .B(B[17]), .Ci(CTMP[16]), .S(S[17]), .Co(CTMP[17]) );
  FA_155 FAI_17 ( .A(A[18]), .B(B[18]), .Ci(CTMP[17]), .S(S[18]), .Co(Co) );
endmodule


module RCA_GEN_NO_C_N19_5 ( A, B, S, Co );
  input [18:0] A;
  input [18:0] B;
  output [18:0] S;
  output Co;

  wire   [17:0] CTMP;

  HA_5 HA_INST ( .A(A[0]), .B(B[0]), .S(S[0]), .Co(CTMP[0]) );
  FA_154 FAI_0 ( .A(A[1]), .B(B[1]), .Ci(CTMP[0]), .S(S[1]), .Co(CTMP[1]) );
  FA_153 FAI_1 ( .A(A[2]), .B(B[2]), .Ci(CTMP[1]), .S(S[2]), .Co(CTMP[2]) );
  FA_152 FAI_2 ( .A(A[3]), .B(B[3]), .Ci(CTMP[2]), .S(S[3]), .Co(CTMP[3]) );
  FA_151 FAI_3 ( .A(A[4]), .B(B[4]), .Ci(CTMP[3]), .S(S[4]), .Co(CTMP[4]) );
  FA_150 FAI_4 ( .A(A[5]), .B(B[5]), .Ci(CTMP[4]), .S(S[5]), .Co(CTMP[5]) );
  FA_149 FAI_5 ( .A(A[6]), .B(B[6]), .Ci(CTMP[5]), .S(S[6]), .Co(CTMP[6]) );
  FA_148 FAI_6 ( .A(A[7]), .B(B[7]), .Ci(CTMP[6]), .S(S[7]), .Co(CTMP[7]) );
  FA_147 FAI_7 ( .A(A[8]), .B(B[8]), .Ci(CTMP[7]), .S(S[8]), .Co(CTMP[8]) );
  FA_146 FAI_8 ( .A(A[9]), .B(B[9]), .Ci(CTMP[8]), .S(S[9]), .Co(CTMP[9]) );
  FA_145 FAI_9 ( .A(A[10]), .B(B[10]), .Ci(CTMP[9]), .S(S[10]), .Co(CTMP[10])
         );
  FA_144 FAI_10 ( .A(A[11]), .B(B[11]), .Ci(CTMP[10]), .S(S[11]), .Co(CTMP[11]) );
  FA_143 FAI_11 ( .A(A[12]), .B(B[12]), .Ci(CTMP[11]), .S(S[12]), .Co(CTMP[12]) );
  FA_142 FAI_12 ( .A(A[13]), .B(B[13]), .Ci(CTMP[12]), .S(S[13]), .Co(CTMP[13]) );
  FA_141 FAI_13 ( .A(A[14]), .B(B[14]), .Ci(CTMP[13]), .S(S[14]), .Co(CTMP[14]) );
  FA_140 FAI_14 ( .A(A[15]), .B(B[15]), .Ci(CTMP[14]), .S(S[15]), .Co(CTMP[15]) );
  FA_139 FAI_15 ( .A(A[16]), .B(B[16]), .Ci(CTMP[15]), .S(S[16]), .Co(CTMP[16]) );
  FA_138 FAI_16 ( .A(A[17]), .B(B[17]), .Ci(CTMP[16]), .S(S[17]), .Co(CTMP[17]) );
  FA_137 FAI_17 ( .A(A[18]), .B(B[18]), .Ci(CTMP[17]), .S(S[18]), .Co(Co) );
endmodule


module RCA_GEN_NO_C_N19_4 ( A, B, S, Co );
  input [18:0] A;
  input [18:0] B;
  output [18:0] S;
  output Co;

  wire   [17:0] CTMP;

  HA_4 HA_INST ( .A(A[0]), .B(B[0]), .S(S[0]), .Co(CTMP[0]) );
  FA_136 FAI_0 ( .A(A[1]), .B(B[1]), .Ci(CTMP[0]), .S(S[1]), .Co(CTMP[1]) );
  FA_135 FAI_1 ( .A(A[2]), .B(B[2]), .Ci(CTMP[1]), .S(S[2]), .Co(CTMP[2]) );
  FA_134 FAI_2 ( .A(A[3]), .B(B[3]), .Ci(CTMP[2]), .S(S[3]), .Co(CTMP[3]) );
  FA_133 FAI_3 ( .A(A[4]), .B(B[4]), .Ci(CTMP[3]), .S(S[4]), .Co(CTMP[4]) );
  FA_132 FAI_4 ( .A(A[5]), .B(B[5]), .Ci(CTMP[4]), .S(S[5]), .Co(CTMP[5]) );
  FA_131 FAI_5 ( .A(A[6]), .B(B[6]), .Ci(CTMP[5]), .S(S[6]), .Co(CTMP[6]) );
  FA_130 FAI_6 ( .A(A[7]), .B(B[7]), .Ci(CTMP[6]), .S(S[7]), .Co(CTMP[7]) );
  FA_129 FAI_7 ( .A(A[8]), .B(B[8]), .Ci(CTMP[7]), .S(S[8]), .Co(CTMP[8]) );
  FA_128 FAI_8 ( .A(A[9]), .B(B[9]), .Ci(CTMP[8]), .S(S[9]), .Co(CTMP[9]) );
  FA_127 FAI_9 ( .A(A[10]), .B(B[10]), .Ci(CTMP[9]), .S(S[10]), .Co(CTMP[10])
         );
  FA_126 FAI_10 ( .A(A[11]), .B(B[11]), .Ci(CTMP[10]), .S(S[11]), .Co(CTMP[11]) );
  FA_125 FAI_11 ( .A(A[12]), .B(B[12]), .Ci(CTMP[11]), .S(S[12]), .Co(CTMP[12]) );
  FA_124 FAI_12 ( .A(A[13]), .B(B[13]), .Ci(CTMP[12]), .S(S[13]), .Co(CTMP[13]) );
  FA_123 FAI_13 ( .A(A[14]), .B(B[14]), .Ci(CTMP[13]), .S(S[14]), .Co(CTMP[14]) );
  FA_122 FAI_14 ( .A(A[15]), .B(B[15]), .Ci(CTMP[14]), .S(S[15]), .Co(CTMP[15]) );
  FA_121 FAI_15 ( .A(A[16]), .B(B[16]), .Ci(CTMP[15]), .S(S[16]), .Co(CTMP[16]) );
  FA_120 FAI_16 ( .A(A[17]), .B(B[17]), .Ci(CTMP[16]), .S(S[17]), .Co(CTMP[17]) );
  FA_119 FAI_17 ( .A(A[18]), .B(B[18]), .Ci(CTMP[17]), .S(S[18]), .Co(Co) );
endmodule


module RCA_GEN_NO_C_N19_3 ( A, B, S, Co );
  input [18:0] A;
  input [18:0] B;
  output [18:0] S;
  output Co;

  wire   [17:0] CTMP;

  HA_3 HA_INST ( .A(A[0]), .B(B[0]), .S(S[0]), .Co(CTMP[0]) );
  FA_118 FAI_0 ( .A(A[1]), .B(B[1]), .Ci(CTMP[0]), .S(S[1]), .Co(CTMP[1]) );
  FA_117 FAI_1 ( .A(A[2]), .B(B[2]), .Ci(CTMP[1]), .S(S[2]), .Co(CTMP[2]) );
  FA_116 FAI_2 ( .A(A[3]), .B(B[3]), .Ci(CTMP[2]), .S(S[3]), .Co(CTMP[3]) );
  FA_115 FAI_3 ( .A(A[4]), .B(B[4]), .Ci(CTMP[3]), .S(S[4]), .Co(CTMP[4]) );
  FA_114 FAI_4 ( .A(A[5]), .B(B[5]), .Ci(CTMP[4]), .S(S[5]), .Co(CTMP[5]) );
  FA_113 FAI_5 ( .A(A[6]), .B(B[6]), .Ci(CTMP[5]), .S(S[6]), .Co(CTMP[6]) );
  FA_112 FAI_6 ( .A(A[7]), .B(B[7]), .Ci(CTMP[6]), .S(S[7]), .Co(CTMP[7]) );
  FA_111 FAI_7 ( .A(A[8]), .B(B[8]), .Ci(CTMP[7]), .S(S[8]), .Co(CTMP[8]) );
  FA_110 FAI_8 ( .A(A[9]), .B(B[9]), .Ci(CTMP[8]), .S(S[9]), .Co(CTMP[9]) );
  FA_109 FAI_9 ( .A(A[10]), .B(B[10]), .Ci(CTMP[9]), .S(S[10]), .Co(CTMP[10])
         );
  FA_108 FAI_10 ( .A(A[11]), .B(B[11]), .Ci(CTMP[10]), .S(S[11]), .Co(CTMP[11]) );
  FA_107 FAI_11 ( .A(A[12]), .B(B[12]), .Ci(CTMP[11]), .S(S[12]), .Co(CTMP[12]) );
  FA_106 FAI_12 ( .A(A[13]), .B(B[13]), .Ci(CTMP[12]), .S(S[13]), .Co(CTMP[13]) );
  FA_105 FAI_13 ( .A(A[14]), .B(B[14]), .Ci(CTMP[13]), .S(S[14]), .Co(CTMP[14]) );
  FA_104 FAI_14 ( .A(A[15]), .B(B[15]), .Ci(CTMP[14]), .S(S[15]), .Co(CTMP[15]) );
  FA_103 FAI_15 ( .A(A[16]), .B(B[16]), .Ci(CTMP[15]), .S(S[16]), .Co(CTMP[16]) );
  FA_102 FAI_16 ( .A(A[17]), .B(B[17]), .Ci(CTMP[16]), .S(S[17]), .Co(CTMP[17]) );
  FA_101 FAI_17 ( .A(A[18]), .B(B[18]), .Ci(CTMP[17]), .S(S[18]), .Co(Co) );
endmodule


module RCA_GEN_NO_C_N19_2 ( A, B, S, Co );
  input [18:0] A;
  input [18:0] B;
  output [18:0] S;
  output Co;

  wire   [17:0] CTMP;

  HA_2 HA_INST ( .A(A[0]), .B(B[0]), .S(S[0]), .Co(CTMP[0]) );
  FA_100 FAI_0 ( .A(A[1]), .B(B[1]), .Ci(CTMP[0]), .S(S[1]), .Co(CTMP[1]) );
  FA_99 FAI_1 ( .A(A[2]), .B(B[2]), .Ci(CTMP[1]), .S(S[2]), .Co(CTMP[2]) );
  FA_98 FAI_2 ( .A(A[3]), .B(B[3]), .Ci(CTMP[2]), .S(S[3]), .Co(CTMP[3]) );
  FA_97 FAI_3 ( .A(A[4]), .B(B[4]), .Ci(CTMP[3]), .S(S[4]), .Co(CTMP[4]) );
  FA_96 FAI_4 ( .A(A[5]), .B(B[5]), .Ci(CTMP[4]), .S(S[5]), .Co(CTMP[5]) );
  FA_95 FAI_5 ( .A(A[6]), .B(B[6]), .Ci(CTMP[5]), .S(S[6]), .Co(CTMP[6]) );
  FA_94 FAI_6 ( .A(A[7]), .B(B[7]), .Ci(CTMP[6]), .S(S[7]), .Co(CTMP[7]) );
  FA_93 FAI_7 ( .A(A[8]), .B(B[8]), .Ci(CTMP[7]), .S(S[8]), .Co(CTMP[8]) );
  FA_92 FAI_8 ( .A(A[9]), .B(B[9]), .Ci(CTMP[8]), .S(S[9]), .Co(CTMP[9]) );
  FA_91 FAI_9 ( .A(A[10]), .B(B[10]), .Ci(CTMP[9]), .S(S[10]), .Co(CTMP[10])
         );
  FA_90 FAI_10 ( .A(A[11]), .B(B[11]), .Ci(CTMP[10]), .S(S[11]), .Co(CTMP[11])
         );
  FA_89 FAI_11 ( .A(A[12]), .B(B[12]), .Ci(CTMP[11]), .S(S[12]), .Co(CTMP[12])
         );
  FA_88 FAI_12 ( .A(A[13]), .B(B[13]), .Ci(CTMP[12]), .S(S[13]), .Co(CTMP[13])
         );
  FA_87 FAI_13 ( .A(A[14]), .B(B[14]), .Ci(CTMP[13]), .S(S[14]), .Co(CTMP[14])
         );
  FA_86 FAI_14 ( .A(A[15]), .B(B[15]), .Ci(CTMP[14]), .S(S[15]), .Co(CTMP[15])
         );
  FA_85 FAI_15 ( .A(A[16]), .B(B[16]), .Ci(CTMP[15]), .S(S[16]), .Co(CTMP[16])
         );
  FA_84 FAI_16 ( .A(A[17]), .B(B[17]), .Ci(CTMP[16]), .S(S[17]), .Co(CTMP[17])
         );
  FA_83 FAI_17 ( .A(A[18]), .B(B[18]), .Ci(CTMP[17]), .S(S[18]), .Co(Co) );
endmodule


module RCA_GEN_NO_C_N19_1 ( A, B, S, Co );
  input [18:0] A;
  input [18:0] B;
  output [18:0] S;
  output Co;

  wire   [17:0] CTMP;

  HA_1 HA_INST ( .A(A[0]), .B(B[0]), .S(S[0]), .Co(CTMP[0]) );
  FA_82 FAI_0 ( .A(A[1]), .B(B[1]), .Ci(CTMP[0]), .S(S[1]), .Co(CTMP[1]) );
  FA_81 FAI_1 ( .A(A[2]), .B(B[2]), .Ci(CTMP[1]), .S(S[2]), .Co(CTMP[2]) );
  FA_80 FAI_2 ( .A(A[3]), .B(B[3]), .Ci(CTMP[2]), .S(S[3]), .Co(CTMP[3]) );
  FA_79 FAI_3 ( .A(A[4]), .B(B[4]), .Ci(CTMP[3]), .S(S[4]), .Co(CTMP[4]) );
  FA_78 FAI_4 ( .A(A[5]), .B(B[5]), .Ci(CTMP[4]), .S(S[5]), .Co(CTMP[5]) );
  FA_77 FAI_5 ( .A(A[6]), .B(B[6]), .Ci(CTMP[5]), .S(S[6]), .Co(CTMP[6]) );
  FA_76 FAI_6 ( .A(A[7]), .B(B[7]), .Ci(CTMP[6]), .S(S[7]), .Co(CTMP[7]) );
  FA_75 FAI_7 ( .A(A[8]), .B(B[8]), .Ci(CTMP[7]), .S(S[8]), .Co(CTMP[8]) );
  FA_74 FAI_8 ( .A(A[9]), .B(B[9]), .Ci(CTMP[8]), .S(S[9]), .Co(CTMP[9]) );
  FA_73 FAI_9 ( .A(A[10]), .B(B[10]), .Ci(CTMP[9]), .S(S[10]), .Co(CTMP[10])
         );
  FA_72 FAI_10 ( .A(A[11]), .B(B[11]), .Ci(CTMP[10]), .S(S[11]), .Co(CTMP[11])
         );
  FA_71 FAI_11 ( .A(A[12]), .B(B[12]), .Ci(CTMP[11]), .S(S[12]), .Co(CTMP[12])
         );
  FA_70 FAI_12 ( .A(A[13]), .B(B[13]), .Ci(CTMP[12]), .S(S[13]), .Co(CTMP[13])
         );
  FA_69 FAI_13 ( .A(A[14]), .B(B[14]), .Ci(CTMP[13]), .S(S[14]), .Co(CTMP[14])
         );
  FA_68 FAI_14 ( .A(A[15]), .B(B[15]), .Ci(CTMP[14]), .S(S[15]), .Co(CTMP[15])
         );
  FA_67 FAI_15 ( .A(A[16]), .B(B[16]), .Ci(CTMP[15]), .S(S[16]), .Co(CTMP[16])
         );
  FA_66 FAI_16 ( .A(A[17]), .B(B[17]), .Ci(CTMP[16]), .S(S[17]), .Co(CTMP[17])
         );
  FA_65 FAI_17 ( .A(A[18]), .B(B[18]), .Ci(CTMP[17]), .S(S[18]), .Co(Co) );
endmodule


module MUX51_GEN_N19_7 ( A, B, C, D, E, SEL, Y );
  input [18:0] A;
  input [18:0] B;
  input [18:0] C;
  input [18:0] D;
  input [18:0] E;
  input [2:0] SEL;
  output [18:0] Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99;

  BUF_X8 U1 ( .A(n93), .Z(n4) );
  AOI22_X2 U2 ( .A1(n94), .A2(E[1]), .B1(n93), .B2(B[1]), .ZN(n19) );
  NOR2_X2 U3 ( .A1(n14), .A2(n13), .ZN(n94) );
  NAND3_X2 U4 ( .A1(n16), .A2(n17), .A3(n18), .ZN(Y[0]) );
  AOI22_X4 U5 ( .A1(E[0]), .A2(n1), .B1(B[0]), .B2(n4), .ZN(n16) );
  NAND3_X1 U6 ( .A1(n19), .A2(n20), .A3(n21), .ZN(Y[1]) );
  INV_X1 U7 ( .A(n92), .ZN(n5) );
  AOI22_X1 U8 ( .A1(C[0]), .A2(n25), .B1(A[0]), .B2(n96), .ZN(n18) );
  INV_X2 U9 ( .A(n5), .ZN(n6) );
  NOR2_X1 U10 ( .A1(n14), .A2(n13), .ZN(n1) );
  INV_X1 U11 ( .A(n11), .ZN(n2) );
  INV_X2 U12 ( .A(n15), .ZN(n93) );
  NAND2_X2 U13 ( .A1(n12), .A2(n32), .ZN(n14) );
  NAND2_X2 U14 ( .A1(n15), .A2(n6), .ZN(n13) );
  NAND2_X2 U15 ( .A1(n2), .A2(n8), .ZN(n12) );
  INV_X4 U16 ( .A(n12), .ZN(n96) );
  INV_X1 U17 ( .A(n32), .ZN(n3) );
  AOI211_X1 U18 ( .C1(E[7]), .C2(n7), .A(n42), .B(n9), .ZN(n43) );
  NAND3_X1 U19 ( .A1(SEL[2]), .A2(n11), .A3(n10), .ZN(n92) );
  CLKBUF_X1 U20 ( .A(n1), .Z(n7) );
  INV_X1 U21 ( .A(n32), .ZN(n95) );
  INV_X1 U22 ( .A(n32), .ZN(n25) );
  INV_X1 U23 ( .A(n6), .ZN(n50) );
  INV_X1 U24 ( .A(n6), .ZN(n55) );
  INV_X1 U25 ( .A(n6), .ZN(n60) );
  INV_X1 U26 ( .A(n6), .ZN(n65) );
  INV_X1 U27 ( .A(n6), .ZN(n70) );
  INV_X1 U28 ( .A(n6), .ZN(n83) );
  NAND3_X1 U29 ( .A1(n2), .A2(SEL[2]), .A3(n10), .ZN(n32) );
  INV_X1 U30 ( .A(SEL[0]), .ZN(n11) );
  AND2_X1 U31 ( .A1(SEL[2]), .A2(SEL[1]), .ZN(n8) );
  NOR2_X1 U32 ( .A1(n6), .A2(n41), .ZN(n42) );
  AND2_X1 U33 ( .A1(B[7]), .A2(n4), .ZN(n9) );
  AOI22_X1 U34 ( .A1(C[2]), .A2(n95), .B1(A[2]), .B2(n96), .ZN(n24) );
  AOI22_X1 U35 ( .A1(E[2]), .A2(n1), .B1(B[2]), .B2(n4), .ZN(n22) );
  AOI22_X1 U36 ( .A1(C[3]), .A2(n95), .B1(A[3]), .B2(n96), .ZN(n28) );
  AOI22_X1 U37 ( .A1(E[3]), .A2(n1), .B1(B[3]), .B2(n4), .ZN(n26) );
  AOI22_X1 U38 ( .A1(E[4]), .A2(n1), .B1(B[4]), .B2(n4), .ZN(n29) );
  AOI22_X1 U39 ( .A1(C[4]), .A2(n95), .B1(A[4]), .B2(n96), .ZN(n31) );
  AOI22_X1 U40 ( .A1(C[1]), .A2(n3), .B1(A[1]), .B2(n96), .ZN(n21) );
  AOI22_X1 U41 ( .A1(E[6]), .A2(n7), .B1(B[6]), .B2(n4), .ZN(n38) );
  AOI22_X1 U42 ( .A1(A[6]), .A2(n96), .B1(C[6]), .B2(n95), .ZN(n40) );
  NAND4_X1 U43 ( .A1(n91), .A2(n90), .A3(n89), .A4(n88), .ZN(Y[17]) );
  AOI22_X1 U44 ( .A1(D[17]), .A2(n83), .B1(B[17]), .B2(n93), .ZN(n91) );
  NAND4_X1 U45 ( .A1(n87), .A2(n86), .A3(n85), .A4(n84), .ZN(Y[16]) );
  AOI22_X1 U46 ( .A1(D[16]), .A2(n83), .B1(B[16]), .B2(n93), .ZN(n87) );
  NAND4_X1 U47 ( .A1(n54), .A2(n53), .A3(n52), .A4(n51), .ZN(Y[9]) );
  AOI22_X1 U48 ( .A1(D[9]), .A2(n50), .B1(B[9]), .B2(n4), .ZN(n54) );
  NAND4_X1 U49 ( .A1(n59), .A2(n58), .A3(n57), .A4(n56), .ZN(Y[10]) );
  AOI22_X1 U50 ( .A1(D[10]), .A2(n55), .B1(B[10]), .B2(n4), .ZN(n59) );
  NAND4_X1 U51 ( .A1(n64), .A2(n63), .A3(n62), .A4(n61), .ZN(Y[11]) );
  AOI22_X1 U52 ( .A1(D[11]), .A2(n60), .B1(B[11]), .B2(n4), .ZN(n64) );
  NAND4_X1 U53 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(Y[12]) );
  AOI22_X1 U54 ( .A1(D[12]), .A2(n65), .B1(B[12]), .B2(n4), .ZN(n69) );
  NAND4_X1 U55 ( .A1(n74), .A2(n73), .A3(n72), .A4(n71), .ZN(Y[13]) );
  AOI22_X1 U56 ( .A1(D[13]), .A2(n70), .B1(B[13]), .B2(n4), .ZN(n74) );
  NAND4_X1 U57 ( .A1(n78), .A2(n77), .A3(n76), .A4(n75), .ZN(Y[14]) );
  AOI22_X1 U58 ( .A1(D[14]), .A2(n83), .B1(B[14]), .B2(n4), .ZN(n78) );
  NAND4_X1 U59 ( .A1(n82), .A2(n81), .A3(n80), .A4(n79), .ZN(Y[15]) );
  AOI22_X1 U60 ( .A1(D[15]), .A2(n83), .B1(B[15]), .B2(n93), .ZN(n82) );
  NAND4_X1 U61 ( .A1(n49), .A2(n48), .A3(n47), .A4(n46), .ZN(Y[8]) );
  AOI22_X1 U62 ( .A1(D[8]), .A2(n50), .B1(B[8]), .B2(n4), .ZN(n49) );
  AOI22_X1 U63 ( .A1(D[18]), .A2(n83), .B1(B[18]), .B2(n93), .ZN(n99) );
  AOI22_X1 U64 ( .A1(A[18]), .A2(n96), .B1(C[18]), .B2(n95), .ZN(n97) );
  INV_X1 U65 ( .A(SEL[1]), .ZN(n10) );
  INV_X1 U66 ( .A(n6), .ZN(n37) );
  NAND2_X1 U67 ( .A1(D[0]), .A2(n37), .ZN(n17) );
  NAND2_X1 U68 ( .A1(n11), .A2(n8), .ZN(n15) );
  NAND2_X1 U69 ( .A1(D[1]), .A2(n37), .ZN(n20) );
  NAND2_X1 U70 ( .A1(D[2]), .A2(n37), .ZN(n23) );
  NAND3_X1 U71 ( .A1(n24), .A2(n23), .A3(n22), .ZN(Y[2]) );
  NAND2_X1 U72 ( .A1(D[3]), .A2(n37), .ZN(n27) );
  NAND3_X1 U73 ( .A1(n28), .A2(n27), .A3(n26), .ZN(Y[3]) );
  NAND2_X1 U74 ( .A1(D[4]), .A2(n37), .ZN(n30) );
  NAND3_X1 U75 ( .A1(n31), .A2(n30), .A3(n29), .ZN(Y[4]) );
  NAND2_X1 U76 ( .A1(E[5]), .A2(n1), .ZN(n36) );
  NAND2_X1 U77 ( .A1(B[5]), .A2(n4), .ZN(n35) );
  NAND2_X1 U78 ( .A1(D[5]), .A2(n37), .ZN(n34) );
  AOI22_X1 U79 ( .A1(C[5]), .A2(n95), .B1(A[5]), .B2(n96), .ZN(n33) );
  NAND4_X1 U80 ( .A1(n36), .A2(n35), .A3(n34), .A4(n33), .ZN(Y[5]) );
  NAND2_X1 U81 ( .A1(D[6]), .A2(n37), .ZN(n39) );
  NAND3_X1 U82 ( .A1(n40), .A2(n39), .A3(n38), .ZN(Y[6]) );
  NAND2_X1 U83 ( .A1(A[7]), .A2(n96), .ZN(n45) );
  NAND2_X1 U84 ( .A1(C[7]), .A2(n95), .ZN(n44) );
  INV_X1 U85 ( .A(D[7]), .ZN(n41) );
  NAND3_X1 U86 ( .A1(n45), .A2(n44), .A3(n43), .ZN(Y[7]) );
  NAND2_X1 U87 ( .A1(E[8]), .A2(n7), .ZN(n48) );
  NAND2_X1 U88 ( .A1(C[8]), .A2(n95), .ZN(n47) );
  NAND2_X1 U89 ( .A1(A[8]), .A2(n96), .ZN(n46) );
  NAND2_X1 U90 ( .A1(E[9]), .A2(n7), .ZN(n53) );
  NAND2_X1 U91 ( .A1(C[9]), .A2(n95), .ZN(n52) );
  NAND2_X1 U92 ( .A1(A[9]), .A2(n96), .ZN(n51) );
  NAND2_X1 U93 ( .A1(E[10]), .A2(n7), .ZN(n58) );
  NAND2_X1 U94 ( .A1(C[10]), .A2(n95), .ZN(n57) );
  NAND2_X1 U95 ( .A1(A[10]), .A2(n96), .ZN(n56) );
  NAND2_X1 U96 ( .A1(E[11]), .A2(n7), .ZN(n63) );
  NAND2_X1 U97 ( .A1(C[11]), .A2(n95), .ZN(n62) );
  NAND2_X1 U98 ( .A1(A[11]), .A2(n96), .ZN(n61) );
  NAND2_X1 U99 ( .A1(E[12]), .A2(n7), .ZN(n68) );
  NAND2_X1 U100 ( .A1(C[12]), .A2(n95), .ZN(n67) );
  NAND2_X1 U101 ( .A1(A[12]), .A2(n96), .ZN(n66) );
  NAND2_X1 U102 ( .A1(E[13]), .A2(n7), .ZN(n73) );
  NAND2_X1 U103 ( .A1(C[13]), .A2(n95), .ZN(n72) );
  NAND2_X1 U104 ( .A1(A[13]), .A2(n96), .ZN(n71) );
  NAND2_X1 U105 ( .A1(E[14]), .A2(n7), .ZN(n77) );
  NAND2_X1 U106 ( .A1(C[14]), .A2(n95), .ZN(n76) );
  NAND2_X1 U107 ( .A1(A[14]), .A2(n96), .ZN(n75) );
  NAND2_X1 U108 ( .A1(E[15]), .A2(n7), .ZN(n81) );
  NAND2_X1 U109 ( .A1(C[15]), .A2(n95), .ZN(n80) );
  NAND2_X1 U110 ( .A1(A[15]), .A2(n96), .ZN(n79) );
  NAND2_X1 U111 ( .A1(E[16]), .A2(n7), .ZN(n86) );
  NAND2_X1 U112 ( .A1(C[16]), .A2(n95), .ZN(n85) );
  NAND2_X1 U113 ( .A1(A[16]), .A2(n96), .ZN(n84) );
  NAND2_X1 U114 ( .A1(E[17]), .A2(n7), .ZN(n90) );
  NAND2_X1 U115 ( .A1(C[17]), .A2(n95), .ZN(n89) );
  NAND2_X1 U116 ( .A1(A[17]), .A2(n96), .ZN(n88) );
  NAND2_X1 U117 ( .A1(E[18]), .A2(n7), .ZN(n98) );
  NAND3_X1 U118 ( .A1(n99), .A2(n98), .A3(n97), .ZN(Y[18]) );
endmodule


module MUX51_GEN_N19_6 ( A, B, C, D, E, SEL, Y );
  input [18:0] A;
  input [18:0] B;
  input [18:0] C;
  input [18:0] D;
  input [18:0] E;
  input [2:0] SEL;
  output [18:0] Y;
  wire   n1, n2, n3, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104;

  NAND2_X1 U46 ( .A1(n104), .A2(n103), .ZN(Y[9]) );
  NAND2_X1 U47 ( .A1(n97), .A2(n96), .ZN(Y[8]) );
  NAND2_X1 U48 ( .A1(n95), .A2(n94), .ZN(Y[7]) );
  NAND2_X1 U49 ( .A1(n93), .A2(n92), .ZN(Y[6]) );
  NAND2_X1 U50 ( .A1(n91), .A2(n90), .ZN(Y[5]) );
  NAND2_X1 U51 ( .A1(n89), .A2(n88), .ZN(Y[4]) );
  NAND2_X1 U52 ( .A1(n87), .A2(n86), .ZN(Y[3]) );
  NAND2_X1 U53 ( .A1(n85), .A2(n84), .ZN(Y[2]) );
  NAND2_X1 U54 ( .A1(n83), .A2(n82), .ZN(Y[1]) );
  NAND2_X1 U55 ( .A1(n81), .A2(n80), .ZN(Y[18]) );
  NAND2_X1 U56 ( .A1(n79), .A2(n78), .ZN(Y[17]) );
  NAND2_X1 U57 ( .A1(n77), .A2(n76), .ZN(Y[16]) );
  NAND2_X1 U58 ( .A1(n75), .A2(n74), .ZN(Y[15]) );
  NAND2_X1 U59 ( .A1(n73), .A2(n72), .ZN(Y[14]) );
  NAND2_X1 U60 ( .A1(n71), .A2(n70), .ZN(Y[13]) );
  NAND2_X1 U61 ( .A1(n69), .A2(n68), .ZN(Y[12]) );
  NAND2_X1 U62 ( .A1(n67), .A2(n66), .ZN(Y[11]) );
  NAND2_X1 U63 ( .A1(n65), .A2(n64), .ZN(Y[10]) );
  NAND2_X1 U64 ( .A1(n63), .A2(n62), .ZN(Y[0]) );
  AOI222_X4 U1 ( .A1(E[18]), .A2(n59), .B1(B[18]), .B2(n57), .C1(D[18]), .C2(
        n55), .ZN(n80) );
  AOI222_X1 U2 ( .A1(E[17]), .A2(n59), .B1(B[17]), .B2(n101), .C1(D[17]), .C2(
        n100), .ZN(n78) );
  AOI222_X4 U3 ( .A1(E[14]), .A2(n59), .B1(B[14]), .B2(n101), .C1(D[14]), .C2(
        n100), .ZN(n72) );
  AOI222_X4 U4 ( .A1(E[16]), .A2(n59), .B1(B[16]), .B2(n58), .C1(D[16]), .C2(
        n56), .ZN(n76) );
  AOI222_X4 U5 ( .A1(E[13]), .A2(n59), .B1(B[13]), .B2(n58), .C1(D[13]), .C2(
        n56), .ZN(n70) );
  AOI222_X4 U6 ( .A1(E[12]), .A2(n59), .B1(B[12]), .B2(n57), .C1(D[12]), .C2(
        n55), .ZN(n68) );
  AOI222_X4 U7 ( .A1(E[9]), .A2(n59), .B1(B[9]), .B2(n57), .C1(D[9]), .C2(n55), 
        .ZN(n103) );
  AOI222_X1 U8 ( .A1(E[7]), .A2(n59), .B1(B[7]), .B2(n58), .C1(D[7]), .C2(n56), 
        .ZN(n94) );
  CLKBUF_X1 U9 ( .A(n98), .Z(n52) );
  CLKBUF_X1 U10 ( .A(n98), .Z(n51) );
  CLKBUF_X1 U11 ( .A(n98), .Z(n53) );
  CLKBUF_X1 U12 ( .A(n98), .Z(n49) );
  CLKBUF_X1 U13 ( .A(n98), .Z(n3) );
  CLKBUF_X1 U14 ( .A(n98), .Z(n54) );
  BUF_X1 U15 ( .A(n98), .Z(n50) );
  BUF_X1 U16 ( .A(n102), .Z(n59) );
  NOR4_X1 U17 ( .A1(n56), .A2(n58), .A3(n2), .A4(n50), .ZN(n102) );
  AND3_X1 U18 ( .A1(SEL[1]), .A2(n61), .A3(SEL[2]), .ZN(n57) );
  AND3_X1 U19 ( .A1(SEL[1]), .A2(n61), .A3(SEL[2]), .ZN(n101) );
  AND3_X1 U20 ( .A1(SEL[1]), .A2(n61), .A3(SEL[2]), .ZN(n58) );
  INV_X1 U21 ( .A(SEL[1]), .ZN(n60) );
  AND3_X1 U22 ( .A1(SEL[2]), .A2(n60), .A3(SEL[0]), .ZN(n1) );
  AND3_X1 U23 ( .A1(SEL[2]), .A2(n60), .A3(SEL[0]), .ZN(n99) );
  AND3_X1 U24 ( .A1(SEL[2]), .A2(n60), .A3(SEL[0]), .ZN(n2) );
  AND3_X1 U25 ( .A1(n61), .A2(n60), .A3(SEL[2]), .ZN(n55) );
  AND3_X1 U26 ( .A1(n61), .A2(n60), .A3(SEL[2]), .ZN(n100) );
  AND3_X1 U27 ( .A1(n61), .A2(n60), .A3(SEL[2]), .ZN(n56) );
  INV_X1 U28 ( .A(SEL[0]), .ZN(n61) );
  AND3_X1 U29 ( .A1(SEL[2]), .A2(SEL[1]), .A3(SEL[0]), .ZN(n98) );
  AOI22_X1 U30 ( .A1(C[5]), .A2(n99), .B1(A[5]), .B2(n54), .ZN(n91) );
  AOI222_X1 U31 ( .A1(E[5]), .A2(n59), .B1(B[5]), .B2(n101), .C1(D[5]), .C2(
        n100), .ZN(n90) );
  AOI22_X1 U32 ( .A1(C[3]), .A2(n1), .B1(A[3]), .B2(n49), .ZN(n87) );
  AOI222_X1 U33 ( .A1(E[3]), .A2(n59), .B1(B[3]), .B2(n57), .C1(D[3]), .C2(n55), .ZN(n86) );
  AOI22_X1 U34 ( .A1(C[4]), .A2(n2), .B1(A[4]), .B2(n53), .ZN(n89) );
  AOI222_X1 U35 ( .A1(E[4]), .A2(n59), .B1(B[4]), .B2(n58), .C1(D[4]), .C2(n56), .ZN(n88) );
  AOI22_X1 U36 ( .A1(C[2]), .A2(n99), .B1(A[2]), .B2(n53), .ZN(n85) );
  AOI222_X1 U37 ( .A1(E[2]), .A2(n59), .B1(B[2]), .B2(n101), .C1(D[2]), .C2(
        n100), .ZN(n84) );
  AOI222_X1 U38 ( .A1(E[15]), .A2(n59), .B1(B[15]), .B2(n57), .C1(D[15]), .C2(
        n55), .ZN(n74) );
  AOI22_X1 U39 ( .A1(C[15]), .A2(n1), .B1(A[15]), .B2(n52), .ZN(n75) );
  AOI22_X1 U40 ( .A1(C[16]), .A2(n2), .B1(A[16]), .B2(n49), .ZN(n77) );
  AOI22_X1 U41 ( .A1(C[17]), .A2(n99), .B1(A[17]), .B2(n50), .ZN(n79) );
  AOI22_X1 U42 ( .A1(C[9]), .A2(n1), .B1(A[9]), .B2(n51), .ZN(n104) );
  AOI222_X1 U43 ( .A1(E[10]), .A2(n59), .B1(B[10]), .B2(n101), .C1(D[10]), 
        .C2(n100), .ZN(n64) );
  AOI22_X1 U44 ( .A1(C[10]), .A2(n99), .B1(A[10]), .B2(n52), .ZN(n65) );
  AOI222_X1 U45 ( .A1(E[11]), .A2(n59), .B1(B[11]), .B2(n101), .C1(D[11]), 
        .C2(n100), .ZN(n66) );
  AOI22_X1 U65 ( .A1(C[11]), .A2(n99), .B1(A[11]), .B2(n53), .ZN(n67) );
  AOI22_X1 U66 ( .A1(C[12]), .A2(n1), .B1(A[12]), .B2(n54), .ZN(n69) );
  AOI22_X1 U67 ( .A1(C[13]), .A2(n2), .B1(A[13]), .B2(n3), .ZN(n71) );
  AOI22_X1 U68 ( .A1(C[14]), .A2(n99), .B1(A[14]), .B2(n3), .ZN(n73) );
  AOI222_X1 U69 ( .A1(E[8]), .A2(n59), .B1(B[8]), .B2(n101), .C1(D[8]), .C2(
        n100), .ZN(n96) );
  AOI22_X1 U70 ( .A1(C[8]), .A2(n99), .B1(A[8]), .B2(n50), .ZN(n97) );
  AOI22_X1 U71 ( .A1(C[7]), .A2(n2), .B1(A[7]), .B2(n49), .ZN(n95) );
  AOI222_X1 U72 ( .A1(E[6]), .A2(n59), .B1(B[6]), .B2(n57), .C1(D[6]), .C2(n55), .ZN(n92) );
  AOI22_X1 U73 ( .A1(C[6]), .A2(n1), .B1(A[6]), .B2(n3), .ZN(n93) );
  AOI22_X1 U74 ( .A1(C[18]), .A2(n1), .B1(A[18]), .B2(n51), .ZN(n81) );
  AOI22_X1 U75 ( .A1(C[0]), .A2(n1), .B1(A[0]), .B2(n51), .ZN(n63) );
  AOI222_X1 U76 ( .A1(E[0]), .A2(n59), .B1(B[0]), .B2(n57), .C1(D[0]), .C2(n55), .ZN(n62) );
  AOI22_X1 U77 ( .A1(C[1]), .A2(n2), .B1(A[1]), .B2(n52), .ZN(n83) );
  AOI222_X1 U78 ( .A1(E[1]), .A2(n59), .B1(B[1]), .B2(n58), .C1(D[1]), .C2(n56), .ZN(n82) );
endmodule


module MUX51_GEN_N19_5 ( A, B, C, D, E, SEL, Y );
  input [18:0] A;
  input [18:0] B;
  input [18:0] C;
  input [18:0] D;
  input [18:0] E;
  input [2:0] SEL;
  output [18:0] Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93;

  NAND2_X2 U1 ( .A1(n21), .A2(n19), .ZN(n1) );
  INV_X4 U2 ( .A(n21), .ZN(n89) );
  AOI22_X1 U3 ( .A1(C[0]), .A2(n15), .B1(A[0]), .B2(n87), .ZN(n24) );
  INV_X1 U4 ( .A(n17), .ZN(n87) );
  INV_X1 U5 ( .A(SEL[0]), .ZN(n18) );
  CLKBUF_X1 U6 ( .A(n90), .Z(n2) );
  AOI22_X2 U7 ( .A1(n90), .A2(E[0]), .B1(B[0]), .B2(n89), .ZN(n22) );
  INV_X2 U8 ( .A(n18), .ZN(n3) );
  NAND3_X1 U9 ( .A1(n22), .A2(n23), .A3(n24), .ZN(Y[0]) );
  NAND2_X2 U10 ( .A1(n3), .A2(n11), .ZN(n17) );
  NAND2_X2 U11 ( .A1(n18), .A2(n11), .ZN(n21) );
  NAND3_X2 U12 ( .A1(n26), .A2(n27), .A3(n28), .ZN(Y[1]) );
  INV_X1 U13 ( .A(n17), .ZN(n4) );
  INV_X2 U14 ( .A(n19), .ZN(n88) );
  AOI22_X1 U15 ( .A1(C[2]), .A2(n65), .B1(A[2]), .B2(n87), .ZN(n32) );
  AOI22_X4 U16 ( .A1(n9), .A2(E[1]), .B1(B[1]), .B2(n89), .ZN(n26) );
  CLKBUF_X1 U17 ( .A(n2), .Z(n5) );
  NOR2_X2 U18 ( .A1(n20), .A2(n1), .ZN(n9) );
  AOI22_X2 U19 ( .A1(C[1]), .A2(n10), .B1(A[1]), .B2(n87), .ZN(n28) );
  INV_X1 U20 ( .A(n10), .ZN(n6) );
  AND3_X4 U21 ( .A1(n3), .A2(n16), .A3(SEL[2]), .ZN(n10) );
  AND2_X2 U22 ( .A1(SEL[1]), .A2(SEL[2]), .ZN(n11) );
  NAND2_X2 U23 ( .A1(n6), .A2(n17), .ZN(n20) );
  INV_X1 U24 ( .A(n5), .ZN(n7) );
  INV_X1 U25 ( .A(n7), .ZN(n8) );
  INV_X1 U26 ( .A(n12), .ZN(n15) );
  INV_X1 U27 ( .A(n13), .ZN(n33) );
  INV_X1 U28 ( .A(n13), .ZN(n47) );
  INV_X1 U29 ( .A(n13), .ZN(n51) );
  INV_X1 U30 ( .A(n13), .ZN(n65) );
  INV_X1 U31 ( .A(n13), .ZN(n79) );
  INV_X1 U32 ( .A(n13), .ZN(n83) );
  INV_X1 U33 ( .A(n14), .ZN(n25) );
  INV_X1 U34 ( .A(n14), .ZN(n29) );
  INV_X1 U35 ( .A(n14), .ZN(n43) );
  INV_X1 U36 ( .A(n14), .ZN(n58) );
  INV_X1 U37 ( .A(n14), .ZN(n75) );
  INV_X1 U38 ( .A(n10), .ZN(n12) );
  INV_X1 U39 ( .A(n10), .ZN(n13) );
  INV_X1 U40 ( .A(n10), .ZN(n14) );
  NOR2_X1 U41 ( .A1(n20), .A2(n1), .ZN(n90) );
  AOI22_X1 U42 ( .A1(C[17]), .A2(n75), .B1(A[17]), .B2(n4), .ZN(n86) );
  AOI22_X1 U43 ( .A1(E[17]), .A2(n8), .B1(B[17]), .B2(n89), .ZN(n84) );
  AOI22_X1 U44 ( .A1(C[18]), .A2(n75), .B1(A[18]), .B2(n4), .ZN(n93) );
  AOI22_X1 U45 ( .A1(E[18]), .A2(n8), .B1(B[18]), .B2(n89), .ZN(n91) );
  AOI22_X1 U46 ( .A1(n90), .A2(E[2]), .B1(B[2]), .B2(n89), .ZN(n30) );
  AOI22_X1 U47 ( .A1(C[3]), .A2(n51), .B1(A[3]), .B2(n4), .ZN(n36) );
  AOI22_X1 U48 ( .A1(E[3]), .A2(n2), .B1(B[3]), .B2(n89), .ZN(n34) );
  AOI22_X1 U49 ( .A1(C[4]), .A2(n47), .B1(A[4]), .B2(n4), .ZN(n39) );
  AOI22_X1 U50 ( .A1(E[4]), .A2(n5), .B1(B[4]), .B2(n89), .ZN(n37) );
  AOI22_X1 U51 ( .A1(C[5]), .A2(n33), .B1(A[5]), .B2(n4), .ZN(n42) );
  AOI22_X1 U52 ( .A1(E[5]), .A2(n5), .B1(B[5]), .B2(n89), .ZN(n40) );
  AOI22_X1 U53 ( .A1(C[6]), .A2(n33), .B1(A[6]), .B2(n4), .ZN(n46) );
  AOI22_X1 U54 ( .A1(E[6]), .A2(n5), .B1(B[6]), .B2(n89), .ZN(n44) );
  AOI22_X1 U55 ( .A1(C[7]), .A2(n47), .B1(A[7]), .B2(n4), .ZN(n50) );
  AOI22_X1 U56 ( .A1(E[7]), .A2(n5), .B1(B[7]), .B2(n89), .ZN(n48) );
  AOI22_X1 U57 ( .A1(C[8]), .A2(n51), .B1(A[8]), .B2(n4), .ZN(n54) );
  AOI22_X1 U58 ( .A1(E[8]), .A2(n8), .B1(B[8]), .B2(n89), .ZN(n52) );
  AOI22_X1 U59 ( .A1(C[9]), .A2(n65), .B1(A[9]), .B2(n4), .ZN(n57) );
  AOI22_X1 U60 ( .A1(E[9]), .A2(n8), .B1(B[9]), .B2(n89), .ZN(n55) );
  AOI22_X1 U61 ( .A1(C[10]), .A2(n79), .B1(A[10]), .B2(n4), .ZN(n61) );
  AOI22_X1 U62 ( .A1(E[10]), .A2(n8), .B1(B[10]), .B2(n89), .ZN(n59) );
  AOI22_X1 U63 ( .A1(C[11]), .A2(n83), .B1(A[11]), .B2(n4), .ZN(n64) );
  AOI22_X1 U64 ( .A1(E[11]), .A2(n8), .B1(B[11]), .B2(n89), .ZN(n62) );
  AOI22_X1 U65 ( .A1(C[12]), .A2(n25), .B1(A[12]), .B2(n4), .ZN(n68) );
  AOI22_X1 U66 ( .A1(E[12]), .A2(n8), .B1(B[12]), .B2(n89), .ZN(n66) );
  AOI22_X1 U67 ( .A1(C[13]), .A2(n29), .B1(A[13]), .B2(n4), .ZN(n71) );
  AOI22_X1 U68 ( .A1(E[13]), .A2(n8), .B1(B[13]), .B2(n89), .ZN(n69) );
  AOI22_X1 U69 ( .A1(C[14]), .A2(n43), .B1(A[14]), .B2(n4), .ZN(n74) );
  AOI22_X1 U70 ( .A1(E[14]), .A2(n8), .B1(B[14]), .B2(n89), .ZN(n72) );
  AOI22_X1 U71 ( .A1(C[15]), .A2(n58), .B1(A[15]), .B2(n4), .ZN(n78) );
  AOI22_X1 U72 ( .A1(E[15]), .A2(n8), .B1(B[15]), .B2(n89), .ZN(n76) );
  AOI22_X1 U73 ( .A1(C[16]), .A2(n75), .B1(A[16]), .B2(n4), .ZN(n82) );
  AOI22_X1 U74 ( .A1(E[16]), .A2(n8), .B1(B[16]), .B2(n89), .ZN(n80) );
  INV_X1 U75 ( .A(SEL[1]), .ZN(n16) );
  NAND3_X1 U76 ( .A1(n16), .A2(n18), .A3(SEL[2]), .ZN(n19) );
  NAND2_X1 U77 ( .A1(D[0]), .A2(n88), .ZN(n23) );
  NAND2_X1 U78 ( .A1(D[1]), .A2(n88), .ZN(n27) );
  NAND2_X1 U79 ( .A1(D[2]), .A2(n88), .ZN(n31) );
  NAND3_X1 U80 ( .A1(n32), .A2(n31), .A3(n30), .ZN(Y[2]) );
  NAND2_X1 U81 ( .A1(D[3]), .A2(n88), .ZN(n35) );
  NAND3_X1 U82 ( .A1(n36), .A2(n35), .A3(n34), .ZN(Y[3]) );
  NAND2_X1 U83 ( .A1(D[4]), .A2(n88), .ZN(n38) );
  NAND3_X1 U84 ( .A1(n39), .A2(n38), .A3(n37), .ZN(Y[4]) );
  NAND2_X1 U85 ( .A1(D[5]), .A2(n88), .ZN(n41) );
  NAND3_X1 U86 ( .A1(n42), .A2(n41), .A3(n40), .ZN(Y[5]) );
  NAND2_X1 U87 ( .A1(D[6]), .A2(n88), .ZN(n45) );
  NAND3_X1 U88 ( .A1(n46), .A2(n45), .A3(n44), .ZN(Y[6]) );
  NAND2_X1 U89 ( .A1(D[7]), .A2(n88), .ZN(n49) );
  NAND3_X1 U90 ( .A1(n50), .A2(n49), .A3(n48), .ZN(Y[7]) );
  NAND2_X1 U91 ( .A1(D[8]), .A2(n88), .ZN(n53) );
  NAND3_X1 U92 ( .A1(n54), .A2(n53), .A3(n52), .ZN(Y[8]) );
  NAND2_X1 U93 ( .A1(D[9]), .A2(n88), .ZN(n56) );
  NAND3_X1 U94 ( .A1(n57), .A2(n56), .A3(n55), .ZN(Y[9]) );
  NAND2_X1 U95 ( .A1(D[10]), .A2(n88), .ZN(n60) );
  NAND3_X1 U96 ( .A1(n61), .A2(n60), .A3(n59), .ZN(Y[10]) );
  NAND2_X1 U97 ( .A1(D[11]), .A2(n88), .ZN(n63) );
  NAND3_X1 U98 ( .A1(n64), .A2(n63), .A3(n62), .ZN(Y[11]) );
  NAND2_X1 U99 ( .A1(D[12]), .A2(n88), .ZN(n67) );
  NAND3_X1 U100 ( .A1(n68), .A2(n67), .A3(n66), .ZN(Y[12]) );
  NAND2_X1 U101 ( .A1(D[13]), .A2(n88), .ZN(n70) );
  NAND3_X1 U102 ( .A1(n71), .A2(n70), .A3(n69), .ZN(Y[13]) );
  NAND2_X1 U103 ( .A1(D[14]), .A2(n88), .ZN(n73) );
  NAND3_X1 U104 ( .A1(n74), .A2(n73), .A3(n72), .ZN(Y[14]) );
  NAND2_X1 U105 ( .A1(D[15]), .A2(n88), .ZN(n77) );
  NAND3_X1 U106 ( .A1(n78), .A2(n77), .A3(n76), .ZN(Y[15]) );
  NAND2_X1 U107 ( .A1(D[16]), .A2(n88), .ZN(n81) );
  NAND3_X1 U108 ( .A1(n82), .A2(n81), .A3(n80), .ZN(Y[16]) );
  NAND2_X1 U109 ( .A1(D[17]), .A2(n88), .ZN(n85) );
  NAND3_X1 U110 ( .A1(n86), .A2(n85), .A3(n84), .ZN(Y[17]) );
  NAND2_X1 U111 ( .A1(D[18]), .A2(n88), .ZN(n92) );
  NAND3_X1 U112 ( .A1(n93), .A2(n92), .A3(n91), .ZN(Y[18]) );
endmodule


module MUX51_GEN_N19_4 ( A, B, C, D, E, SEL, Y );
  input [18:0] A;
  input [18:0] B;
  input [18:0] C;
  input [18:0] D;
  input [18:0] E;
  input [2:0] SEL;
  output [18:0] Y;
  wire   n1, n2, n3, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104;

  NAND2_X1 U46 ( .A1(n104), .A2(n103), .ZN(Y[9]) );
  NAND2_X1 U47 ( .A1(n97), .A2(n96), .ZN(Y[8]) );
  NAND2_X1 U48 ( .A1(n95), .A2(n94), .ZN(Y[7]) );
  NAND2_X1 U50 ( .A1(n91), .A2(n90), .ZN(Y[5]) );
  NAND2_X1 U51 ( .A1(n89), .A2(n88), .ZN(Y[4]) );
  NAND2_X1 U52 ( .A1(n87), .A2(n86), .ZN(Y[3]) );
  NAND2_X1 U53 ( .A1(n85), .A2(n84), .ZN(Y[2]) );
  NAND2_X1 U55 ( .A1(n81), .A2(n80), .ZN(Y[18]) );
  NAND2_X1 U56 ( .A1(n79), .A2(n78), .ZN(Y[17]) );
  NAND2_X1 U57 ( .A1(n77), .A2(n76), .ZN(Y[16]) );
  NAND2_X1 U58 ( .A1(n75), .A2(n74), .ZN(Y[15]) );
  NAND2_X1 U59 ( .A1(n73), .A2(n72), .ZN(Y[14]) );
  NAND2_X1 U60 ( .A1(n71), .A2(n70), .ZN(Y[13]) );
  NAND2_X1 U61 ( .A1(n69), .A2(n68), .ZN(Y[12]) );
  NAND2_X1 U62 ( .A1(n67), .A2(n66), .ZN(Y[11]) );
  NAND2_X1 U63 ( .A1(n65), .A2(n64), .ZN(Y[10]) );
  NAND2_X1 U64 ( .A1(n63), .A2(n62), .ZN(Y[0]) );
  NAND2_X1 U1 ( .A1(n93), .A2(n92), .ZN(Y[6]) );
  BUF_X1 U2 ( .A(n102), .Z(n59) );
  NAND2_X1 U3 ( .A1(n83), .A2(n82), .ZN(Y[1]) );
  CLKBUF_X1 U4 ( .A(n98), .Z(n52) );
  CLKBUF_X1 U5 ( .A(n98), .Z(n51) );
  CLKBUF_X1 U6 ( .A(n98), .Z(n53) );
  CLKBUF_X1 U7 ( .A(n98), .Z(n49) );
  CLKBUF_X1 U8 ( .A(n98), .Z(n3) );
  CLKBUF_X1 U9 ( .A(n98), .Z(n54) );
  BUF_X1 U10 ( .A(n98), .Z(n50) );
  NOR4_X1 U11 ( .A1(n56), .A2(n58), .A3(n2), .A4(n50), .ZN(n102) );
  AND3_X1 U12 ( .A1(SEL[1]), .A2(n61), .A3(SEL[2]), .ZN(n101) );
  AND3_X1 U13 ( .A1(SEL[1]), .A2(n61), .A3(SEL[2]), .ZN(n57) );
  AND3_X1 U14 ( .A1(SEL[1]), .A2(n61), .A3(SEL[2]), .ZN(n58) );
  INV_X1 U15 ( .A(SEL[1]), .ZN(n60) );
  AND3_X1 U16 ( .A1(SEL[2]), .A2(n60), .A3(SEL[0]), .ZN(n99) );
  AND3_X1 U17 ( .A1(SEL[2]), .A2(n60), .A3(SEL[0]), .ZN(n1) );
  AND3_X1 U18 ( .A1(SEL[2]), .A2(n60), .A3(SEL[0]), .ZN(n2) );
  AND3_X1 U19 ( .A1(n61), .A2(n60), .A3(SEL[2]), .ZN(n100) );
  AND3_X1 U20 ( .A1(n61), .A2(n60), .A3(SEL[2]), .ZN(n55) );
  AND3_X1 U21 ( .A1(n61), .A2(n60), .A3(SEL[2]), .ZN(n56) );
  INV_X1 U22 ( .A(SEL[0]), .ZN(n61) );
  AND3_X1 U23 ( .A1(SEL[2]), .A2(SEL[1]), .A3(SEL[0]), .ZN(n98) );
  AOI22_X1 U24 ( .A1(C[3]), .A2(n1), .B1(A[3]), .B2(n49), .ZN(n87) );
  AOI222_X1 U25 ( .A1(E[3]), .A2(n59), .B1(B[3]), .B2(n57), .C1(D[3]), .C2(n55), .ZN(n86) );
  AOI22_X1 U26 ( .A1(C[4]), .A2(n2), .B1(A[4]), .B2(n53), .ZN(n89) );
  AOI222_X1 U27 ( .A1(E[4]), .A2(n59), .B1(B[4]), .B2(n58), .C1(D[4]), .C2(n56), .ZN(n88) );
  AOI22_X1 U28 ( .A1(C[5]), .A2(n99), .B1(A[5]), .B2(n54), .ZN(n91) );
  AOI222_X1 U29 ( .A1(E[5]), .A2(n59), .B1(B[5]), .B2(n101), .C1(D[5]), .C2(
        n100), .ZN(n90) );
  AOI22_X1 U30 ( .A1(C[6]), .A2(n1), .B1(A[6]), .B2(n3), .ZN(n93) );
  AOI222_X1 U31 ( .A1(E[6]), .A2(n59), .B1(B[6]), .B2(n57), .C1(D[6]), .C2(n55), .ZN(n92) );
  AOI22_X1 U32 ( .A1(C[7]), .A2(n2), .B1(A[7]), .B2(n49), .ZN(n95) );
  AOI222_X1 U33 ( .A1(E[7]), .A2(n59), .B1(B[7]), .B2(n58), .C1(D[7]), .C2(n56), .ZN(n94) );
  AOI22_X1 U34 ( .A1(C[8]), .A2(n99), .B1(A[8]), .B2(n50), .ZN(n97) );
  AOI222_X1 U35 ( .A1(E[8]), .A2(n59), .B1(B[8]), .B2(n101), .C1(D[8]), .C2(
        n100), .ZN(n96) );
  AOI22_X1 U36 ( .A1(C[9]), .A2(n1), .B1(A[9]), .B2(n51), .ZN(n104) );
  AOI222_X1 U37 ( .A1(E[9]), .A2(n59), .B1(B[9]), .B2(n57), .C1(D[9]), .C2(n55), .ZN(n103) );
  AOI22_X1 U38 ( .A1(C[10]), .A2(n99), .B1(A[10]), .B2(n52), .ZN(n65) );
  AOI222_X1 U39 ( .A1(E[10]), .A2(n59), .B1(B[10]), .B2(n101), .C1(D[10]), 
        .C2(n100), .ZN(n64) );
  AOI22_X1 U40 ( .A1(C[11]), .A2(n99), .B1(A[11]), .B2(n53), .ZN(n67) );
  AOI222_X1 U41 ( .A1(E[11]), .A2(n59), .B1(B[11]), .B2(n101), .C1(D[11]), 
        .C2(n100), .ZN(n66) );
  AOI22_X1 U42 ( .A1(C[12]), .A2(n1), .B1(A[12]), .B2(n54), .ZN(n69) );
  AOI222_X1 U43 ( .A1(E[12]), .A2(n59), .B1(B[12]), .B2(n57), .C1(D[12]), .C2(
        n55), .ZN(n68) );
  AOI22_X1 U44 ( .A1(C[13]), .A2(n2), .B1(A[13]), .B2(n3), .ZN(n71) );
  AOI222_X1 U45 ( .A1(E[13]), .A2(n59), .B1(B[13]), .B2(n58), .C1(D[13]), .C2(
        n56), .ZN(n70) );
  AOI22_X1 U49 ( .A1(C[14]), .A2(n99), .B1(A[14]), .B2(n3), .ZN(n73) );
  AOI222_X1 U54 ( .A1(E[14]), .A2(n59), .B1(B[14]), .B2(n101), .C1(D[14]), 
        .C2(n100), .ZN(n72) );
  AOI22_X1 U65 ( .A1(C[15]), .A2(n1), .B1(A[15]), .B2(n52), .ZN(n75) );
  AOI222_X1 U66 ( .A1(E[15]), .A2(n59), .B1(B[15]), .B2(n57), .C1(D[15]), .C2(
        n55), .ZN(n74) );
  AOI22_X1 U67 ( .A1(C[16]), .A2(n2), .B1(A[16]), .B2(n49), .ZN(n77) );
  AOI222_X1 U68 ( .A1(E[16]), .A2(n59), .B1(B[16]), .B2(n58), .C1(D[16]), .C2(
        n56), .ZN(n76) );
  AOI22_X1 U69 ( .A1(C[2]), .A2(n99), .B1(A[2]), .B2(n53), .ZN(n85) );
  AOI222_X1 U70 ( .A1(E[2]), .A2(n59), .B1(B[2]), .B2(n101), .C1(D[2]), .C2(
        n100), .ZN(n84) );
  AOI22_X1 U71 ( .A1(C[0]), .A2(n1), .B1(A[0]), .B2(n51), .ZN(n63) );
  AOI222_X1 U72 ( .A1(E[0]), .A2(n59), .B1(B[0]), .B2(n57), .C1(D[0]), .C2(n55), .ZN(n62) );
  AOI22_X1 U73 ( .A1(C[1]), .A2(n2), .B1(A[1]), .B2(n52), .ZN(n83) );
  AOI222_X1 U74 ( .A1(E[1]), .A2(n59), .B1(B[1]), .B2(n58), .C1(D[1]), .C2(n56), .ZN(n82) );
  AOI22_X1 U75 ( .A1(C[18]), .A2(n1), .B1(A[18]), .B2(n51), .ZN(n81) );
  AOI222_X1 U76 ( .A1(E[18]), .A2(n59), .B1(B[18]), .B2(n57), .C1(D[18]), .C2(
        n55), .ZN(n80) );
  AOI22_X1 U77 ( .A1(C[17]), .A2(n99), .B1(A[17]), .B2(n50), .ZN(n79) );
  AOI222_X1 U78 ( .A1(E[17]), .A2(n59), .B1(B[17]), .B2(n101), .C1(D[17]), 
        .C2(n100), .ZN(n78) );
endmodule


module MUX51_GEN_N19_3 ( A, B, C, D, E, SEL, Y );
  input [18:0] A;
  input [18:0] B;
  input [18:0] C;
  input [18:0] D;
  input [18:0] E;
  input [2:0] SEL;
  output [18:0] Y;
  wire   n1, n2, n3, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104;

  NAND2_X1 U46 ( .A1(n104), .A2(n103), .ZN(Y[9]) );
  NAND2_X1 U47 ( .A1(n97), .A2(n96), .ZN(Y[8]) );
  NAND2_X1 U48 ( .A1(n95), .A2(n94), .ZN(Y[7]) );
  NAND2_X1 U49 ( .A1(n93), .A2(n92), .ZN(Y[6]) );
  NAND2_X1 U50 ( .A1(n91), .A2(n90), .ZN(Y[5]) );
  NAND2_X1 U51 ( .A1(n89), .A2(n88), .ZN(Y[4]) );
  NAND2_X1 U52 ( .A1(n87), .A2(n86), .ZN(Y[3]) );
  NAND2_X1 U53 ( .A1(n85), .A2(n84), .ZN(Y[2]) );
  NAND2_X1 U54 ( .A1(n83), .A2(n82), .ZN(Y[1]) );
  NAND2_X1 U55 ( .A1(n81), .A2(n80), .ZN(Y[18]) );
  NAND2_X1 U56 ( .A1(n79), .A2(n78), .ZN(Y[17]) );
  NAND2_X1 U57 ( .A1(n77), .A2(n76), .ZN(Y[16]) );
  NAND2_X1 U58 ( .A1(n75), .A2(n74), .ZN(Y[15]) );
  NAND2_X1 U59 ( .A1(n73), .A2(n72), .ZN(Y[14]) );
  NAND2_X1 U60 ( .A1(n71), .A2(n70), .ZN(Y[13]) );
  NAND2_X1 U61 ( .A1(n69), .A2(n68), .ZN(Y[12]) );
  NAND2_X1 U62 ( .A1(n67), .A2(n66), .ZN(Y[11]) );
  NAND2_X1 U63 ( .A1(n65), .A2(n64), .ZN(Y[10]) );
  NAND2_X1 U64 ( .A1(n63), .A2(n62), .ZN(Y[0]) );
  BUF_X1 U1 ( .A(n98), .Z(n50) );
  BUF_X1 U2 ( .A(n98), .Z(n49) );
  BUF_X1 U3 ( .A(n98), .Z(n51) );
  BUF_X1 U4 ( .A(n98), .Z(n53) );
  BUF_X1 U5 ( .A(n98), .Z(n3) );
  BUF_X1 U6 ( .A(n98), .Z(n52) );
  BUF_X1 U7 ( .A(n102), .Z(n59) );
  NOR4_X1 U8 ( .A1(n56), .A2(n58), .A3(n2), .A4(n50), .ZN(n102) );
  BUF_X1 U9 ( .A(n98), .Z(n54) );
  AND3_X1 U10 ( .A1(SEL[1]), .A2(n61), .A3(SEL[2]), .ZN(n57) );
  AND3_X1 U11 ( .A1(SEL[1]), .A2(n61), .A3(SEL[2]), .ZN(n101) );
  AND3_X1 U12 ( .A1(SEL[1]), .A2(n61), .A3(SEL[2]), .ZN(n58) );
  INV_X1 U13 ( .A(SEL[1]), .ZN(n60) );
  AND3_X1 U14 ( .A1(SEL[2]), .A2(n60), .A3(SEL[0]), .ZN(n1) );
  AND3_X1 U15 ( .A1(SEL[2]), .A2(n60), .A3(SEL[0]), .ZN(n99) );
  AND3_X1 U16 ( .A1(SEL[2]), .A2(n60), .A3(SEL[0]), .ZN(n2) );
  AND3_X1 U17 ( .A1(n61), .A2(n60), .A3(SEL[2]), .ZN(n55) );
  AND3_X1 U18 ( .A1(n61), .A2(n60), .A3(SEL[2]), .ZN(n100) );
  AND3_X1 U19 ( .A1(n61), .A2(n60), .A3(SEL[2]), .ZN(n56) );
  INV_X1 U20 ( .A(SEL[0]), .ZN(n61) );
  AND3_X1 U21 ( .A1(SEL[2]), .A2(SEL[1]), .A3(SEL[0]), .ZN(n98) );
  AOI22_X1 U22 ( .A1(C[3]), .A2(n1), .B1(A[3]), .B2(n49), .ZN(n87) );
  AOI222_X1 U23 ( .A1(E[3]), .A2(n59), .B1(B[3]), .B2(n57), .C1(D[3]), .C2(n55), .ZN(n86) );
  AOI22_X1 U24 ( .A1(C[4]), .A2(n2), .B1(A[4]), .B2(n53), .ZN(n89) );
  AOI222_X1 U25 ( .A1(E[4]), .A2(n59), .B1(B[4]), .B2(n58), .C1(D[4]), .C2(n56), .ZN(n88) );
  AOI22_X1 U26 ( .A1(C[5]), .A2(n99), .B1(A[5]), .B2(n54), .ZN(n91) );
  AOI222_X1 U27 ( .A1(E[5]), .A2(n59), .B1(B[5]), .B2(n101), .C1(D[5]), .C2(
        n100), .ZN(n90) );
  AOI22_X1 U28 ( .A1(C[6]), .A2(n1), .B1(A[6]), .B2(n3), .ZN(n93) );
  AOI222_X1 U29 ( .A1(E[6]), .A2(n59), .B1(B[6]), .B2(n57), .C1(D[6]), .C2(n55), .ZN(n92) );
  AOI22_X1 U30 ( .A1(C[7]), .A2(n2), .B1(A[7]), .B2(n49), .ZN(n95) );
  AOI222_X1 U31 ( .A1(E[7]), .A2(n59), .B1(B[7]), .B2(n58), .C1(D[7]), .C2(n56), .ZN(n94) );
  AOI22_X1 U32 ( .A1(C[8]), .A2(n99), .B1(A[8]), .B2(n50), .ZN(n97) );
  AOI222_X1 U33 ( .A1(E[8]), .A2(n59), .B1(B[8]), .B2(n101), .C1(D[8]), .C2(
        n100), .ZN(n96) );
  AOI22_X1 U34 ( .A1(C[9]), .A2(n1), .B1(A[9]), .B2(n51), .ZN(n104) );
  AOI222_X1 U35 ( .A1(E[9]), .A2(n59), .B1(B[9]), .B2(n57), .C1(D[9]), .C2(n55), .ZN(n103) );
  AOI22_X1 U36 ( .A1(C[10]), .A2(n99), .B1(A[10]), .B2(n52), .ZN(n65) );
  AOI222_X1 U37 ( .A1(E[10]), .A2(n59), .B1(B[10]), .B2(n101), .C1(D[10]), 
        .C2(n100), .ZN(n64) );
  AOI22_X1 U38 ( .A1(C[11]), .A2(n99), .B1(A[11]), .B2(n53), .ZN(n67) );
  AOI222_X1 U39 ( .A1(E[11]), .A2(n59), .B1(B[11]), .B2(n101), .C1(D[11]), 
        .C2(n100), .ZN(n66) );
  AOI22_X1 U40 ( .A1(C[12]), .A2(n1), .B1(A[12]), .B2(n54), .ZN(n69) );
  AOI222_X1 U41 ( .A1(E[12]), .A2(n59), .B1(B[12]), .B2(n57), .C1(D[12]), .C2(
        n55), .ZN(n68) );
  AOI22_X1 U42 ( .A1(C[2]), .A2(n99), .B1(A[2]), .B2(n53), .ZN(n85) );
  AOI222_X1 U43 ( .A1(E[2]), .A2(n59), .B1(B[2]), .B2(n101), .C1(D[2]), .C2(
        n100), .ZN(n84) );
  AOI22_X1 U44 ( .A1(C[0]), .A2(n1), .B1(A[0]), .B2(n51), .ZN(n63) );
  AOI222_X1 U45 ( .A1(E[0]), .A2(n59), .B1(B[0]), .B2(n57), .C1(D[0]), .C2(n55), .ZN(n62) );
  AOI22_X1 U65 ( .A1(C[1]), .A2(n2), .B1(A[1]), .B2(n52), .ZN(n83) );
  AOI222_X1 U66 ( .A1(E[1]), .A2(n59), .B1(B[1]), .B2(n58), .C1(D[1]), .C2(n56), .ZN(n82) );
  AOI22_X1 U67 ( .A1(C[18]), .A2(n1), .B1(A[18]), .B2(n51), .ZN(n81) );
  AOI222_X1 U68 ( .A1(E[18]), .A2(n59), .B1(B[18]), .B2(n57), .C1(D[18]), .C2(
        n55), .ZN(n80) );
  AOI22_X1 U69 ( .A1(C[17]), .A2(n99), .B1(A[17]), .B2(n50), .ZN(n79) );
  AOI222_X1 U70 ( .A1(E[17]), .A2(n59), .B1(B[17]), .B2(n101), .C1(D[17]), 
        .C2(n100), .ZN(n78) );
  AOI22_X1 U71 ( .A1(C[16]), .A2(n2), .B1(A[16]), .B2(n49), .ZN(n77) );
  AOI222_X1 U72 ( .A1(E[16]), .A2(n59), .B1(B[16]), .B2(n58), .C1(D[16]), .C2(
        n56), .ZN(n76) );
  AOI22_X1 U73 ( .A1(C[13]), .A2(n2), .B1(A[13]), .B2(n3), .ZN(n71) );
  AOI222_X1 U74 ( .A1(E[13]), .A2(n59), .B1(B[13]), .B2(n58), .C1(D[13]), .C2(
        n56), .ZN(n70) );
  AOI22_X1 U75 ( .A1(C[14]), .A2(n99), .B1(A[14]), .B2(n3), .ZN(n73) );
  AOI222_X1 U76 ( .A1(E[14]), .A2(n59), .B1(B[14]), .B2(n101), .C1(D[14]), 
        .C2(n100), .ZN(n72) );
  AOI22_X1 U77 ( .A1(C[15]), .A2(n1), .B1(A[15]), .B2(n52), .ZN(n75) );
  AOI222_X1 U78 ( .A1(E[15]), .A2(n59), .B1(B[15]), .B2(n57), .C1(D[15]), .C2(
        n55), .ZN(n74) );
endmodule


module MUX51_GEN_N19_2 ( A, B, C, D, E, SEL, Y );
  input [18:0] A;
  input [18:0] B;
  input [18:0] C;
  input [18:0] D;
  input [18:0] E;
  input [2:0] SEL;
  output [18:0] Y;
  wire   n1, n2, n3, n7, n10, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98;

  NAND2_X1 U46 ( .A1(n98), .A2(n97), .ZN(Y[9]) );
  NAND2_X1 U47 ( .A1(n93), .A2(n92), .ZN(Y[8]) );
  NAND2_X1 U48 ( .A1(n91), .A2(n90), .ZN(Y[7]) );
  NAND2_X1 U49 ( .A1(n89), .A2(n88), .ZN(Y[6]) );
  NAND2_X1 U50 ( .A1(n87), .A2(n86), .ZN(Y[5]) );
  NAND2_X1 U51 ( .A1(n85), .A2(n84), .ZN(Y[4]) );
  NAND2_X1 U52 ( .A1(n83), .A2(n82), .ZN(Y[3]) );
  NAND2_X1 U53 ( .A1(n81), .A2(n80), .ZN(Y[2]) );
  NAND2_X1 U55 ( .A1(n77), .A2(n76), .ZN(Y[18]) );
  NAND2_X1 U56 ( .A1(n75), .A2(n74), .ZN(Y[17]) );
  NAND2_X1 U57 ( .A1(n73), .A2(n72), .ZN(Y[16]) );
  NAND2_X1 U58 ( .A1(n71), .A2(n70), .ZN(Y[15]) );
  NAND2_X1 U59 ( .A1(n69), .A2(n68), .ZN(Y[14]) );
  NAND2_X1 U60 ( .A1(n67), .A2(n66), .ZN(Y[13]) );
  NAND2_X1 U61 ( .A1(n65), .A2(n64), .ZN(Y[12]) );
  NAND2_X1 U62 ( .A1(n63), .A2(n62), .ZN(Y[11]) );
  NAND2_X1 U63 ( .A1(n61), .A2(n60), .ZN(Y[10]) );
  NAND2_X1 U64 ( .A1(n59), .A2(n58), .ZN(Y[0]) );
  INV_X8 U1 ( .A(n2), .ZN(n96) );
  AND3_X1 U2 ( .A1(SEL[1]), .A2(SEL[2]), .A3(SEL[0]), .ZN(n1) );
  NAND2_X2 U3 ( .A1(n78), .A2(n79), .ZN(Y[1]) );
  AND3_X2 U4 ( .A1(SEL[2]), .A2(n56), .A3(SEL[0]), .ZN(n7) );
  INV_X2 U5 ( .A(SEL[0]), .ZN(n57) );
  INV_X2 U6 ( .A(SEL[1]), .ZN(n56) );
  OR4_X4 U7 ( .A1(n53), .A2(n55), .A3(n7), .A4(n1), .ZN(n2) );
  AOI222_X2 U8 ( .A1(E[1]), .A2(n96), .B1(B[1]), .B2(n55), .C1(D[1]), .C2(n53), 
        .ZN(n78) );
  AND3_X2 U9 ( .A1(SEL[1]), .A2(n57), .A3(SEL[2]), .ZN(n55) );
  AND3_X2 U10 ( .A1(n57), .A2(n56), .A3(SEL[2]), .ZN(n53) );
  CLKBUF_X1 U11 ( .A(n1), .Z(n51) );
  CLKBUF_X1 U12 ( .A(n1), .Z(n50) );
  CLKBUF_X1 U13 ( .A(n1), .Z(n10) );
  CLKBUF_X1 U14 ( .A(n1), .Z(n49) );
  AND3_X1 U15 ( .A1(SEL[2]), .A2(n56), .A3(SEL[0]), .ZN(n3) );
  AND3_X1 U16 ( .A1(SEL[2]), .A2(n56), .A3(SEL[0]), .ZN(n94) );
  AND3_X1 U17 ( .A1(n57), .A2(n56), .A3(SEL[2]), .ZN(n52) );
  AND3_X1 U18 ( .A1(n57), .A2(n56), .A3(SEL[2]), .ZN(n95) );
  AOI22_X1 U19 ( .A1(C[17]), .A2(n94), .B1(A[17]), .B2(n10), .ZN(n75) );
  AOI222_X1 U20 ( .A1(E[17]), .A2(n96), .B1(B[17]), .B2(n54), .C1(D[17]), .C2(
        n95), .ZN(n74) );
  AOI22_X1 U21 ( .A1(C[4]), .A2(n7), .B1(A[4]), .B2(n51), .ZN(n85) );
  AOI222_X1 U22 ( .A1(E[4]), .A2(n96), .B1(B[4]), .B2(n55), .C1(D[4]), .C2(n53), .ZN(n84) );
  AOI22_X1 U23 ( .A1(C[3]), .A2(n3), .B1(A[3]), .B2(n10), .ZN(n83) );
  AOI222_X1 U24 ( .A1(E[3]), .A2(n96), .B1(B[3]), .B2(n54), .C1(D[3]), .C2(n52), .ZN(n82) );
  AOI22_X1 U25 ( .A1(C[5]), .A2(n94), .B1(A[5]), .B2(n10), .ZN(n87) );
  AOI222_X1 U26 ( .A1(E[5]), .A2(n96), .B1(B[5]), .B2(n54), .C1(D[5]), .C2(n95), .ZN(n86) );
  AOI22_X1 U27 ( .A1(C[6]), .A2(n3), .B1(A[6]), .B2(n10), .ZN(n89) );
  AOI222_X1 U28 ( .A1(E[6]), .A2(n96), .B1(B[6]), .B2(n54), .C1(D[6]), .C2(n52), .ZN(n88) );
  AOI22_X1 U29 ( .A1(C[7]), .A2(n7), .B1(A[7]), .B2(n10), .ZN(n91) );
  AOI222_X1 U30 ( .A1(E[7]), .A2(n96), .B1(B[7]), .B2(n55), .C1(D[7]), .C2(n53), .ZN(n90) );
  AOI22_X1 U31 ( .A1(C[8]), .A2(n94), .B1(A[8]), .B2(n10), .ZN(n93) );
  AOI222_X1 U32 ( .A1(E[8]), .A2(n96), .B1(B[8]), .B2(n54), .C1(D[8]), .C2(n95), .ZN(n92) );
  AOI22_X1 U33 ( .A1(C[9]), .A2(n3), .B1(A[9]), .B2(n49), .ZN(n98) );
  AOI222_X1 U34 ( .A1(E[9]), .A2(n96), .B1(B[9]), .B2(n54), .C1(D[9]), .C2(n52), .ZN(n97) );
  AOI22_X1 U35 ( .A1(C[10]), .A2(n94), .B1(A[10]), .B2(n50), .ZN(n61) );
  AOI222_X1 U36 ( .A1(E[10]), .A2(n96), .B1(B[10]), .B2(n54), .C1(D[10]), .C2(
        n95), .ZN(n60) );
  AOI22_X1 U37 ( .A1(C[11]), .A2(n94), .B1(A[11]), .B2(n51), .ZN(n63) );
  AOI222_X1 U38 ( .A1(E[11]), .A2(n96), .B1(B[11]), .B2(n54), .C1(D[11]), .C2(
        n95), .ZN(n62) );
  AOI22_X1 U39 ( .A1(C[12]), .A2(n3), .B1(A[12]), .B2(n10), .ZN(n65) );
  AOI222_X1 U40 ( .A1(E[12]), .A2(n96), .B1(B[12]), .B2(n54), .C1(D[12]), .C2(
        n52), .ZN(n64) );
  AOI22_X1 U41 ( .A1(C[13]), .A2(n7), .B1(A[13]), .B2(n10), .ZN(n67) );
  AOI222_X1 U42 ( .A1(E[13]), .A2(n96), .B1(B[13]), .B2(n55), .C1(D[13]), .C2(
        n53), .ZN(n66) );
  AOI22_X1 U43 ( .A1(C[14]), .A2(n94), .B1(A[14]), .B2(n10), .ZN(n69) );
  AOI222_X1 U44 ( .A1(E[14]), .A2(n96), .B1(B[14]), .B2(n54), .C1(D[14]), .C2(
        n95), .ZN(n68) );
  AOI22_X1 U45 ( .A1(C[15]), .A2(n3), .B1(A[15]), .B2(n50), .ZN(n71) );
  AOI222_X1 U54 ( .A1(E[15]), .A2(n96), .B1(B[15]), .B2(n54), .C1(D[15]), .C2(
        n52), .ZN(n70) );
  AOI22_X1 U65 ( .A1(C[16]), .A2(n7), .B1(A[16]), .B2(n10), .ZN(n73) );
  AOI222_X1 U66 ( .A1(E[16]), .A2(n96), .B1(B[16]), .B2(n55), .C1(D[16]), .C2(
        n53), .ZN(n72) );
  AOI22_X1 U67 ( .A1(C[2]), .A2(n94), .B1(A[2]), .B2(n51), .ZN(n81) );
  AOI222_X1 U68 ( .A1(E[2]), .A2(n96), .B1(B[2]), .B2(n54), .C1(D[2]), .C2(n95), .ZN(n80) );
  AOI22_X1 U69 ( .A1(C[0]), .A2(n3), .B1(A[0]), .B2(n49), .ZN(n59) );
  AOI222_X1 U70 ( .A1(E[0]), .A2(n96), .B1(B[0]), .B2(n54), .C1(D[0]), .C2(n52), .ZN(n58) );
  AOI22_X1 U71 ( .A1(C[1]), .A2(n7), .B1(A[1]), .B2(n50), .ZN(n79) );
  AOI22_X1 U72 ( .A1(C[18]), .A2(n3), .B1(A[18]), .B2(n49), .ZN(n77) );
  AOI222_X1 U73 ( .A1(E[18]), .A2(n96), .B1(B[18]), .B2(n54), .C1(D[18]), .C2(
        n52), .ZN(n76) );
  AND3_X1 U74 ( .A1(SEL[1]), .A2(n57), .A3(SEL[2]), .ZN(n54) );
endmodule


module MUX51_GEN_N19_1 ( A, B, C, D, E, SEL, Y );
  input [18:0] A;
  input [18:0] B;
  input [18:0] C;
  input [18:0] D;
  input [18:0] E;
  input [2:0] SEL;
  output [18:0] Y;
  wire   n1, n2, n3, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104;

  NAND2_X1 U46 ( .A1(n104), .A2(n103), .ZN(Y[9]) );
  NAND2_X1 U47 ( .A1(n97), .A2(n96), .ZN(Y[8]) );
  NAND2_X1 U48 ( .A1(n95), .A2(n94), .ZN(Y[7]) );
  NAND2_X1 U49 ( .A1(n93), .A2(n92), .ZN(Y[6]) );
  NAND2_X1 U50 ( .A1(n91), .A2(n90), .ZN(Y[5]) );
  NAND2_X1 U51 ( .A1(n89), .A2(n88), .ZN(Y[4]) );
  NAND2_X1 U52 ( .A1(n87), .A2(n86), .ZN(Y[3]) );
  NAND2_X1 U53 ( .A1(n85), .A2(n84), .ZN(Y[2]) );
  NAND2_X1 U54 ( .A1(n83), .A2(n82), .ZN(Y[1]) );
  NAND2_X1 U55 ( .A1(n81), .A2(n80), .ZN(Y[18]) );
  NAND2_X1 U56 ( .A1(n79), .A2(n78), .ZN(Y[17]) );
  NAND2_X1 U57 ( .A1(n77), .A2(n76), .ZN(Y[16]) );
  NAND2_X1 U58 ( .A1(n75), .A2(n74), .ZN(Y[15]) );
  NAND2_X1 U59 ( .A1(n73), .A2(n72), .ZN(Y[14]) );
  NAND2_X1 U60 ( .A1(n71), .A2(n70), .ZN(Y[13]) );
  NAND2_X1 U61 ( .A1(n69), .A2(n68), .ZN(Y[12]) );
  NAND2_X1 U62 ( .A1(n67), .A2(n66), .ZN(Y[11]) );
  NAND2_X1 U63 ( .A1(n65), .A2(n64), .ZN(Y[10]) );
  NAND2_X1 U64 ( .A1(n63), .A2(n62), .ZN(Y[0]) );
  CLKBUF_X1 U1 ( .A(n98), .Z(n52) );
  CLKBUF_X1 U2 ( .A(n98), .Z(n51) );
  CLKBUF_X1 U3 ( .A(n98), .Z(n53) );
  CLKBUF_X1 U4 ( .A(n98), .Z(n49) );
  CLKBUF_X1 U5 ( .A(n98), .Z(n3) );
  CLKBUF_X1 U6 ( .A(n98), .Z(n54) );
  BUF_X1 U7 ( .A(n98), .Z(n50) );
  BUF_X1 U8 ( .A(n102), .Z(n59) );
  NOR4_X1 U9 ( .A1(n56), .A2(n58), .A3(n2), .A4(n50), .ZN(n102) );
  AND3_X1 U10 ( .A1(SEL[1]), .A2(n61), .A3(SEL[2]), .ZN(n101) );
  AND3_X1 U11 ( .A1(SEL[1]), .A2(n61), .A3(SEL[2]), .ZN(n57) );
  AND3_X1 U12 ( .A1(SEL[1]), .A2(n61), .A3(SEL[2]), .ZN(n58) );
  INV_X1 U13 ( .A(SEL[1]), .ZN(n60) );
  AND3_X1 U14 ( .A1(SEL[2]), .A2(n60), .A3(SEL[0]), .ZN(n99) );
  AND3_X1 U15 ( .A1(SEL[2]), .A2(n60), .A3(SEL[0]), .ZN(n1) );
  AND3_X1 U16 ( .A1(SEL[2]), .A2(n60), .A3(SEL[0]), .ZN(n2) );
  AND3_X1 U17 ( .A1(n61), .A2(n60), .A3(SEL[2]), .ZN(n100) );
  AND3_X1 U18 ( .A1(n61), .A2(n60), .A3(SEL[2]), .ZN(n55) );
  AND3_X1 U19 ( .A1(n61), .A2(n60), .A3(SEL[2]), .ZN(n56) );
  INV_X1 U20 ( .A(SEL[0]), .ZN(n61) );
  AND3_X1 U21 ( .A1(SEL[2]), .A2(SEL[1]), .A3(SEL[0]), .ZN(n98) );
  AOI22_X1 U22 ( .A1(C[1]), .A2(n2), .B1(A[1]), .B2(n52), .ZN(n83) );
  AOI222_X1 U23 ( .A1(E[1]), .A2(n59), .B1(B[1]), .B2(n58), .C1(D[1]), .C2(n56), .ZN(n82) );
  AOI22_X1 U24 ( .A1(C[3]), .A2(n1), .B1(A[3]), .B2(n49), .ZN(n87) );
  AOI222_X1 U25 ( .A1(E[3]), .A2(n59), .B1(B[3]), .B2(n57), .C1(D[3]), .C2(n55), .ZN(n86) );
  AOI22_X1 U26 ( .A1(C[4]), .A2(n2), .B1(A[4]), .B2(n53), .ZN(n89) );
  AOI222_X1 U27 ( .A1(E[4]), .A2(n59), .B1(B[4]), .B2(n58), .C1(D[4]), .C2(n56), .ZN(n88) );
  AOI22_X1 U28 ( .A1(C[7]), .A2(n2), .B1(A[7]), .B2(n49), .ZN(n95) );
  AOI222_X1 U29 ( .A1(E[7]), .A2(n59), .B1(B[7]), .B2(n58), .C1(D[7]), .C2(n56), .ZN(n94) );
  AOI22_X1 U30 ( .A1(C[12]), .A2(n1), .B1(A[12]), .B2(n54), .ZN(n69) );
  AOI222_X1 U31 ( .A1(E[12]), .A2(n59), .B1(B[12]), .B2(n57), .C1(D[12]), .C2(
        n55), .ZN(n68) );
  AOI22_X1 U32 ( .A1(C[6]), .A2(n1), .B1(A[6]), .B2(n3), .ZN(n93) );
  AOI222_X1 U33 ( .A1(E[6]), .A2(n59), .B1(B[6]), .B2(n57), .C1(D[6]), .C2(n55), .ZN(n92) );
  AOI22_X1 U34 ( .A1(C[8]), .A2(n99), .B1(A[8]), .B2(n50), .ZN(n97) );
  AOI222_X1 U35 ( .A1(E[8]), .A2(n59), .B1(B[8]), .B2(n101), .C1(D[8]), .C2(
        n100), .ZN(n96) );
  AOI22_X1 U36 ( .A1(C[13]), .A2(n2), .B1(A[13]), .B2(n3), .ZN(n71) );
  AOI222_X1 U37 ( .A1(E[13]), .A2(n59), .B1(B[13]), .B2(n58), .C1(D[13]), .C2(
        n56), .ZN(n70) );
  AOI22_X1 U38 ( .A1(C[5]), .A2(n99), .B1(A[5]), .B2(n54), .ZN(n91) );
  AOI222_X1 U39 ( .A1(E[5]), .A2(n59), .B1(B[5]), .B2(n101), .C1(D[5]), .C2(
        n100), .ZN(n90) );
  AOI22_X1 U40 ( .A1(C[9]), .A2(n1), .B1(A[9]), .B2(n51), .ZN(n104) );
  AOI222_X1 U41 ( .A1(E[9]), .A2(n59), .B1(B[9]), .B2(n57), .C1(D[9]), .C2(n55), .ZN(n103) );
  AOI22_X1 U42 ( .A1(C[10]), .A2(n99), .B1(A[10]), .B2(n52), .ZN(n65) );
  AOI222_X1 U43 ( .A1(E[10]), .A2(n59), .B1(B[10]), .B2(n101), .C1(D[10]), 
        .C2(n100), .ZN(n64) );
  AOI22_X1 U44 ( .A1(C[11]), .A2(n99), .B1(A[11]), .B2(n53), .ZN(n67) );
  AOI222_X1 U45 ( .A1(E[11]), .A2(n59), .B1(B[11]), .B2(n101), .C1(D[11]), 
        .C2(n100), .ZN(n66) );
  AOI22_X1 U65 ( .A1(C[14]), .A2(n99), .B1(A[14]), .B2(n3), .ZN(n73) );
  AOI222_X1 U66 ( .A1(E[14]), .A2(n59), .B1(B[14]), .B2(n101), .C1(D[14]), 
        .C2(n100), .ZN(n72) );
  AOI22_X1 U67 ( .A1(C[2]), .A2(n99), .B1(A[2]), .B2(n53), .ZN(n85) );
  AOI222_X1 U68 ( .A1(E[2]), .A2(n59), .B1(B[2]), .B2(n101), .C1(D[2]), .C2(
        n100), .ZN(n84) );
  AOI22_X1 U69 ( .A1(C[0]), .A2(n1), .B1(A[0]), .B2(n51), .ZN(n63) );
  AOI222_X1 U70 ( .A1(E[0]), .A2(n59), .B1(B[0]), .B2(n57), .C1(D[0]), .C2(n55), .ZN(n62) );
  AOI22_X1 U71 ( .A1(C[15]), .A2(n1), .B1(A[15]), .B2(n52), .ZN(n75) );
  AOI222_X1 U72 ( .A1(E[15]), .A2(n59), .B1(B[15]), .B2(n57), .C1(D[15]), .C2(
        n55), .ZN(n74) );
  AOI22_X1 U73 ( .A1(C[16]), .A2(n2), .B1(A[16]), .B2(n49), .ZN(n77) );
  AOI222_X1 U74 ( .A1(E[16]), .A2(n59), .B1(B[16]), .B2(n58), .C1(D[16]), .C2(
        n56), .ZN(n76) );
  AOI22_X1 U75 ( .A1(C[18]), .A2(n1), .B1(A[18]), .B2(n51), .ZN(n81) );
  AOI222_X1 U76 ( .A1(E[18]), .A2(n59), .B1(B[18]), .B2(n57), .C1(D[18]), .C2(
        n55), .ZN(n80) );
  AOI22_X1 U77 ( .A1(C[17]), .A2(n99), .B1(A[17]), .B2(n50), .ZN(n79) );
  AOI222_X1 U78 ( .A1(E[17]), .A2(n59), .B1(B[17]), .B2(n101), .C1(D[17]), 
        .C2(n100), .ZN(n78) );
endmodule


module PG_BLOCK_26 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_26 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_26 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_25 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_25 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_25 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_24 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_24 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_24 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_23 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_23 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_23 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_22 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_22 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_22 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_21 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_21 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_21 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_20 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_20 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_20 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_19 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_19 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_19 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_18 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_18 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_18 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_17 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_17 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_17 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_16 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_16 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_16 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_15 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_15 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_15 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_14 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_14 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_14 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_13 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_13 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_13 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_12 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_12 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_12 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_11 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_11 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_11 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_10 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_10 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_10 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_9 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_9 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_9 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_8 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_8 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_8 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_7 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_7 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_7 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_6 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_6 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_6 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_5 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_5 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_5 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_4 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_4 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_4 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_3 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_3 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_3 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_2 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_2 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_2 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module PG_BLOCK_1 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_1 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_1 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module GENERAL_GENERATE_36 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_481 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_241 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_35 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_480 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_240 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_34 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_479 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_239 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_33 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_478 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_238 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_32 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_477 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_237 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_31 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_476 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_236 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_30 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_475 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_235 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_29 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_474 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_234 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_28 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_442 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_218 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_27 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_441 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_217 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_26 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_439 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_216 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_25 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_437 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_215 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_24 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_435 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_214 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_23 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_433 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_213 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_22 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_431 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_212 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_21 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_429 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_211 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_20 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_427 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_210 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_19 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_425 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_209 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_18 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_423 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_208 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_17 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_421 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_207 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_16 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_419 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_206 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_15 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_417 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_205 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_14 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_415 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_204 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_13 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_413 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_203 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_12 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_411 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_202 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_11 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_409 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_201 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_10 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_407 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_200 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_9 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_405 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_199 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_8 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_403 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_198 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_7 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_401 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_197 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_6 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_399 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_196 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_5 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_397 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_195 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_4 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_395 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_194 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_3 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_393 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_193 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_2 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_391 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_192 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module GENERAL_GENERATE_1 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_389 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_191 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module REG_N16_5 ( D, Q, EN, RST, CLK );
  input [15:0] D;
  output [15:0] Q;
  input EN, RST, CLK;
  wire   n1, n2;

  FD_107 FF_0 ( .D(D[0]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[0]) );
  FD_106 FF_1 ( .D(D[1]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[1]) );
  FD_105 FF_2 ( .D(D[2]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[2]) );
  FD_104 FF_3 ( .D(D[3]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[3]) );
  FD_103 FF_4 ( .D(D[4]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[4]) );
  FD_102 FF_5 ( .D(D[5]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[5]) );
  FD_101 FF_6 ( .D(D[6]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[6]) );
  FD_100 FF_7 ( .D(D[7]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[7]) );
  FD_99 FF_8 ( .D(D[8]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[8]) );
  FD_98 FF_9 ( .D(D[9]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[9]) );
  FD_97 FF_10 ( .D(D[10]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[10]) );
  FD_96 FF_11 ( .D(D[11]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[11]) );
  FD_95 FF_12 ( .D(D[12]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[12]) );
  FD_94 FF_13 ( .D(D[13]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[13]) );
  FD_93 FF_14 ( .D(D[14]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[14]) );
  FD_92 FF_15 ( .D(D[15]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[15]) );
  BUF_X1 U1 ( .A(RST), .Z(n1) );
  BUF_X1 U2 ( .A(RST), .Z(n2) );
endmodule


module REG_N16_4 ( D, Q, EN, RST, CLK );
  input [15:0] D;
  output [15:0] Q;
  input EN, RST, CLK;
  wire   n1, n2;

  FD_91 FF_0 ( .D(D[0]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[0]) );
  FD_90 FF_1 ( .D(D[1]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[1]) );
  FD_89 FF_2 ( .D(D[2]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[2]) );
  FD_88 FF_3 ( .D(D[3]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[3]) );
  FD_87 FF_4 ( .D(D[4]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[4]) );
  FD_86 FF_5 ( .D(D[5]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[5]) );
  FD_85 FF_6 ( .D(D[6]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[6]) );
  FD_84 FF_7 ( .D(D[7]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[7]) );
  FD_83 FF_8 ( .D(D[8]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[8]) );
  FD_82 FF_9 ( .D(D[9]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[9]) );
  FD_81 FF_10 ( .D(D[10]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[10]) );
  FD_80 FF_11 ( .D(D[11]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[11]) );
  FD_79 FF_12 ( .D(D[12]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[12]) );
  FD_78 FF_13 ( .D(D[13]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[13]) );
  FD_77 FF_14 ( .D(D[14]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[14]) );
  FD_76 FF_15 ( .D(D[15]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[15]) );
  BUF_X1 U1 ( .A(RST), .Z(n1) );
  BUF_X1 U2 ( .A(RST), .Z(n2) );
endmodule


module REG_N16_3 ( D, Q, EN, RST, CLK );
  input [15:0] D;
  output [15:0] Q;
  input EN, RST, CLK;
  wire   n1, n2;

  FD_48 FF_0 ( .D(D[0]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[0]) );
  FD_47 FF_1 ( .D(D[1]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[1]) );
  FD_46 FF_2 ( .D(D[2]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[2]) );
  FD_45 FF_3 ( .D(D[3]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[3]) );
  FD_44 FF_4 ( .D(D[4]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[4]) );
  FD_43 FF_5 ( .D(D[5]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[5]) );
  FD_42 FF_6 ( .D(D[6]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[6]) );
  FD_41 FF_7 ( .D(D[7]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[7]) );
  FD_40 FF_8 ( .D(D[8]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[8]) );
  FD_39 FF_9 ( .D(D[9]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[9]) );
  FD_38 FF_10 ( .D(D[10]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[10]) );
  FD_37 FF_11 ( .D(D[11]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[11]) );
  FD_36 FF_12 ( .D(D[12]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[12]) );
  FD_35 FF_13 ( .D(D[13]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[13]) );
  FD_34 FF_14 ( .D(D[14]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[14]) );
  FD_33 FF_15 ( .D(D[15]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[15]) );
  BUF_X1 U1 ( .A(RST), .Z(n1) );
  BUF_X1 U2 ( .A(RST), .Z(n2) );
endmodule


module REG_N16_2 ( D, Q, EN, RST, CLK );
  input [15:0] D;
  output [15:0] Q;
  input EN, RST, CLK;
  wire   n1, n2;

  FD_32 FF_0 ( .D(D[0]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[0]) );
  FD_31 FF_1 ( .D(D[1]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[1]) );
  FD_30 FF_2 ( .D(D[2]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[2]) );
  FD_29 FF_3 ( .D(D[3]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[3]) );
  FD_28 FF_4 ( .D(D[4]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[4]) );
  FD_27 FF_5 ( .D(D[5]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[5]) );
  FD_26 FF_6 ( .D(D[6]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[6]) );
  FD_25 FF_7 ( .D(D[7]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[7]) );
  FD_24 FF_8 ( .D(D[8]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[8]) );
  FD_23 FF_9 ( .D(D[9]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[9]) );
  FD_22 FF_10 ( .D(D[10]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[10]) );
  FD_21 FF_11 ( .D(D[11]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[11]) );
  FD_20 FF_12 ( .D(D[12]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[12]) );
  FD_19 FF_13 ( .D(D[13]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[13]) );
  FD_18 FF_14 ( .D(D[14]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[14]) );
  FD_17 FF_15 ( .D(D[15]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[15]) );
  BUF_X1 U1 ( .A(RST), .Z(n1) );
  BUF_X1 U2 ( .A(RST), .Z(n2) );
endmodule


module REG_N16_1 ( D, Q, EN, RST, CLK );
  input [15:0] D;
  output [15:0] Q;
  input EN, RST, CLK;
  wire   n1, n2;

  FD_16 FF_0 ( .D(D[0]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[0]) );
  FD_15 FF_1 ( .D(D[1]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[1]) );
  FD_14 FF_2 ( .D(D[2]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[2]) );
  FD_13 FF_3 ( .D(D[3]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[3]) );
  FD_12 FF_4 ( .D(D[4]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[4]) );
  FD_11 FF_5 ( .D(D[5]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[5]) );
  FD_10 FF_6 ( .D(D[6]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[6]) );
  FD_9 FF_7 ( .D(D[7]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[7]) );
  FD_8 FF_8 ( .D(D[8]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[8]) );
  FD_7 FF_9 ( .D(D[9]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[9]) );
  FD_6 FF_10 ( .D(D[10]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[10]) );
  FD_5 FF_11 ( .D(D[11]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[11]) );
  FD_4 FF_12 ( .D(D[12]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[12]) );
  FD_3 FF_13 ( .D(D[13]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[13]) );
  FD_2 FF_14 ( .D(D[14]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[14]) );
  FD_1 FF_15 ( .D(D[15]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[15]) );
  BUF_X1 U1 ( .A(RST), .Z(n1) );
  BUF_X1 U2 ( .A(RST), .Z(n2) );
endmodule


module REG_N17_1 ( D, Q, EN, RST, CLK );
  input [16:0] D;
  output [16:0] Q;
  input EN, RST, CLK;
  wire   n1, n2;

  FD_65 FF_0 ( .D(D[0]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[0]) );
  FD_64 FF_1 ( .D(D[1]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[1]) );
  FD_63 FF_2 ( .D(D[2]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[2]) );
  FD_62 FF_3 ( .D(D[3]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[3]) );
  FD_61 FF_4 ( .D(D[4]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[4]) );
  FD_60 FF_5 ( .D(D[5]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[5]) );
  FD_59 FF_6 ( .D(D[6]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[6]) );
  FD_58 FF_7 ( .D(D[7]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[7]) );
  FD_57 FF_8 ( .D(D[8]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[8]) );
  FD_56 FF_9 ( .D(D[9]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[9]) );
  FD_55 FF_10 ( .D(D[10]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[10]) );
  FD_54 FF_11 ( .D(D[11]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[11]) );
  FD_53 FF_12 ( .D(D[12]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[12]) );
  FD_52 FF_13 ( .D(D[13]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[13]) );
  FD_51 FF_14 ( .D(D[14]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[14]) );
  FD_50 FF_15 ( .D(D[15]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[15]) );
  FD_49 FF_16 ( .D(D[16]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[16]) );
  BUF_X1 U1 ( .A(RST), .Z(n1) );
  BUF_X1 U2 ( .A(RST), .Z(n2) );
endmodule


module MUX21_GEN_N7_3 ( A, B, SEL, Y );
  input [6:0] A;
  input [6:0] B;
  output [6:0] Y;
  input SEL;
  wire   SB;
  wire   [6:0] Y1;
  wire   [6:0] Y2;

  INV_1_22 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_495 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_494 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_493 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_492 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_491 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_490 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_489 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_488 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_487 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_486 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_485 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_484 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_483 UND1_4 ( .A(A[4]), .B(SEL), .Y(Y1[4]) );
  NAND_GATE_482 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  NAND_GATE_481 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_480 UND1_5 ( .A(A[5]), .B(SEL), .Y(Y1[5]) );
  NAND_GATE_479 UND2_5 ( .A(B[5]), .B(SB), .Y(Y2[5]) );
  NAND_GATE_478 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_477 UND1_6 ( .A(A[6]), .B(SEL), .Y(Y1[6]) );
  NAND_GATE_476 UND2_6 ( .A(B[6]), .B(SB), .Y(Y2[6]) );
  NAND_GATE_475 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
endmodule


module MUX21_GEN_N7_2 ( A, B, SEL, Y );
  input [6:0] A;
  input [6:0] B;
  output [6:0] Y;
  input SEL;
  wire   SB;
  wire   [6:0] Y1;
  wire   [6:0] Y2;

  INV_1_17 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_378 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_377 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_376 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_375 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_374 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_373 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_372 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_371 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_370 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_369 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_368 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_367 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_366 UND1_4 ( .A(A[4]), .B(SEL), .Y(Y1[4]) );
  NAND_GATE_365 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  NAND_GATE_364 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_363 UND1_5 ( .A(A[5]), .B(SEL), .Y(Y1[5]) );
  NAND_GATE_362 UND2_5 ( .A(B[5]), .B(SB), .Y(Y2[5]) );
  NAND_GATE_361 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_360 UND1_6 ( .A(A[6]), .B(SEL), .Y(Y1[6]) );
  NAND_GATE_359 UND2_6 ( .A(B[6]), .B(SB), .Y(Y2[6]) );
  NAND_GATE_358 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
endmodule


module MUX21_GEN_N7_1 ( A, B, SEL, Y );
  input [6:0] A;
  input [6:0] B;
  output [6:0] Y;
  input SEL;
  wire   SB;
  wire   [6:0] Y1;
  wire   [6:0] Y2;

  INV_1_12 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_261 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_260 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_259 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_258 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_257 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_256 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_255 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_254 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_253 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_252 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_251 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_250 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_249 UND1_4 ( .A(A[4]), .B(SEL), .Y(Y1[4]) );
  NAND_GATE_248 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  NAND_GATE_247 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_246 UND1_5 ( .A(A[5]), .B(SEL), .Y(Y1[5]) );
  NAND_GATE_245 UND2_5 ( .A(B[5]), .B(SB), .Y(Y2[5]) );
  NAND_GATE_244 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_243 UND1_6 ( .A(A[6]), .B(SEL), .Y(Y1[6]) );
  NAND_GATE_242 UND2_6 ( .A(B[6]), .B(SB), .Y(Y2[6]) );
  NAND_GATE_241 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
endmodule


module MUX21_GEN_N8_15 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;
  wire   SB;
  wire   [7:0] Y1;
  wire   [7:0] Y2;

  INV_1_30 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_684 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_683 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_682 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_681 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_680 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_679 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_678 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_677 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_676 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_675 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_674 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_673 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_672 UND1_4 ( .A(A[4]), .B(SEL), .Y(Y1[4]) );
  NAND_GATE_671 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  NAND_GATE_670 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_669 UND1_5 ( .A(A[5]), .B(SEL), .Y(Y1[5]) );
  NAND_GATE_668 UND2_5 ( .A(B[5]), .B(SB), .Y(Y2[5]) );
  NAND_GATE_667 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_666 UND1_6 ( .A(A[6]), .B(SEL), .Y(Y1[6]) );
  NAND_GATE_665 UND2_6 ( .A(B[6]), .B(SB), .Y(Y2[6]) );
  NAND_GATE_664 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_663 UND1_7 ( .A(A[7]), .B(SEL), .Y(Y1[7]) );
  NAND_GATE_662 UND2_7 ( .A(B[7]), .B(SB), .Y(Y2[7]) );
  NAND_GATE_661 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
endmodule


module MUX21_GEN_N8_14 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;
  wire   SB;
  wire   [7:0] Y1;
  wire   [7:0] Y2;

  INV_1_29 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_660 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_659 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_658 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_657 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_656 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_655 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_654 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_653 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_652 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_651 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_650 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_649 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_648 UND1_4 ( .A(A[4]), .B(SEL), .Y(Y1[4]) );
  NAND_GATE_647 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  NAND_GATE_646 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_645 UND1_5 ( .A(A[5]), .B(SEL), .Y(Y1[5]) );
  NAND_GATE_644 UND2_5 ( .A(B[5]), .B(SB), .Y(Y2[5]) );
  NAND_GATE_643 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_642 UND1_6 ( .A(A[6]), .B(SEL), .Y(Y1[6]) );
  NAND_GATE_641 UND2_6 ( .A(B[6]), .B(SB), .Y(Y2[6]) );
  NAND_GATE_640 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_639 UND1_7 ( .A(A[7]), .B(SEL), .Y(Y1[7]) );
  NAND_GATE_638 UND2_7 ( .A(B[7]), .B(SB), .Y(Y2[7]) );
  NAND_GATE_637 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
endmodule


module MUX21_GEN_N8_13 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;
  wire   SB;
  wire   [7:0] Y1;
  wire   [7:0] Y2;

  INV_1_28 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_636 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_635 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_634 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_633 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_632 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_631 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_630 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_629 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_628 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_627 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_626 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_625 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_624 UND1_4 ( .A(A[4]), .B(SEL), .Y(Y1[4]) );
  NAND_GATE_623 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  NAND_GATE_622 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_621 UND1_5 ( .A(A[5]), .B(SEL), .Y(Y1[5]) );
  NAND_GATE_620 UND2_5 ( .A(B[5]), .B(SB), .Y(Y2[5]) );
  NAND_GATE_619 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_618 UND1_6 ( .A(A[6]), .B(SEL), .Y(Y1[6]) );
  NAND_GATE_617 UND2_6 ( .A(B[6]), .B(SB), .Y(Y2[6]) );
  NAND_GATE_616 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_615 UND1_7 ( .A(A[7]), .B(SEL), .Y(Y1[7]) );
  NAND_GATE_614 UND2_7 ( .A(B[7]), .B(SB), .Y(Y2[7]) );
  NAND_GATE_613 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
endmodule


module MUX21_GEN_N8_12 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;
  wire   SB;
  wire   [7:0] Y1;
  wire   [7:0] Y2;

  INV_1_26 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_591 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_590 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_589 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_588 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_587 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_586 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_585 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_584 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_583 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_582 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_581 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_580 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_579 UND1_4 ( .A(A[4]), .B(SEL), .Y(Y1[4]) );
  NAND_GATE_578 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  NAND_GATE_577 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_576 UND1_5 ( .A(A[5]), .B(SEL), .Y(Y1[5]) );
  NAND_GATE_575 UND2_5 ( .A(B[5]), .B(SB), .Y(Y2[5]) );
  NAND_GATE_574 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_573 UND1_6 ( .A(A[6]), .B(SEL), .Y(Y1[6]) );
  NAND_GATE_572 UND2_6 ( .A(B[6]), .B(SB), .Y(Y2[6]) );
  NAND_GATE_571 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_570 UND1_7 ( .A(A[7]), .B(SEL), .Y(Y1[7]) );
  NAND_GATE_569 UND2_7 ( .A(B[7]), .B(SB), .Y(Y2[7]) );
  NAND_GATE_568 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
endmodule


module MUX21_GEN_N8_11 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;
  wire   SB;
  wire   [7:0] Y1;
  wire   [7:0] Y2;

  INV_1_25 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_567 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_566 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_565 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_564 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_563 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_562 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_561 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_560 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_559 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_558 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_557 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_556 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_555 UND1_4 ( .A(A[4]), .B(SEL), .Y(Y1[4]) );
  NAND_GATE_554 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  NAND_GATE_553 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_552 UND1_5 ( .A(A[5]), .B(SEL), .Y(Y1[5]) );
  NAND_GATE_551 UND2_5 ( .A(B[5]), .B(SB), .Y(Y2[5]) );
  NAND_GATE_550 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_549 UND1_6 ( .A(A[6]), .B(SEL), .Y(Y1[6]) );
  NAND_GATE_548 UND2_6 ( .A(B[6]), .B(SB), .Y(Y2[6]) );
  NAND_GATE_547 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_546 UND1_7 ( .A(A[7]), .B(SEL), .Y(Y1[7]) );
  NAND_GATE_545 UND2_7 ( .A(B[7]), .B(SB), .Y(Y2[7]) );
  NAND_GATE_544 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
endmodule


module MUX21_GEN_N8_10 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;
  wire   SB;
  wire   [7:0] Y1;
  wire   [7:0] Y2;

  INV_1_24 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_543 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_542 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_541 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_540 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_539 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_538 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_537 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_536 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_535 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_534 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_533 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_532 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_531 UND1_4 ( .A(A[4]), .B(SEL), .Y(Y1[4]) );
  NAND_GATE_530 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  NAND_GATE_529 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_528 UND1_5 ( .A(A[5]), .B(SEL), .Y(Y1[5]) );
  NAND_GATE_527 UND2_5 ( .A(B[5]), .B(SB), .Y(Y2[5]) );
  NAND_GATE_526 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_525 UND1_6 ( .A(A[6]), .B(SEL), .Y(Y1[6]) );
  NAND_GATE_524 UND2_6 ( .A(B[6]), .B(SB), .Y(Y2[6]) );
  NAND_GATE_523 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_522 UND1_7 ( .A(A[7]), .B(SEL), .Y(Y1[7]) );
  NAND_GATE_521 UND2_7 ( .A(B[7]), .B(SB), .Y(Y2[7]) );
  NAND_GATE_520 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
endmodule


module MUX21_GEN_N8_9 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;
  wire   SB;
  wire   [7:0] Y1;
  wire   [7:0] Y2;

  INV_1_23 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_519 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_518 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_517 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_516 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_515 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_514 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_513 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_512 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_511 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_510 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_509 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_508 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_507 UND1_4 ( .A(A[4]), .B(SEL), .Y(Y1[4]) );
  NAND_GATE_506 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  NAND_GATE_505 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_504 UND1_5 ( .A(A[5]), .B(SEL), .Y(Y1[5]) );
  NAND_GATE_503 UND2_5 ( .A(B[5]), .B(SB), .Y(Y2[5]) );
  NAND_GATE_502 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_501 UND1_6 ( .A(A[6]), .B(SEL), .Y(Y1[6]) );
  NAND_GATE_500 UND2_6 ( .A(B[6]), .B(SB), .Y(Y2[6]) );
  NAND_GATE_499 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_498 UND1_7 ( .A(A[7]), .B(SEL), .Y(Y1[7]) );
  NAND_GATE_497 UND2_7 ( .A(B[7]), .B(SB), .Y(Y2[7]) );
  NAND_GATE_496 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
endmodule


module MUX21_GEN_N8_8 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;
  wire   SB;
  wire   [7:0] Y1;
  wire   [7:0] Y2;

  INV_1_21 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_474 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_473 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_472 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_471 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_470 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_469 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_468 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_467 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_466 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_465 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_464 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_463 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_462 UND1_4 ( .A(A[4]), .B(SEL), .Y(Y1[4]) );
  NAND_GATE_461 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  NAND_GATE_460 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_459 UND1_5 ( .A(A[5]), .B(SEL), .Y(Y1[5]) );
  NAND_GATE_458 UND2_5 ( .A(B[5]), .B(SB), .Y(Y2[5]) );
  NAND_GATE_457 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_456 UND1_6 ( .A(A[6]), .B(SEL), .Y(Y1[6]) );
  NAND_GATE_455 UND2_6 ( .A(B[6]), .B(SB), .Y(Y2[6]) );
  NAND_GATE_454 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_453 UND1_7 ( .A(A[7]), .B(SEL), .Y(Y1[7]) );
  NAND_GATE_452 UND2_7 ( .A(B[7]), .B(SB), .Y(Y2[7]) );
  NAND_GATE_451 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
endmodule


module MUX21_GEN_N8_7 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;
  wire   SB;
  wire   [7:0] Y1;
  wire   [7:0] Y2;

  INV_1_20 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_450 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_449 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_448 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_447 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_446 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_445 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_444 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_443 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_442 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_441 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_440 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_439 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_438 UND1_4 ( .A(A[4]), .B(SEL), .Y(Y1[4]) );
  NAND_GATE_437 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  NAND_GATE_436 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_435 UND1_5 ( .A(A[5]), .B(SEL), .Y(Y1[5]) );
  NAND_GATE_434 UND2_5 ( .A(B[5]), .B(SB), .Y(Y2[5]) );
  NAND_GATE_433 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_432 UND1_6 ( .A(A[6]), .B(SEL), .Y(Y1[6]) );
  NAND_GATE_431 UND2_6 ( .A(B[6]), .B(SB), .Y(Y2[6]) );
  NAND_GATE_430 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_429 UND1_7 ( .A(A[7]), .B(SEL), .Y(Y1[7]) );
  NAND_GATE_428 UND2_7 ( .A(B[7]), .B(SB), .Y(Y2[7]) );
  NAND_GATE_427 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
endmodule


module MUX21_GEN_N8_6 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;
  wire   SB;
  wire   [7:0] Y1;
  wire   [7:0] Y2;

  INV_1_19 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_426 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_425 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_424 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_423 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_422 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_421 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_420 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_419 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_418 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_417 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_416 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_415 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_414 UND1_4 ( .A(A[4]), .B(SEL), .Y(Y1[4]) );
  NAND_GATE_413 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  NAND_GATE_412 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_411 UND1_5 ( .A(A[5]), .B(SEL), .Y(Y1[5]) );
  NAND_GATE_410 UND2_5 ( .A(B[5]), .B(SB), .Y(Y2[5]) );
  NAND_GATE_409 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_408 UND1_6 ( .A(A[6]), .B(SEL), .Y(Y1[6]) );
  NAND_GATE_407 UND2_6 ( .A(B[6]), .B(SB), .Y(Y2[6]) );
  NAND_GATE_406 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_405 UND1_7 ( .A(A[7]), .B(SEL), .Y(Y1[7]) );
  NAND_GATE_404 UND2_7 ( .A(B[7]), .B(SB), .Y(Y2[7]) );
  NAND_GATE_403 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
endmodule


module MUX21_GEN_N8_5 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;
  wire   SB;
  wire   [7:0] Y1;
  wire   [7:0] Y2;

  INV_1_18 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_402 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_401 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_400 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_399 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_398 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_397 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_396 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_395 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_394 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_393 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_392 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_391 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_390 UND1_4 ( .A(A[4]), .B(SEL), .Y(Y1[4]) );
  NAND_GATE_389 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  NAND_GATE_388 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_387 UND1_5 ( .A(A[5]), .B(SEL), .Y(Y1[5]) );
  NAND_GATE_386 UND2_5 ( .A(B[5]), .B(SB), .Y(Y2[5]) );
  NAND_GATE_385 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_384 UND1_6 ( .A(A[6]), .B(SEL), .Y(Y1[6]) );
  NAND_GATE_383 UND2_6 ( .A(B[6]), .B(SB), .Y(Y2[6]) );
  NAND_GATE_382 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_381 UND1_7 ( .A(A[7]), .B(SEL), .Y(Y1[7]) );
  NAND_GATE_380 UND2_7 ( .A(B[7]), .B(SB), .Y(Y2[7]) );
  NAND_GATE_379 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
endmodule


module MUX21_GEN_N8_4 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;
  wire   SB;
  wire   [7:0] Y1;
  wire   [7:0] Y2;

  INV_1_16 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_357 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_356 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_355 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_354 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_353 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_352 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_351 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_350 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_349 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_348 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_347 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_346 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_345 UND1_4 ( .A(A[4]), .B(SEL), .Y(Y1[4]) );
  NAND_GATE_344 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  NAND_GATE_343 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_342 UND1_5 ( .A(A[5]), .B(SEL), .Y(Y1[5]) );
  NAND_GATE_341 UND2_5 ( .A(B[5]), .B(SB), .Y(Y2[5]) );
  NAND_GATE_340 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_339 UND1_6 ( .A(A[6]), .B(SEL), .Y(Y1[6]) );
  NAND_GATE_338 UND2_6 ( .A(B[6]), .B(SB), .Y(Y2[6]) );
  NAND_GATE_337 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_336 UND1_7 ( .A(A[7]), .B(SEL), .Y(Y1[7]) );
  NAND_GATE_335 UND2_7 ( .A(B[7]), .B(SB), .Y(Y2[7]) );
  NAND_GATE_334 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
endmodule


module MUX21_GEN_N8_3 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;
  wire   SB;
  wire   [7:0] Y1;
  wire   [7:0] Y2;

  INV_1_15 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_333 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_332 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_331 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_330 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_329 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_328 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_327 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_326 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_325 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_324 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_323 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_322 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_321 UND1_4 ( .A(A[4]), .B(SEL), .Y(Y1[4]) );
  NAND_GATE_320 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  NAND_GATE_319 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_318 UND1_5 ( .A(A[5]), .B(SEL), .Y(Y1[5]) );
  NAND_GATE_317 UND2_5 ( .A(B[5]), .B(SB), .Y(Y2[5]) );
  NAND_GATE_316 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_315 UND1_6 ( .A(A[6]), .B(SEL), .Y(Y1[6]) );
  NAND_GATE_314 UND2_6 ( .A(B[6]), .B(SB), .Y(Y2[6]) );
  NAND_GATE_313 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_312 UND1_7 ( .A(A[7]), .B(SEL), .Y(Y1[7]) );
  NAND_GATE_311 UND2_7 ( .A(B[7]), .B(SB), .Y(Y2[7]) );
  NAND_GATE_310 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
endmodule


module MUX21_GEN_N8_2 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;
  wire   SB;
  wire   [7:0] Y1;
  wire   [7:0] Y2;

  INV_1_14 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_309 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_308 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_307 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_306 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_305 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_304 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_303 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_302 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_301 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_300 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_299 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_298 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_297 UND1_4 ( .A(A[4]), .B(SEL), .Y(Y1[4]) );
  NAND_GATE_296 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  NAND_GATE_295 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_294 UND1_5 ( .A(A[5]), .B(SEL), .Y(Y1[5]) );
  NAND_GATE_293 UND2_5 ( .A(B[5]), .B(SB), .Y(Y2[5]) );
  NAND_GATE_292 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_291 UND1_6 ( .A(A[6]), .B(SEL), .Y(Y1[6]) );
  NAND_GATE_290 UND2_6 ( .A(B[6]), .B(SB), .Y(Y2[6]) );
  NAND_GATE_289 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_288 UND1_7 ( .A(A[7]), .B(SEL), .Y(Y1[7]) );
  NAND_GATE_287 UND2_7 ( .A(B[7]), .B(SB), .Y(Y2[7]) );
  NAND_GATE_286 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
endmodule


module MUX21_GEN_N8_1 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;
  wire   SB;
  wire   [7:0] Y1;
  wire   [7:0] Y2;

  INV_1_13 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_285 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_284 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_283 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_282 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_281 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_280 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_279 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_278 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_277 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_276 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_275 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_274 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_273 UND1_4 ( .A(A[4]), .B(SEL), .Y(Y1[4]) );
  NAND_GATE_272 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  NAND_GATE_271 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_270 UND1_5 ( .A(A[5]), .B(SEL), .Y(Y1[5]) );
  NAND_GATE_269 UND2_5 ( .A(B[5]), .B(SB), .Y(Y2[5]) );
  NAND_GATE_268 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_267 UND1_6 ( .A(A[6]), .B(SEL), .Y(Y1[6]) );
  NAND_GATE_266 UND2_6 ( .A(B[6]), .B(SB), .Y(Y2[6]) );
  NAND_GATE_265 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_264 UND1_7 ( .A(A[7]), .B(SEL), .Y(Y1[7]) );
  NAND_GATE_263 UND2_7 ( .A(B[7]), .B(SB), .Y(Y2[7]) );
  NAND_GATE_262 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
endmodule


module N_NAND_N4_31 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_30 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_29 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_28 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_27 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_26 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_25 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_24 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_23 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_22 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_21 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_20 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_19 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_18 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_17 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_16 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_15 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_14 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_13 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_12 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_11 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_10 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_9 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_8 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_7 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_6 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_5 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_4 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_3 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_2 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N4_1 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N3_127 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_126 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_125 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_124 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_123 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_122 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_121 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_120 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_119 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_118 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_117 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_116 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_115 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_114 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_113 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_112 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_111 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_110 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_109 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_108 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_107 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_106 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_105 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_104 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_103 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_102 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_101 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_100 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_99 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_98 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_97 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_96 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_95 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_94 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_93 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_92 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_91 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_90 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_89 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_88 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_87 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_86 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_85 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_84 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_83 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_82 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_81 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_80 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_79 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_78 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_77 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_76 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_75 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_74 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_73 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_72 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_71 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_70 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_69 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_68 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_67 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_66 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_65 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_64 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_63 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_62 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_61 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_60 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_59 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_58 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_57 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_56 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_55 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_54 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_53 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_52 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_51 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_50 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_49 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_48 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_47 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_46 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_45 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_44 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_43 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_42 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_41 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_40 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_39 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_38 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_37 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_36 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_35 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_34 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_33 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_32 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_31 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_30 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_29 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_28 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_27 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_26 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_25 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_24 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_23 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_22 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_21 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_20 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_19 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_18 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_17 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_16 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_15 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_14 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_13 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_12 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_11 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_10 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_9 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_8 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_7 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_6 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_5 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_4 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_3 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_2 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module N_NAND_N3_1 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module NOR_GATE_337 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_336 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_335 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_334 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_333 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_332 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_331 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_330 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_329 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_328 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_327 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_326 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_325 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_324 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_323 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_322 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_321 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_320 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_319 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_318 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_317 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_316 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_315 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_314 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_313 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_312 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_311 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_310 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_309 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_308 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_307 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_306 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_305 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_304 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_303 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_302 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_301 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_300 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_299 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_298 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_297 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_296 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_295 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_294 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_293 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_292 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_291 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_290 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_289 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_288 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_287 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_286 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_285 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_284 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_283 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_282 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_281 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_280 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_279 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_278 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_277 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_276 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_275 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_274 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_273 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_272 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_271 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_270 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_269 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_268 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_267 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_266 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_265 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_264 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_263 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_262 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_261 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_260 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_259 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_258 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_257 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_256 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_255 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_254 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_253 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_252 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_251 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_250 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_249 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_248 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_247 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_246 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_245 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_244 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_243 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_242 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_241 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_240 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_239 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_238 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_237 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_236 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_235 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_234 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_233 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_232 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_231 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_230 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_229 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_228 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_227 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_226 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_225 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_224 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_223 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_222 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_221 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_220 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_219 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_218 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_217 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_216 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_215 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_214 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_213 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_212 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_211 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_210 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_209 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_208 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_207 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_206 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_205 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_204 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_203 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_202 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_201 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_200 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_199 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_198 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_197 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_196 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_195 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_194 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_193 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_192 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_191 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_190 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_189 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_188 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_187 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_186 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_185 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_184 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_183 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_182 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_181 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_180 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_179 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_178 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_177 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_176 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_175 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_174 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_173 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_172 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_171 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_170 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_169 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_168 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_167 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_166 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_165 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_164 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_163 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_162 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_161 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_160 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_159 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_158 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_157 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_156 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_155 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_154 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_153 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_152 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_151 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_150 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_149 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_148 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_147 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_146 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_145 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_144 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_143 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_142 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_141 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_140 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_139 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_138 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_137 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_136 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_135 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_134 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_133 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_132 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_131 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_130 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_129 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_128 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_127 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_126 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_125 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_124 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_123 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_122 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_121 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_120 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_119 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_118 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_117 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_116 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_115 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_114 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_113 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_112 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_111 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_110 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_109 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_108 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_107 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_106 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_105 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_104 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_103 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_102 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_101 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_100 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_99 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_98 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_97 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_96 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_95 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_94 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_93 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_92 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_91 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_90 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_89 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_88 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_87 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_86 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_85 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_84 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_83 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_82 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_81 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_80 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_79 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_78 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_77 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_76 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_75 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_74 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_73 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_72 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_71 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_70 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_69 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_68 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_67 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_66 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_65 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_64 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_63 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_62 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_61 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_60 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_59 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_58 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_57 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_56 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_55 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_54 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_53 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_52 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_51 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_50 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_49 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_48 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_47 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_46 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_45 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_44 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_43 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_42 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_41 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_40 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_39 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_38 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_37 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_36 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_35 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_34 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_33 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_32 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_31 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_30 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_29 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_28 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_27 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_26 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_25 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_24 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_23 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_22 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_21 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_20 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_19 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_18 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_17 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_16 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_15 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_14 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_13 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_12 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_11 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_10 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_9 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_8 ( A, B, Y );
  input A, B;
  output Y;
  wire   n2;

  BUF_X1 U1 ( .A(n2), .Z(Y) );
  NOR2_X1 U2 ( .A1(B), .A2(A), .ZN(n2) );
endmodule


module NOR_GATE_7 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_6 ( A, B, Y );
  input A, B;
  output Y;
  wire   n2;

  BUF_X1 U1 ( .A(n2), .Z(Y) );
  NOR2_X1 U2 ( .A1(B), .A2(A), .ZN(n2) );
endmodule


module NOR_GATE_5 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_4 ( A, B, Y );
  input A, B;
  output Y;
  wire   n2;

  BUF_X1 U1 ( .A(n2), .Z(Y) );
  NOR2_X1 U2 ( .A1(B), .A2(A), .ZN(n2) );
endmodule


module NOR_GATE_3 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NOR_GATE_2 ( A, B, Y );
  input A, B;
  output Y;
  wire   n2;

  BUF_X1 U1 ( .A(n2), .Z(Y) );
  NOR2_X1 U2 ( .A1(B), .A2(A), .ZN(n2) );
endmodule


module NOR_GATE_1 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module N_AND_N32_4 ( A, Y );
  input [31:0] A;
  output Y;
  wire   n11, n12, n13, n14, n15, n16, n17, n18, n19, n20;

  NAND4_X1 U1 ( .A1(A[23]), .A2(A[22]), .A3(A[21]), .A4(A[20]), .ZN(n15) );
  NAND4_X1 U2 ( .A1(A[9]), .A2(A[8]), .A3(A[7]), .A4(A[6]), .ZN(n11) );
  NAND4_X1 U3 ( .A1(A[1]), .A2(A[19]), .A3(A[18]), .A4(A[17]), .ZN(n16) );
  NAND4_X1 U4 ( .A1(A[5]), .A2(A[4]), .A3(A[3]), .A4(A[31]), .ZN(n12) );
  NAND4_X1 U5 ( .A1(A[16]), .A2(A[15]), .A3(A[14]), .A4(A[13]), .ZN(n17) );
  NAND4_X1 U6 ( .A1(A[30]), .A2(A[2]), .A3(A[29]), .A4(A[28]), .ZN(n13) );
  NAND4_X1 U7 ( .A1(A[12]), .A2(A[11]), .A3(A[10]), .A4(A[0]), .ZN(n18) );
  NAND4_X1 U8 ( .A1(A[27]), .A2(A[26]), .A3(A[25]), .A4(A[24]), .ZN(n14) );
  AND2_X1 U9 ( .A1(n20), .A2(n19), .ZN(Y) );
  NOR4_X1 U10 ( .A1(n14), .A2(n13), .A3(n12), .A4(n11), .ZN(n20) );
  NOR4_X1 U11 ( .A1(n18), .A2(n17), .A3(n16), .A4(n15), .ZN(n19) );
endmodule


module N_AND_N32_3 ( A, Y );
  input [31:0] A;
  output Y;
  wire   n11, n12, n13, n14, n15, n16, n17, n18, n19, n20;

  NAND4_X1 U1 ( .A1(A[23]), .A2(A[22]), .A3(A[21]), .A4(A[20]), .ZN(n15) );
  NAND4_X1 U2 ( .A1(A[9]), .A2(A[8]), .A3(A[7]), .A4(A[6]), .ZN(n11) );
  NAND4_X1 U3 ( .A1(A[1]), .A2(A[19]), .A3(A[18]), .A4(A[17]), .ZN(n16) );
  NAND4_X1 U4 ( .A1(A[5]), .A2(A[4]), .A3(A[3]), .A4(A[31]), .ZN(n12) );
  NAND4_X1 U5 ( .A1(A[16]), .A2(A[15]), .A3(A[14]), .A4(A[13]), .ZN(n17) );
  NAND4_X1 U6 ( .A1(A[30]), .A2(A[2]), .A3(A[29]), .A4(A[28]), .ZN(n13) );
  NAND4_X1 U7 ( .A1(A[12]), .A2(A[11]), .A3(A[10]), .A4(A[0]), .ZN(n18) );
  NAND4_X1 U8 ( .A1(A[27]), .A2(A[26]), .A3(A[25]), .A4(A[24]), .ZN(n14) );
  AND2_X1 U9 ( .A1(n20), .A2(n19), .ZN(Y) );
  NOR4_X1 U10 ( .A1(n14), .A2(n13), .A3(n12), .A4(n11), .ZN(n20) );
  NOR4_X1 U11 ( .A1(n18), .A2(n17), .A3(n16), .A4(n15), .ZN(n19) );
endmodule


module N_AND_N32_2 ( A, Y );
  input [31:0] A;
  output Y;
  wire   n11, n12, n13, n14, n15, n16, n17, n18, n19, n20;

  NAND4_X1 U1 ( .A1(A[23]), .A2(A[22]), .A3(A[21]), .A4(A[20]), .ZN(n15) );
  NAND4_X1 U2 ( .A1(A[9]), .A2(A[8]), .A3(A[7]), .A4(A[6]), .ZN(n11) );
  NAND4_X1 U3 ( .A1(A[1]), .A2(A[19]), .A3(A[18]), .A4(A[17]), .ZN(n16) );
  NAND4_X1 U4 ( .A1(A[5]), .A2(A[4]), .A3(A[3]), .A4(A[31]), .ZN(n12) );
  NAND4_X1 U5 ( .A1(A[16]), .A2(A[15]), .A3(A[14]), .A4(A[13]), .ZN(n17) );
  NAND4_X1 U6 ( .A1(A[30]), .A2(A[2]), .A3(A[29]), .A4(A[28]), .ZN(n13) );
  NAND4_X1 U7 ( .A1(A[12]), .A2(A[11]), .A3(A[10]), .A4(A[0]), .ZN(n18) );
  NAND4_X1 U8 ( .A1(A[27]), .A2(A[26]), .A3(A[25]), .A4(A[24]), .ZN(n14) );
  AND2_X1 U9 ( .A1(n20), .A2(n19), .ZN(Y) );
  NOR4_X1 U10 ( .A1(n14), .A2(n13), .A3(n12), .A4(n11), .ZN(n20) );
  NOR4_X1 U11 ( .A1(n18), .A2(n17), .A3(n16), .A4(n15), .ZN(n19) );
endmodule


module N_AND_N32_1 ( A, Y );
  input [31:0] A;
  output Y;
  wire   n11, n12, n13, n14, n15, n16, n17, n18, n19, n20;

  AND2_X1 U1 ( .A1(n20), .A2(n19), .ZN(Y) );
  NOR4_X1 U2 ( .A1(n18), .A2(n17), .A3(n16), .A4(n15), .ZN(n19) );
  NOR4_X1 U3 ( .A1(n14), .A2(n13), .A3(n12), .A4(n11), .ZN(n20) );
  NAND4_X1 U4 ( .A1(A[12]), .A2(A[11]), .A3(A[10]), .A4(A[0]), .ZN(n18) );
  NAND4_X1 U5 ( .A1(A[9]), .A2(A[8]), .A3(A[7]), .A4(A[6]), .ZN(n11) );
  NAND4_X1 U6 ( .A1(A[23]), .A2(A[22]), .A3(A[21]), .A4(A[20]), .ZN(n15) );
  NAND4_X1 U7 ( .A1(A[5]), .A2(A[4]), .A3(A[3]), .A4(A[31]), .ZN(n12) );
  NAND4_X1 U8 ( .A1(A[1]), .A2(A[19]), .A3(A[18]), .A4(A[17]), .ZN(n16) );
  NAND4_X1 U9 ( .A1(A[30]), .A2(A[2]), .A3(A[29]), .A4(A[28]), .ZN(n13) );
  NAND4_X1 U10 ( .A1(A[16]), .A2(A[15]), .A3(A[14]), .A4(A[13]), .ZN(n17) );
  NAND4_X1 U11 ( .A1(A[27]), .A2(A[26]), .A3(A[25]), .A4(A[24]), .ZN(n14) );
endmodule


module FFT_6 ( T, CLK, EN, RST, Q );
  input T, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 TMP_reg ( .D(n1), .CK(CLK), .Q(Q) );
  XOR2_X1 U4 ( .A(n4), .B(Q), .Z(n5) );
  NAND2_X1 U5 ( .A1(T), .A2(EN), .ZN(n4) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
endmodule


module FFT_5 ( T, CLK, EN, RST, Q );
  input T, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 TMP_reg ( .D(n1), .CK(CLK), .Q(Q) );
  XOR2_X1 U4 ( .A(n4), .B(Q), .Z(n5) );
  NAND2_X1 U5 ( .A1(T), .A2(EN), .ZN(n4) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
endmodule


module FFT_4 ( T, CLK, EN, RST, Q );
  input T, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 TMP_reg ( .D(n1), .CK(CLK), .Q(Q) );
  XOR2_X1 U4 ( .A(n4), .B(Q), .Z(n5) );
  NAND2_X1 U5 ( .A1(T), .A2(EN), .ZN(n4) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
endmodule


module FFT_3 ( T, CLK, EN, RST, Q );
  input T, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 TMP_reg ( .D(n1), .CK(CLK), .Q(Q) );
  XOR2_X1 U4 ( .A(n4), .B(Q), .Z(n5) );
  NAND2_X1 U5 ( .A1(T), .A2(EN), .ZN(n4) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
endmodule


module FFT_2 ( T, CLK, EN, RST, Q );
  input T, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 TMP_reg ( .D(n1), .CK(CLK), .Q(Q) );
  XOR2_X1 U4 ( .A(n4), .B(Q), .Z(n5) );
  NAND2_X1 U5 ( .A1(T), .A2(EN), .ZN(n4) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
endmodule


module FFT_1 ( T, CLK, EN, RST, Q );
  input T, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 TMP_reg ( .D(n1), .CK(CLK), .Q(Q) );
  XOR2_X1 U4 ( .A(n4), .B(Q), .Z(n5) );
  NAND2_X1 U5 ( .A1(T), .A2(EN), .ZN(n4) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
endmodule


module N_AND_N5_6 ( A, Y );
  input [4:0] A;
  output Y;
  wire   n2;

  AND3_X1 U1 ( .A1(A[4]), .A2(A[3]), .A3(n2), .ZN(Y) );
  AND3_X1 U2 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(n2) );
endmodule


module N_AND_N5_5 ( A, Y );
  input [4:0] A;
  output Y;
  wire   n2;

  AND3_X1 U1 ( .A1(A[4]), .A2(A[3]), .A3(n2), .ZN(Y) );
  AND3_X1 U2 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(n2) );
endmodule


module N_AND_N5_4 ( A, Y );
  input [4:0] A;
  output Y;
  wire   n2;

  AND3_X1 U1 ( .A1(A[4]), .A2(A[3]), .A3(n2), .ZN(Y) );
  AND3_X1 U2 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(n2) );
endmodule


module N_AND_N5_3 ( A, Y );
  input [4:0] A;
  output Y;
  wire   n2;

  AND3_X1 U1 ( .A1(A[4]), .A2(A[3]), .A3(n2), .ZN(Y) );
  AND3_X1 U2 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(n2) );
endmodule


module N_AND_N5_2 ( A, Y );
  input [4:0] A;
  output Y;
  wire   n2;

  AND3_X1 U1 ( .A1(A[4]), .A2(A[3]), .A3(n2), .ZN(Y) );
  AND3_X1 U2 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(n2) );
endmodule


module N_AND_N5_1 ( A, Y );
  input [4:0] A;
  output Y;
  wire   n2;

  AND3_X1 U1 ( .A1(A[4]), .A2(A[3]), .A3(n2), .ZN(Y) );
  AND3_X1 U2 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(n2) );
endmodule


module XNOR_GATE_217 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_216 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_215 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_214 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_213 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_212 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_211 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_210 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_209 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_208 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_207 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_206 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_205 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_204 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_203 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_202 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_201 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_200 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_199 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_198 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_197 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_196 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_195 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_194 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_193 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_192 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_191 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_190 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_189 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_188 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_187 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_186 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_185 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_184 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_183 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_182 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_181 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_180 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_179 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_178 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_177 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_176 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_175 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_174 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_173 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_172 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_171 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_170 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_169 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_168 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_167 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_166 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_165 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_164 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_163 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_162 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_161 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_160 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_159 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_158 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_157 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_156 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_155 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_154 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_153 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_152 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_151 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_150 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_149 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_148 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_147 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_146 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_145 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_144 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_143 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_142 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_141 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_140 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_139 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_138 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_137 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_136 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_135 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_134 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_133 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_132 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_131 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_130 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_129 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_128 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_127 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_126 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_125 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_124 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_123 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_122 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_121 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_120 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_119 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_118 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_117 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_116 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_115 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_114 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_113 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_112 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_111 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_110 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_109 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_108 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_107 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_106 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_105 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_104 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_103 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_102 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_101 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_100 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_99 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_98 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_97 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_96 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_95 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_94 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_93 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_92 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_91 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_90 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_89 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_88 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_87 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_86 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_85 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_84 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_83 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_82 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_81 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_80 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_79 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_78 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_77 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_76 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_75 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_74 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_73 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_72 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_71 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_70 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_69 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_68 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_67 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_66 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_65 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_64 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_63 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_62 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_61 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_60 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_59 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_58 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_57 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_56 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_55 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_54 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_53 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_52 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_51 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_50 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_49 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_48 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_47 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_46 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_45 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_44 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_43 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_42 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_41 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_40 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_39 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_38 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_37 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_36 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_35 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_34 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_33 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_32 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_31 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_30 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_29 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_28 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_27 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_26 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_25 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_24 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_23 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_22 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_21 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_20 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_19 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_18 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_17 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_16 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_15 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_14 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_13 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_12 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_11 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_10 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_9 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_8 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_7 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_6 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_5 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_4 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_3 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_2 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XNOR_GATE_1 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module XOR_GATE_1_669 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_668 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_667 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_666 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_665 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_664 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_663 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_662 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_661 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_660 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_659 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_658 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_657 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_656 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_655 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_654 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_653 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_652 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_651 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_650 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_649 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_648 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_647 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_646 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_645 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_644 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_643 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_642 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_641 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_640 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_639 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_638 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_637 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1;

  XNOR2_X2 U1 ( .A(A), .B(n1), .ZN(Y) );
  INV_X1 U2 ( .A(B), .ZN(n1) );
endmodule


module XOR_GATE_1_636 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_635 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_634 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_633 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_632 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_631 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_630 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_629 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_628 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_627 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_626 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_625 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_624 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_623 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_622 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_621 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_620 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_619 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_618 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_617 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_616 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_615 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_614 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_613 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_612 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_611 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_610 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_609 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_608 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_607 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_606 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_605 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_604 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_603 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_602 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_601 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_600 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_599 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_598 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_597 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_596 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_595 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_594 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_593 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_592 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_591 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_590 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_589 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_588 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_587 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_586 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_585 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_584 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_583 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_582 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2, n3, n4;

  NAND2_X1 U1 ( .A1(B), .A2(n2), .ZN(n3) );
  NAND2_X1 U2 ( .A1(n1), .A2(A), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n3), .A2(n4), .ZN(Y) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  INV_X1 U5 ( .A(A), .ZN(n2) );
endmodule


module XOR_GATE_1_581 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_580 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2, n3, n4;

  INV_X1 U1 ( .A(B), .ZN(n1) );
  NAND2_X1 U2 ( .A1(n3), .A2(n4), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n2), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n1), .A2(A), .ZN(n4) );
  INV_X1 U5 ( .A(A), .ZN(n2) );
endmodule


module XOR_GATE_1_579 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_578 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_577 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_576 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_575 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_574 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_573 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_572 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_571 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_570 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_569 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_568 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_567 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_566 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_565 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_564 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_563 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_562 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_561 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_560 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_559 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_558 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_557 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_556 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_555 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_554 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_553 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_552 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_551 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_550 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_549 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_548 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_547 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_546 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_545 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_544 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_543 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_542 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_541 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_540 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_539 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_538 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_537 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_536 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_535 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_534 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_533 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_532 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_531 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_530 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_529 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_528 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_527 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_526 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_525 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_524 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_523 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_522 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_521 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_520 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_519 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_518 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_517 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_516 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_515 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_514 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_513 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_512 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_511 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_510 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_509 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_508 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_507 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_506 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_505 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_504 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_503 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_502 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_501 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_500 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_499 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_498 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_497 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_496 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_495 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_494 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_493 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_492 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_491 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_490 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_489 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_488 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_487 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_486 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_485 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_484 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_483 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_482 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_481 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_480 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_479 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_478 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_477 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_476 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_475 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_474 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_473 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_472 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_471 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_470 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_469 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_468 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_467 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_466 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_465 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_464 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_463 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_462 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_461 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_460 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_459 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_458 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_457 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_456 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_455 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_454 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_453 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_452 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_451 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_450 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_449 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_448 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_447 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_446 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_445 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_444 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_443 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_442 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_441 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_440 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_439 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_438 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_437 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_436 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_435 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_434 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_433 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_432 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_431 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_430 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_429 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_428 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_427 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_426 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_425 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_424 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_423 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_422 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_421 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_420 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_419 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_418 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_417 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1;

  XNOR2_X2 U1 ( .A(A), .B(n1), .ZN(Y) );
  INV_X32 U2 ( .A(B), .ZN(n1) );
endmodule


module XOR_GATE_1_416 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_415 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_414 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_413 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_412 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2, n3, n4;

  NAND2_X1 U1 ( .A1(n3), .A2(n4), .ZN(Y) );
  NAND2_X1 U2 ( .A1(B), .A2(n2), .ZN(n3) );
  NAND2_X1 U3 ( .A1(n1), .A2(A), .ZN(n4) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  INV_X1 U5 ( .A(A), .ZN(n2) );
endmodule


module XOR_GATE_1_411 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_410 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_409 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_408 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_407 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_406 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_405 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_404 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_403 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_402 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_401 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_400 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_399 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_398 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_397 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_396 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_395 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_394 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_393 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_392 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X2 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_391 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_390 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_389 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_388 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2, n3, n4;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  NAND2_X4 U2 ( .A1(B), .A2(n2), .ZN(n3) );
  NAND2_X2 U3 ( .A1(n1), .A2(A), .ZN(n4) );
  NAND2_X4 U4 ( .A1(n3), .A2(n4), .ZN(Y) );
  INV_X1 U5 ( .A(B), .ZN(n1) );
endmodule


module XOR_GATE_1_387 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_386 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_385 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_384 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_383 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_382 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2, n3, n4;

  NAND2_X1 U1 ( .A1(A), .A2(n2), .ZN(n3) );
  NAND2_X1 U2 ( .A1(n1), .A2(B), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n3), .A2(n4), .ZN(Y) );
  INV_X1 U4 ( .A(A), .ZN(n1) );
  INV_X1 U5 ( .A(B), .ZN(n2) );
endmodule


module XOR_GATE_1_381 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_380 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_379 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_378 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_377 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2, n3, n4;

  NAND2_X1 U1 ( .A1(n3), .A2(n4), .ZN(Y) );
  NAND2_X1 U2 ( .A1(B), .A2(n2), .ZN(n3) );
  NAND2_X1 U3 ( .A1(n1), .A2(A), .ZN(n4) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  INV_X1 U5 ( .A(A), .ZN(n2) );
endmodule


module XOR_GATE_1_376 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_375 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2, n3, n4;

  NAND2_X1 U1 ( .A1(n3), .A2(n4), .ZN(Y) );
  NAND2_X1 U2 ( .A1(B), .A2(n2), .ZN(n3) );
  NAND2_X1 U3 ( .A1(n1), .A2(A), .ZN(n4) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  INV_X1 U5 ( .A(A), .ZN(n2) );
endmodule


module XOR_GATE_1_374 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_373 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_372 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_371 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2, n3, n4;

  NAND2_X1 U1 ( .A1(n3), .A2(n4), .ZN(Y) );
  NAND2_X1 U2 ( .A1(B), .A2(n2), .ZN(n3) );
  NAND2_X1 U3 ( .A1(n1), .A2(A), .ZN(n4) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  INV_X1 U5 ( .A(A), .ZN(n2) );
endmodule


module XOR_GATE_1_370 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_369 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_368 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2, n3, n4;

  NAND2_X1 U1 ( .A1(n3), .A2(n4), .ZN(Y) );
  NAND2_X1 U2 ( .A1(A), .A2(n2), .ZN(n3) );
  NAND2_X1 U3 ( .A1(n1), .A2(B), .ZN(n4) );
  INV_X1 U4 ( .A(A), .ZN(n1) );
  INV_X1 U5 ( .A(B), .ZN(n2) );
endmodule


module XOR_GATE_1_367 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_366 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_365 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_364 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_363 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X2 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_362 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_361 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_360 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_359 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2, n3, n4;

  NAND2_X1 U1 ( .A1(n3), .A2(n4), .ZN(Y) );
  NAND2_X1 U2 ( .A1(B), .A2(n2), .ZN(n3) );
  NAND2_X1 U3 ( .A1(n1), .A2(A), .ZN(n4) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  INV_X1 U5 ( .A(A), .ZN(n2) );
endmodule


module XOR_GATE_1_358 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_357 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X2 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_356 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_355 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2, n3, n4;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  NAND2_X2 U2 ( .A1(B), .A2(n2), .ZN(n3) );
  NAND2_X2 U3 ( .A1(n1), .A2(A), .ZN(n4) );
  NAND2_X2 U4 ( .A1(n3), .A2(n4), .ZN(Y) );
  INV_X1 U5 ( .A(B), .ZN(n1) );
endmodule


module XOR_GATE_1_354 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_353 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X2 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_352 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_351 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2, n3, n4;

  NAND2_X2 U1 ( .A1(n3), .A2(n4), .ZN(Y) );
  NAND2_X1 U2 ( .A1(B), .A2(n2), .ZN(n3) );
  NAND2_X1 U3 ( .A1(n1), .A2(A), .ZN(n4) );
  INV_X1 U4 ( .A(A), .ZN(n2) );
  INV_X1 U5 ( .A(B), .ZN(n1) );
endmodule


module XOR_GATE_1_350 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_349 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_348 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_347 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_346 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_345 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(n1), .ZN(Y) );
  INV_X1 U2 ( .A(B), .ZN(n1) );
endmodule


module XOR_GATE_1_344 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_343 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2, n3, n4;

  NAND2_X1 U1 ( .A1(n3), .A2(n4), .ZN(Y) );
  NAND2_X1 U2 ( .A1(n1), .A2(B), .ZN(n4) );
  NAND2_X1 U3 ( .A1(A), .A2(n2), .ZN(n3) );
  INV_X1 U4 ( .A(A), .ZN(n1) );
  INV_X1 U5 ( .A(B), .ZN(n2) );
endmodule


module XOR_GATE_1_342 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_341 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_340 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_339 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2, n3, n4;

  NAND2_X1 U1 ( .A1(n3), .A2(n4), .ZN(Y) );
  NAND2_X1 U2 ( .A1(n1), .A2(B), .ZN(n4) );
  NAND2_X1 U3 ( .A1(A), .A2(n2), .ZN(n3) );
  INV_X1 U4 ( .A(A), .ZN(n1) );
  INV_X1 U5 ( .A(B), .ZN(n2) );
endmodule


module XOR_GATE_1_338 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_337 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_336 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_335 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_334 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_333 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_332 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_331 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1;

  INV_X1 U1 ( .A(B), .ZN(n1) );
  XNOR2_X2 U2 ( .A(A), .B(n1), .ZN(Y) );
endmodule


module XOR_GATE_1_330 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_329 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_328 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_327 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_326 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_325 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X2 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_324 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_323 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1;

  INV_X1 U1 ( .A(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(A), .B(n1), .ZN(Y) );
endmodule


module XOR_GATE_1_322 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_321 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1;

  XNOR2_X2 U1 ( .A(A), .B(n1), .ZN(Y) );
  INV_X1 U2 ( .A(B), .ZN(n1) );
endmodule


module XOR_GATE_1_320 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_319 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1;

  XNOR2_X2 U1 ( .A(A), .B(n1), .ZN(Y) );
  INV_X1 U2 ( .A(B), .ZN(n1) );
endmodule


module XOR_GATE_1_318 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_317 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_316 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_315 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_314 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2, n3, n4;

  INV_X1 U1 ( .A(B), .ZN(n1) );
  NAND2_X1 U2 ( .A1(B), .A2(n2), .ZN(n3) );
  NAND2_X1 U3 ( .A1(n1), .A2(A), .ZN(n4) );
  NAND2_X1 U4 ( .A1(n4), .A2(n3), .ZN(Y) );
  INV_X1 U5 ( .A(A), .ZN(n2) );
endmodule


module XOR_GATE_1_313 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_312 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1;

  XNOR2_X2 U1 ( .A(B), .B(n1), .ZN(Y) );
  INV_X1 U2 ( .A(A), .ZN(n1) );
endmodule


module XOR_GATE_1_311 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_310 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_309 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_308 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_307 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2, n3, n4;

  NAND2_X1 U1 ( .A1(n3), .A2(n4), .ZN(Y) );
  NAND2_X1 U2 ( .A1(B), .A2(n2), .ZN(n3) );
  NAND2_X1 U3 ( .A1(n1), .A2(A), .ZN(n4) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  INV_X1 U5 ( .A(A), .ZN(n2) );
endmodule


module XOR_GATE_1_306 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_305 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_304 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_303 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_302 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_301 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_300 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_299 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_298 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_297 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_296 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_295 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_294 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_293 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_292 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_291 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_290 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_289 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_288 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_287 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_286 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_285 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_284 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_283 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_282 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_281 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_280 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_279 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X2 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_278 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_277 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2, n3, n4;

  NAND2_X2 U1 ( .A1(n3), .A2(n4), .ZN(Y) );
  NAND2_X1 U2 ( .A1(B), .A2(n2), .ZN(n3) );
  NAND2_X1 U3 ( .A1(n1), .A2(A), .ZN(n4) );
  INV_X1 U4 ( .A(A), .ZN(n2) );
  INV_X1 U5 ( .A(B), .ZN(n1) );
endmodule


module XOR_GATE_1_276 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_275 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2, n3, n4;

  INV_X1 U1 ( .A(B), .ZN(n2) );
  NAND2_X1 U2 ( .A1(A), .A2(n2), .ZN(n3) );
  NAND2_X1 U3 ( .A1(n1), .A2(B), .ZN(n4) );
  NAND2_X1 U4 ( .A1(n3), .A2(n4), .ZN(Y) );
  INV_X1 U5 ( .A(A), .ZN(n1) );
endmodule


module XOR_GATE_1_274 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_273 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2, n3, n4;

  NAND2_X1 U1 ( .A1(A), .A2(n2), .ZN(n3) );
  NAND2_X1 U2 ( .A1(n1), .A2(B), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n3), .A2(n4), .ZN(Y) );
  INV_X1 U4 ( .A(A), .ZN(n1) );
  INV_X1 U5 ( .A(B), .ZN(n2) );
endmodule


module XOR_GATE_1_272 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_271 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_270 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_269 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_268 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_267 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_266 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_265 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2, n3, n4;

  NAND2_X1 U1 ( .A1(A), .A2(n2), .ZN(n3) );
  NAND2_X2 U2 ( .A1(n1), .A2(B), .ZN(n4) );
  NAND2_X2 U3 ( .A1(n3), .A2(n4), .ZN(Y) );
  INV_X1 U4 ( .A(A), .ZN(n1) );
  INV_X1 U5 ( .A(B), .ZN(n2) );
endmodule


module XOR_GATE_1_264 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_263 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1;

  XNOR2_X2 U1 ( .A(A), .B(n1), .ZN(Y) );
  INV_X32 U2 ( .A(B), .ZN(n1) );
endmodule


module XOR_GATE_1_262 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_261 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_260 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_259 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(n1), .ZN(Y) );
  INV_X32 U2 ( .A(B), .ZN(n1) );
endmodule


module XOR_GATE_1_258 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_257 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_256 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_255 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_254 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_253 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_252 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_251 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_250 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_249 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1;

  INV_X1 U1 ( .A(B), .ZN(n1) );
  XNOR2_X2 U2 ( .A(A), .B(n1), .ZN(Y) );
endmodule


module XOR_GATE_1_248 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_247 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1;

  XNOR2_X2 U1 ( .A(A), .B(n1), .ZN(Y) );
  INV_X32 U2 ( .A(B), .ZN(n1) );
endmodule


module XOR_GATE_1_246 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_245 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(n1), .ZN(Y) );
  INV_X32 U2 ( .A(B), .ZN(n1) );
endmodule


module XOR_GATE_1_244 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_243 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_242 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X2 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_241 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_240 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X2 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_239 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_238 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_237 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_236 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_235 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_234 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_233 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_232 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2, n3, n4;

  NAND2_X1 U1 ( .A1(A), .A2(n2), .ZN(n3) );
  NAND2_X1 U2 ( .A1(n1), .A2(B), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n3), .A2(n4), .ZN(Y) );
  INV_X1 U4 ( .A(A), .ZN(n1) );
  INV_X1 U5 ( .A(B), .ZN(n2) );
endmodule


module XOR_GATE_1_231 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_230 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1;

  INV_X1 U1 ( .A(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(A), .B(n1), .ZN(Y) );
endmodule


module XOR_GATE_1_229 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_228 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1;

  INV_X1 U1 ( .A(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(A), .B(n1), .ZN(Y) );
endmodule


module XOR_GATE_1_227 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_226 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_225 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_224 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_223 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_222 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_221 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_220 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_219 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_218 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1;

  XNOR2_X2 U1 ( .A(A), .B(n1), .ZN(Y) );
  INV_X32 U2 ( .A(B), .ZN(n1) );
endmodule


module XOR_GATE_1_217 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_216 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_215 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_214 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_213 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_212 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1;

  XNOR2_X2 U1 ( .A(A), .B(n1), .ZN(Y) );
  INV_X1 U2 ( .A(B), .ZN(n1) );
endmodule


module XOR_GATE_1_211 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_210 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1;

  XNOR2_X2 U1 ( .A(A), .B(n1), .ZN(Y) );
  INV_X1 U2 ( .A(B), .ZN(n1) );
endmodule


module XOR_GATE_1_209 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_208 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1;

  INV_X1 U1 ( .A(B), .ZN(n1) );
  XNOR2_X2 U2 ( .A(A), .B(n1), .ZN(Y) );
endmodule


module XOR_GATE_1_207 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_206 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_205 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_204 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_203 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_202 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_201 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_200 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_199 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_198 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_197 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_196 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_195 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_194 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_193 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_192 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_191 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_190 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_189 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_188 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_187 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_186 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_185 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_184 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_183 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_182 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_181 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_180 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_179 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_178 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_177 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_176 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_175 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_174 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_173 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_172 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_171 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_170 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_169 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_168 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_167 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_166 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2, n3, n4;

  NAND2_X2 U1 ( .A1(n3), .A2(n4), .ZN(Y) );
  INV_X1 U2 ( .A(A), .ZN(n2) );
  NAND2_X1 U3 ( .A1(n1), .A2(A), .ZN(n4) );
  NAND2_X1 U4 ( .A1(B), .A2(n2), .ZN(n3) );
  INV_X1 U5 ( .A(B), .ZN(n1) );
endmodule


module XOR_GATE_1_165 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_164 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_163 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_162 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_161 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_160 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(A), .B(B), .Z(Y) );
endmodule


module XOR_GATE_1_159 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_158 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2, n3, n4;

  NAND2_X1 U1 ( .A1(B), .A2(n2), .ZN(n3) );
  NAND2_X1 U2 ( .A1(n1), .A2(A), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n3), .A2(n4), .ZN(Y) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  INV_X1 U5 ( .A(A), .ZN(n2) );
endmodule


module XOR_GATE_1_157 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_156 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_155 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_154 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_153 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_152 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_151 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_150 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_149 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_148 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_147 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_146 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_145 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_144 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_143 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_142 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_141 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_140 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_139 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_138 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_137 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_136 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_135 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_134 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1;

  XNOR2_X1 U1 ( .A(n1), .B(A), .ZN(Y) );
  INV_X32 U2 ( .A(B), .ZN(n1) );
endmodule


module XOR_GATE_1_133 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_132 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_131 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_130 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_129 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X2 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_128 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_127 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_126 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_125 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_124 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_123 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_122 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_121 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_120 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_119 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_118 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_117 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_116 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_115 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_114 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_113 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_112 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_111 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_110 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_109 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_108 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_107 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_106 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_105 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_104 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_103 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_102 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_101 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_100 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_99 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_98 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_97 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_96 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_95 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_94 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_93 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_92 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_91 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_90 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_89 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_88 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_87 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_86 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_85 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_84 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_83 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_82 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_81 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_80 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_79 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_78 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_77 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_76 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_75 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_74 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_73 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_72 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_71 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_70 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_69 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_68 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_67 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_66 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_65 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_64 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_63 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_62 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_61 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_60 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_59 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_58 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_57 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_56 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_55 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_54 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_53 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_52 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_51 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_50 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_49 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_48 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_47 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_46 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_45 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_44 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_43 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_42 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_41 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_40 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_39 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_38 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_37 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_36 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_35 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_34 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_33 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_32 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_31 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_30 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_29 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_28 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_27 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_26 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_25 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_24 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_23 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_22 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_21 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_20 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_19 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_18 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_17 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_16 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_15 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_14 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_13 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_12 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_11 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_10 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_9 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_8 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_7 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_6 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_5 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_4 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_3 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_2 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module XOR_GATE_1_1 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module D_LATCH_168 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_168 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_336 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_335 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_336 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_335 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_167 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_167 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_334 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_333 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_334 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_333 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_166 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_166 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_332 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_331 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_332 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_331 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_165 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_165 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_330 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_329 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_330 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_329 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_164 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_164 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_328 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_327 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_328 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_327 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_163 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_163 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_326 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_325 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_326 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_325 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_162 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_162 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_324 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_323 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_324 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_323 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_161 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_161 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_322 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_321 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_322 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_321 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_160 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_160 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_320 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_319 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_320 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_319 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_159 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_159 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_318 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_317 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_318 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_317 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_158 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_158 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_316 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_315 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_316 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_315 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_157 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_157 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_314 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_313 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_314 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_313 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_156 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_156 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_312 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_311 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_312 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_311 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_155 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_155 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_310 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_309 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_310 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_309 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_154 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_154 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_308 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_307 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_308 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_307 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_153 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_153 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_306 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_305 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_306 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_305 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_152 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_152 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_304 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_303 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_304 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_303 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_151 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_151 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_302 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_301 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_302 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_301 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_150 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_150 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_300 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_299 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_300 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_299 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_149 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_149 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_298 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_297 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_298 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_297 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_148 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_148 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_296 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_295 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_296 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_295 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_147 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_147 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_294 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_293 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_294 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_293 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_146 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_146 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_292 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_291 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_292 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_291 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_145 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_145 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_290 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_289 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_290 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_289 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_144 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_144 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_288 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_287 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_288 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_287 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_143 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_143 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_286 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_285 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_286 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_285 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_142 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_142 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_284 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_283 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_284 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_283 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_141 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_141 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_282 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_281 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_282 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_281 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_140 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_140 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_280 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_279 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_280 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_279 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_139 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_139 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_278 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_277 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_278 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_277 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_138 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_138 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_276 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_275 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_276 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_275 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_137 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_137 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_274 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_273 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_274 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_273 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_136 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_136 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_272 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_271 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_272 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_271 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_135 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_135 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_270 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_269 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_270 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_269 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_134 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_134 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_268 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_267 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_268 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_267 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_133 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_133 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_266 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_265 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_266 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_265 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_132 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_132 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_264 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_263 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_264 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_263 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_131 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_131 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_262 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_261 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_262 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_261 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_130 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_130 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_260 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_259 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_260 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_259 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_129 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_129 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_258 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_257 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_258 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_257 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_128 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_128 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_256 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_255 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_256 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_255 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_127 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_127 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_254 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_253 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_254 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_253 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_126 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_126 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_252 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_251 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_252 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_251 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_125 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_125 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_250 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_249 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_250 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_249 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_124 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_124 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_248 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_247 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_248 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_247 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_123 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_123 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_246 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_245 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_246 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_245 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_122 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_122 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_244 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_243 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_244 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_243 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_121 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_121 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_242 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_241 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_242 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_241 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_120 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_120 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_240 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_239 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_240 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_239 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_119 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_119 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_238 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_237 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_238 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_237 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_118 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_118 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_236 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_235 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_236 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_235 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_117 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_117 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_234 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_233 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_234 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_233 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_116 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_116 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_232 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_231 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_232 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_231 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_115 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_115 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_230 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_229 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_230 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_229 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_114 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_114 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_228 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_227 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_228 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_227 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_113 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_113 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_226 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_225 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_226 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_225 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_112 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_112 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_224 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_223 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_224 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_223 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_111 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_111 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_222 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_221 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_222 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_221 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_110 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_110 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_220 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_219 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_220 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_219 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_109 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_109 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_218 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_217 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_218 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_217 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_108 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_108 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_216 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_215 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_216 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_215 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_107 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_107 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_214 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_213 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_214 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_213 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_106 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_106 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_212 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_211 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_212 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_211 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_105 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_105 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_210 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_209 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_210 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_209 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_104 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_104 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_208 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_207 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_208 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_207 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_103 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_103 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_206 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_205 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_206 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_205 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_102 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_102 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_204 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_203 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_204 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_203 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_101 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_101 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_202 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_201 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_202 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_201 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_100 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_100 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_200 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_199 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_200 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_199 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_99 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_99 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_198 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_197 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_198 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_197 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_98 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_98 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_196 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_195 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_196 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_195 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_97 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_97 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_194 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_193 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_194 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_193 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_96 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_96 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_192 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_191 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_192 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_191 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_95 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_95 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_190 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_189 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_190 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_189 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_94 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_94 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_188 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_187 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_188 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_187 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_93 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_93 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_186 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_185 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_186 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_185 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_92 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_92 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_184 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_183 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_184 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_183 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_91 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_91 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_182 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_181 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_182 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_181 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_90 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_90 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_180 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_179 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_180 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_179 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_89 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_89 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_178 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_177 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_178 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_177 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_88 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_88 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_176 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_175 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_176 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_175 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_87 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_87 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_174 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_173 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_174 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_173 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_86 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_86 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_172 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_171 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_172 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_171 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_85 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_85 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_170 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_169 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_170 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_169 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_84 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_84 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_168 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_167 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_168 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_167 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_83 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_83 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_166 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_165 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_166 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_165 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_82 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_82 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_164 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_163 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_164 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_163 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_81 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_81 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_162 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_161 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_162 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_161 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_80 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_80 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_160 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_159 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_160 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_159 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_79 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_79 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_158 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_157 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_158 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_157 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_78 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_78 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_156 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_155 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_156 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_155 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_77 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_77 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_154 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_153 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_154 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_153 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_76 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_76 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_152 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_151 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_152 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_151 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_75 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_75 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_150 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_149 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_150 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_149 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_74 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_74 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_148 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_147 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_148 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_147 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_73 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_73 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_146 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_145 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_146 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_145 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_72 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_72 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_144 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_143 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_144 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_143 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_71 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_71 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_142 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_141 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_142 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_141 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_70 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_70 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_140 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_139 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_140 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_139 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_69 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_69 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_138 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_137 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_138 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_137 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_68 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_68 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_136 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_135 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_136 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_135 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_67 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_67 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_134 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_133 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_134 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_133 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_66 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_66 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_132 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_131 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_132 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_131 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_65 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_65 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_130 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_129 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_130 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_129 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_64 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_64 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_128 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_127 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_128 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_127 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_63 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_63 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_126 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_125 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_126 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_125 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_62 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_62 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_124 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_123 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_124 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_123 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_61 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_61 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_122 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_121 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_122 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_121 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_60 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_60 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_120 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_119 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_120 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_119 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_59 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_59 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_118 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_117 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_118 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_117 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_58 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_58 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_116 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_115 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_116 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_115 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_57 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_57 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_114 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_113 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_114 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_113 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_56 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_56 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_112 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_111 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_112 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_111 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_55 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_55 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_110 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_109 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_110 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_109 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_54 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_54 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_108 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_107 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_108 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_107 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_53 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_53 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_106 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_105 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_106 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_105 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_52 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_52 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_104 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_103 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_104 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_103 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_51 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_51 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_102 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_101 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_102 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_101 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_50 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_50 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_100 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_99 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_100 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_99 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_49 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_49 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_98 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_97 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_98 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_97 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_48 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_48 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_96 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_95 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_96 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_95 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_47 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_47 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_94 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_93 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_94 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_93 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_46 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_46 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_92 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_91 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_92 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_91 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_45 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_45 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_90 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_89 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_90 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_89 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_44 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_44 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_88 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_87 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_88 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_87 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_43 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_43 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_86 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_85 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_86 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_85 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_42 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_42 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_84 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_83 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_84 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_83 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_41 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_41 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_82 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_81 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_82 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_81 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_40 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_40 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_80 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_79 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_80 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_79 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_39 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_39 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_78 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_77 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_78 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_77 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_38 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_38 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_76 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_75 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_76 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_75 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_37 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_37 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_74 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_73 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_74 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_73 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_36 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_36 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_72 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_71 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_72 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_71 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_35 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_35 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_70 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_69 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_70 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_69 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_34 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_34 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_68 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_67 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_68 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_67 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_33 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_33 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_66 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_65 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_66 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_65 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_32 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_32 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_64 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_63 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_64 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_63 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_31 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_31 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_62 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_61 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_62 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_61 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_30 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_30 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_60 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_59 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_60 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_59 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_29 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_29 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_58 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_57 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_58 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_57 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_28 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_28 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_56 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_55 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_56 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_55 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_27 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_27 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_54 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_53 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_54 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_53 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_26 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_26 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_52 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_51 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_52 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_51 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_25 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_25 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_50 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_49 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_50 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_49 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_24 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_24 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_48 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_47 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_48 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_47 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_23 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_23 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_46 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_45 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_46 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_45 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_22 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_22 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_44 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_43 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_44 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_43 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_21 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_21 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_42 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_41 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_42 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_41 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_20 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_20 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_40 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_39 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_40 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_39 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_19 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_19 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_38 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_37 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_38 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_37 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_18 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_18 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_36 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_35 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_36 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_35 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_17 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_17 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_34 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_33 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_34 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_33 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_16 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_16 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_32 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_31 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_32 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_31 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_15 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_15 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_30 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_29 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_30 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_29 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_14 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_14 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_28 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_27 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_28 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_27 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_13 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_13 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_26 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_25 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_26 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_25 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_12 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_12 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_24 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_23 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_24 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_23 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_11 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_11 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_22 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_21 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_22 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_21 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_10 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_10 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_20 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_19 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_20 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_19 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_9 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_9 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_18 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_17 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_18 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_17 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_8 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_8 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_16 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_15 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_16 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_15 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_7 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_7 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_14 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_13 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_14 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_13 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_6 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_6 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_12 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_11 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_12 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_11 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_5 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_5 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_10 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_9 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_10 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_9 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_4 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_4 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_8 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_7 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_8 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_7 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_3 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_3 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_6 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_5 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_6 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_5 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_2 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_2 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_4 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_3 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_4 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_3 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module D_LATCH_1 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_1 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_2 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_1 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_2 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_1 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module OR_GATE_338 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_337 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_336 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_335 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_334 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_333 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_332 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  INV_X4 U2 ( .A(B), .ZN(n1) );
  NAND2_X4 U3 ( .A1(n1), .A2(n2), .ZN(Y) );
endmodule


module OR_GATE_331 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_330 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_329 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  INV_X4 U2 ( .A(B), .ZN(n1) );
  NAND2_X4 U3 ( .A1(n1), .A2(n2), .ZN(Y) );
endmodule


module OR_GATE_328 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  INV_X4 U2 ( .A(B), .ZN(n1) );
  NAND2_X4 U3 ( .A1(n1), .A2(n2), .ZN(Y) );
endmodule


module OR_GATE_327 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  INV_X4 U2 ( .A(B), .ZN(n1) );
  NAND2_X4 U3 ( .A1(n1), .A2(n2), .ZN(Y) );
endmodule


module OR_GATE_326 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_325 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  INV_X4 U1 ( .A(B), .ZN(n1) );
  INV_X1 U2 ( .A(A), .ZN(n2) );
  NAND2_X4 U3 ( .A1(n1), .A2(n2), .ZN(Y) );
endmodule


module OR_GATE_324 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  INV_X4 U1 ( .A(B), .ZN(n1) );
  INV_X1 U2 ( .A(A), .ZN(n2) );
  NAND2_X4 U3 ( .A1(n1), .A2(n2), .ZN(Y) );
endmodule


module OR_GATE_323 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  INV_X1 U2 ( .A(B), .ZN(n1) );
  NAND2_X4 U3 ( .A1(n1), .A2(n2), .ZN(Y) );
endmodule


module OR_GATE_322 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  NAND2_X2 U1 ( .A1(n1), .A2(n2), .ZN(Y) );
  INV_X1 U2 ( .A(A), .ZN(n2) );
  INV_X1 U3 ( .A(B), .ZN(n1) );
endmodule


module OR_GATE_321 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_320 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_319 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  INV_X2 U1 ( .A(B), .ZN(n1) );
  INV_X1 U2 ( .A(A), .ZN(n2) );
  NAND2_X4 U3 ( .A1(n1), .A2(n2), .ZN(Y) );
endmodule


module OR_GATE_318 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  INV_X4 U2 ( .A(B), .ZN(n1) );
  NAND2_X4 U3 ( .A1(n1), .A2(n2), .ZN(Y) );
endmodule


module OR_GATE_317 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  INV_X4 U2 ( .A(B), .ZN(n1) );
  NAND2_X4 U3 ( .A1(n1), .A2(n2), .ZN(Y) );
endmodule


module OR_GATE_316 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_315 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_314 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  INV_X4 U2 ( .A(B), .ZN(n1) );
  NAND2_X4 U3 ( .A1(n1), .A2(n2), .ZN(Y) );
endmodule


module OR_GATE_313 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  INV_X4 U2 ( .A(B), .ZN(n1) );
  NAND2_X4 U3 ( .A1(n1), .A2(n2), .ZN(Y) );
endmodule


module OR_GATE_312 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_311 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  NAND2_X4 U1 ( .A1(n1), .A2(n2), .ZN(Y) );
  INV_X4 U2 ( .A(B), .ZN(n1) );
  INV_X1 U3 ( .A(A), .ZN(n2) );
endmodule


module OR_GATE_310 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_309 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_308 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_307 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_306 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_305 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_304 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_303 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_302 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_301 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_300 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_299 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_298 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_297 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_296 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_295 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_294 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_293 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_292 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_291 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_290 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_289 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_288 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_287 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_286 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_285 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_284 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_283 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_282 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_281 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_280 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_279 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_278 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_277 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_276 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_275 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_274 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_273 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_272 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_271 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_270 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_269 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_268 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_267 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_266 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_265 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_264 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_263 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_262 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_261 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_260 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_259 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_258 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_257 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_256 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_255 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_254 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_253 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_252 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_251 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_250 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_249 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_248 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_247 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_246 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_245 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_244 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_243 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_242 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_241 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_240 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_239 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_238 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_237 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_236 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_235 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_234 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_233 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_232 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_231 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_230 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_229 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_228 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_227 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_226 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_225 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_224 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_223 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_222 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_221 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_220 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_219 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_218 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_217 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_216 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_215 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_214 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_213 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_212 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_211 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_210 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_209 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_208 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_207 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_206 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_205 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_204 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_203 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_202 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_201 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_200 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_199 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_198 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_197 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_196 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_195 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_194 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_193 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_192 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_191 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_190 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_189 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_188 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_187 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_186 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_185 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_184 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_183 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  INV_X4 U2 ( .A(B), .ZN(n1) );
  NAND2_X4 U3 ( .A1(n1), .A2(n2), .ZN(Y) );
endmodule


module OR_GATE_182 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_181 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_180 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_179 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  INV_X4 U1 ( .A(B), .ZN(n1) );
  NAND2_X4 U2 ( .A1(n1), .A2(n2), .ZN(Y) );
  INV_X32 U3 ( .A(A), .ZN(n2) );
endmodule


module OR_GATE_178 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_177 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_176 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_175 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_174 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_173 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_172 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_171 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  INV_X4 U1 ( .A(B), .ZN(n1) );
  INV_X1 U2 ( .A(A), .ZN(n2) );
  NAND2_X4 U3 ( .A1(n1), .A2(n2), .ZN(Y) );
endmodule


module OR_GATE_170 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_169 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_168 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_167 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  NAND2_X2 U1 ( .A1(n1), .A2(n2), .ZN(Y) );
  INV_X1 U2 ( .A(A), .ZN(n2) );
  INV_X2 U3 ( .A(B), .ZN(n1) );
endmodule


module OR_GATE_166 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n1), .A2(n2), .ZN(Y) );
  INV_X1 U2 ( .A(A), .ZN(n2) );
  INV_X1 U3 ( .A(B), .ZN(n1) );
endmodule


module OR_GATE_165 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n1), .A2(n2), .ZN(Y) );
  INV_X1 U2 ( .A(B), .ZN(n1) );
  INV_X1 U3 ( .A(A), .ZN(n2) );
endmodule


module OR_GATE_164 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n1), .A2(n2), .ZN(Y) );
  INV_X1 U2 ( .A(A), .ZN(n2) );
  INV_X1 U3 ( .A(B), .ZN(n1) );
endmodule


module OR_GATE_163 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_162 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_161 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_160 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  NAND2_X4 U1 ( .A1(n1), .A2(n2), .ZN(Y) );
  INV_X4 U2 ( .A(B), .ZN(n1) );
  INV_X1 U3 ( .A(A), .ZN(n2) );
endmodule


module OR_GATE_159 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_158 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_157 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_156 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_155 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_154 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_153 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  INV_X4 U2 ( .A(B), .ZN(n1) );
  NAND2_X4 U3 ( .A1(n1), .A2(n2), .ZN(Y) );
endmodule


module OR_GATE_152 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_151 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n1), .A2(n2), .ZN(Y) );
  INV_X1 U2 ( .A(A), .ZN(n2) );
  INV_X1 U3 ( .A(B), .ZN(n1) );
endmodule


module OR_GATE_150 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_149 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_148 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_147 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_146 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  NAND2_X4 U1 ( .A1(n1), .A2(n2), .ZN(Y) );
  INV_X4 U2 ( .A(B), .ZN(n1) );
  INV_X32 U3 ( .A(A), .ZN(n2) );
endmodule


module OR_GATE_145 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_144 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_143 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_142 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_141 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_140 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_139 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_138 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_137 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_136 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_135 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_134 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_133 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_132 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_131 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_130 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_129 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  INV_X4 U2 ( .A(B), .ZN(n1) );
  NAND2_X4 U3 ( .A1(n1), .A2(n2), .ZN(Y) );
endmodule


module OR_GATE_128 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_127 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_126 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_125 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_124 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(A), .ZN(n2) );
  INV_X4 U2 ( .A(B), .ZN(n1) );
  NAND2_X4 U3 ( .A1(n1), .A2(n2), .ZN(Y) );
endmodule


module OR_GATE_123 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_122 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_121 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_120 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_119 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_118 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_117 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_116 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_115 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_114 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_113 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_112 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_111 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_110 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_109 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_108 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_107 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_106 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  INV_X2 U1 ( .A(B), .ZN(n1) );
  NAND2_X2 U2 ( .A1(n1), .A2(n2), .ZN(Y) );
  INV_X1 U3 ( .A(A), .ZN(n2) );
endmodule


module OR_GATE_105 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_104 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_103 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_102 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_101 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_100 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module OR_GATE_99 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  NAND2_X2 U1 ( .A1(n1), .A2(n2), .ZN(Y) );
  INV_X4 U2 ( .A(B), .ZN(n2) );
  INV_X1 U3 ( .A(A), .ZN(n1) );
endmodule


module OR_GATE_98 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_97 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_96 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_95 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n1), .A2(n2), .ZN(Y) );
  INV_X1 U2 ( .A(A), .ZN(n1) );
  INV_X1 U3 ( .A(B), .ZN(n2) );
endmodule


module OR_GATE_94 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  NAND2_X2 U1 ( .A1(n1), .A2(n2), .ZN(Y) );
  INV_X4 U2 ( .A(B), .ZN(n2) );
  INV_X1 U3 ( .A(A), .ZN(n1) );
endmodule


module OR_GATE_93 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_92 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_91 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_90 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_89 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_88 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_87 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_86 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_85 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_84 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_83 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_82 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_81 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_80 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_79 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_78 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(A), .ZN(n1) );
  NAND2_X1 U2 ( .A1(n1), .A2(n2), .ZN(Y) );
  INV_X1 U3 ( .A(B), .ZN(n2) );
endmodule


module OR_GATE_77 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_76 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_75 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_74 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_73 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_72 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_71 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_70 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_69 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_68 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n1), .A2(n2), .ZN(Y) );
  INV_X1 U2 ( .A(A), .ZN(n1) );
  INV_X1 U3 ( .A(B), .ZN(n2) );
endmodule


module OR_GATE_67 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(A), .ZN(n1) );
  INV_X4 U2 ( .A(B), .ZN(n2) );
  NAND2_X4 U3 ( .A1(n1), .A2(n2), .ZN(Y) );
endmodule


module OR_GATE_66 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_65 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_64 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_63 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_62 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_61 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_60 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_59 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_58 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_57 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_56 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_55 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_54 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_53 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_52 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_51 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_50 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_49 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_48 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_47 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_46 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_45 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_44 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_43 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_42 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_41 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_40 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_39 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_38 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_37 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_36 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_35 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_34 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_33 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_32 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_31 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_30 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_29 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_28 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_27 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_26 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_25 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_24 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_23 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_22 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_21 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_20 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_19 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_18 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_17 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_16 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_15 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_14 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_13 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_12 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_11 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_10 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_9 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_8 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_7 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_6 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_5 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_4 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_3 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_2 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module OR_GATE_1 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module MUX21_6 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  INV_1_37 UIV ( .A(S), .Y(SB) );
  NAND_GATE_726 UND1 ( .A(A), .B(S), .Y(Y1) );
  NAND_GATE_725 UND2 ( .A(B), .B(SB), .Y(Y2) );
  NAND_GATE_724 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_5 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  INV_1_36 UIV ( .A(S), .Y(SB) );
  NAND_GATE_723 UND1 ( .A(A), .B(S), .Y(Y1) );
  NAND_GATE_722 UND2 ( .A(B), .B(SB), .Y(Y2) );
  NAND_GATE_721 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_4 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  INV_1_35 UIV ( .A(S), .Y(SB) );
  NAND_GATE_720 UND1 ( .A(A), .B(S), .Y(Y1) );
  NAND_GATE_719 UND2 ( .A(B), .B(SB), .Y(Y2) );
  NAND_GATE_718 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_3 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  INV_1_34 UIV ( .A(S), .Y(SB) );
  NAND_GATE_717 UND1 ( .A(A), .B(S), .Y(Y1) );
  NAND_GATE_716 UND2 ( .A(B), .B(SB), .Y(Y2) );
  NAND_GATE_715 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_2 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  INV_1_33 UIV ( .A(S), .Y(SB) );
  NAND_GATE_714 UND1 ( .A(A), .B(S), .Y(Y1) );
  NAND_GATE_713 UND2 ( .A(B), .B(SB), .Y(Y2) );
  NAND_GATE_712 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_1 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  INV_1_32 UIV ( .A(S), .Y(SB) );
  NAND_GATE_711 UND1 ( .A(A), .B(S), .Y(Y1) );
  NAND_GATE_710 UND2 ( .A(B), .B(SB), .Y(Y2) );
  NAND_GATE_709 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GEN_N4_15 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  INV_1_118 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_1005 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_1004 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_1003 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_1002 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_1001 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_1000 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_999 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_998 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_997 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_996 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_995 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_994 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
endmodule


module MUX21_GEN_N4_14 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  INV_1_117 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_993 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_992 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_991 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_990 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_989 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_988 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_987 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_986 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_985 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_984 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_983 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_982 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
endmodule


module MUX21_GEN_N4_13 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  INV_1_116 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_981 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_980 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_979 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_978 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_977 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_976 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_975 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_974 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_973 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_972 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_971 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_970 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
endmodule


module MUX21_GEN_N4_12 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  INV_1_115 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_969 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_968 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_967 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_966 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_965 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_964 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_963 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_962 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_961 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_960 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_959 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_958 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
endmodule


module MUX21_GEN_N4_11 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  INV_1_114 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_957 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_956 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_955 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_954 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_953 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_952 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_951 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_950 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_949 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_948 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_947 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_946 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
endmodule


module MUX21_GEN_N4_10 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  INV_1_113 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_945 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_944 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_943 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_942 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_941 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_940 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_939 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_938 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_937 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_936 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_935 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_934 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
endmodule


module MUX21_GEN_N4_9 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  INV_1_112 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_933 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_932 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_931 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_930 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_929 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_928 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_927 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_926 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_925 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_924 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_923 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_922 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
endmodule


module MUX21_GEN_N4_8 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  INV_1_8 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_96 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_95 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_94 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_93 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_92 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_91 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_90 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_89 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_88 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_87 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_86 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_85 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
endmodule


module MUX21_GEN_N4_7 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  INV_1_7 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_84 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_83 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_82 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_81 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_80 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_79 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_78 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_77 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_76 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_75 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_74 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_73 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
endmodule


module MUX21_GEN_N4_6 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  INV_1_6 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_72 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_71 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_70 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_69 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_68 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_67 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_66 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_65 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_64 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_63 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_62 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_61 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
endmodule


module MUX21_GEN_N4_5 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  INV_1_5 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_60 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_59 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_58 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_57 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_56 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_55 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_54 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_53 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_52 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_51 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_50 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_49 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
endmodule


module MUX21_GEN_N4_4 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  INV_1_4 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_48 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_47 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_46 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_45 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_44 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_43 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_42 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_41 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_40 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_39 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_38 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_37 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
endmodule


module MUX21_GEN_N4_3 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  INV_1_3 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_36 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_35 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_34 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_33 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_32 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_31 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_30 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_29 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_28 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_27 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_26 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_25 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
endmodule


module MUX21_GEN_N4_2 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  INV_1_2 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_24 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_23 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_22 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_21 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_20 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_19 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_18 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_17 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_16 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_15 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_14 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_13 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
endmodule


module MUX21_GEN_N4_1 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  INV_1_1 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_12 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_11 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_10 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_9 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_8 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_7 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_6 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_5 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_4 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_3 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_2 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_1 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
endmodule


module RCA_GEN_N4_31 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_265 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_264 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_263 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_262 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_30 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_261 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_260 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_259 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_258 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_29 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_257 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_256 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_255 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_254 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_28 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_253 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_252 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_251 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_250 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_27 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_249 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_248 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_247 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_246 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_26 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_245 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_244 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_243 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_242 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_25 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_241 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_240 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_239 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_238 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_24 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_237 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_236 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_235 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_234 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_23 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_233 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_232 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_231 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_230 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_22 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_229 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_228 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_227 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_226 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_21 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_225 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_224 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_223 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_222 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_20 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_221 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_220 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_219 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_218 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_19 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_217 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_216 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_215 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_214 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_18 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_213 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_212 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_211 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_210 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_17 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_209 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_208 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_207 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_206 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_16 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_64 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_63 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_62 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_61 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_60 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_59 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_58 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_57 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_56 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_55 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_54 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_53 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_52 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_51 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_50 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_49 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_48 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_47 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_46 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_45 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_44 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_43 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_42 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_41 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_40 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_39 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_38 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_37 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_36 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_35 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_34 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_33 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_32 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_31 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_30 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_29 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_28 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_27 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_26 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_25 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_24 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_23 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_22 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_21 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_20 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_19 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_18 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_17 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_16 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_15 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_14 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_13 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_12 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_11 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_10 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_9 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_8 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_7 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_6 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_5 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_N4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_4 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_3 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_2 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX41_1 ( A, B, C, D, SEL, Y );
  input [1:0] SEL;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n3, n4, n8, n9, n10;

  NAND2_X1 U8 ( .A1(A), .A2(n10), .ZN(n8) );
  INV_X1 U1 ( .A(SEL[0]), .ZN(n1) );
  INV_X1 U2 ( .A(SEL[1]), .ZN(n3) );
  OAI21_X1 U3 ( .B1(n10), .B2(n9), .A(n8), .ZN(Y) );
  NOR2_X1 U4 ( .A1(n3), .A2(n1), .ZN(n10) );
  AOI22_X1 U5 ( .A1(n4), .A2(n3), .B1(B), .B2(SEL[1]), .ZN(n9) );
  INV_X1 U6 ( .A(n2), .ZN(n4) );
  AOI22_X1 U7 ( .A1(C), .A2(SEL[0]), .B1(D), .B2(n1), .ZN(n2) );
endmodule


module EQU_COMPARATOR_N32_4 ( A, B, Y );
  input [31:0] A;
  input [31:0] B;
  output Y;

  wire   [31:0] L;

  XNOR_GATE_128 XNORING_0 ( .A(A[0]), .B(B[0]), .Y(L[0]) );
  XNOR_GATE_127 XNORING_1 ( .A(A[1]), .B(B[1]), .Y(L[1]) );
  XNOR_GATE_126 XNORING_2 ( .A(A[2]), .B(B[2]), .Y(L[2]) );
  XNOR_GATE_125 XNORING_3 ( .A(A[3]), .B(B[3]), .Y(L[3]) );
  XNOR_GATE_124 XNORING_4 ( .A(A[4]), .B(B[4]), .Y(L[4]) );
  XNOR_GATE_123 XNORING_5 ( .A(A[5]), .B(B[5]), .Y(L[5]) );
  XNOR_GATE_122 XNORING_6 ( .A(A[6]), .B(B[6]), .Y(L[6]) );
  XNOR_GATE_121 XNORING_7 ( .A(A[7]), .B(B[7]), .Y(L[7]) );
  XNOR_GATE_120 XNORING_8 ( .A(A[8]), .B(B[8]), .Y(L[8]) );
  XNOR_GATE_119 XNORING_9 ( .A(A[9]), .B(B[9]), .Y(L[9]) );
  XNOR_GATE_118 XNORING_10 ( .A(A[10]), .B(B[10]), .Y(L[10]) );
  XNOR_GATE_117 XNORING_11 ( .A(A[11]), .B(B[11]), .Y(L[11]) );
  XNOR_GATE_116 XNORING_12 ( .A(A[12]), .B(B[12]), .Y(L[12]) );
  XNOR_GATE_115 XNORING_13 ( .A(A[13]), .B(B[13]), .Y(L[13]) );
  XNOR_GATE_114 XNORING_14 ( .A(A[14]), .B(B[14]), .Y(L[14]) );
  XNOR_GATE_113 XNORING_15 ( .A(A[15]), .B(B[15]), .Y(L[15]) );
  XNOR_GATE_112 XNORING_16 ( .A(A[16]), .B(B[16]), .Y(L[16]) );
  XNOR_GATE_111 XNORING_17 ( .A(A[17]), .B(B[17]), .Y(L[17]) );
  XNOR_GATE_110 XNORING_18 ( .A(A[18]), .B(B[18]), .Y(L[18]) );
  XNOR_GATE_109 XNORING_19 ( .A(A[19]), .B(B[19]), .Y(L[19]) );
  XNOR_GATE_108 XNORING_20 ( .A(A[20]), .B(B[20]), .Y(L[20]) );
  XNOR_GATE_107 XNORING_21 ( .A(A[21]), .B(B[21]), .Y(L[21]) );
  XNOR_GATE_106 XNORING_22 ( .A(A[22]), .B(B[22]), .Y(L[22]) );
  XNOR_GATE_105 XNORING_23 ( .A(A[23]), .B(B[23]), .Y(L[23]) );
  XNOR_GATE_104 XNORING_24 ( .A(A[24]), .B(B[24]), .Y(L[24]) );
  XNOR_GATE_103 XNORING_25 ( .A(A[25]), .B(B[25]), .Y(L[25]) );
  XNOR_GATE_102 XNORING_26 ( .A(A[26]), .B(B[26]), .Y(L[26]) );
  XNOR_GATE_101 XNORING_27 ( .A(A[27]), .B(B[27]), .Y(L[27]) );
  XNOR_GATE_100 XNORING_28 ( .A(A[28]), .B(B[28]), .Y(L[28]) );
  XNOR_GATE_99 XNORING_29 ( .A(A[29]), .B(B[29]), .Y(L[29]) );
  XNOR_GATE_98 XNORING_30 ( .A(A[30]), .B(B[30]), .Y(L[30]) );
  XNOR_GATE_97 XNORING_31 ( .A(A[31]), .B(B[31]), .Y(L[31]) );
  N_AND_N32_4 ANDING ( .A(L), .Y(Y) );
endmodule


module EQU_COMPARATOR_N32_3 ( A, B, Y );
  input [31:0] A;
  input [31:0] B;
  output Y;

  wire   [31:0] L;

  XNOR_GATE_96 XNORING_0 ( .A(A[0]), .B(B[0]), .Y(L[0]) );
  XNOR_GATE_95 XNORING_1 ( .A(A[1]), .B(B[1]), .Y(L[1]) );
  XNOR_GATE_94 XNORING_2 ( .A(A[2]), .B(B[2]), .Y(L[2]) );
  XNOR_GATE_93 XNORING_3 ( .A(A[3]), .B(B[3]), .Y(L[3]) );
  XNOR_GATE_92 XNORING_4 ( .A(A[4]), .B(B[4]), .Y(L[4]) );
  XNOR_GATE_91 XNORING_5 ( .A(A[5]), .B(B[5]), .Y(L[5]) );
  XNOR_GATE_90 XNORING_6 ( .A(A[6]), .B(B[6]), .Y(L[6]) );
  XNOR_GATE_89 XNORING_7 ( .A(A[7]), .B(B[7]), .Y(L[7]) );
  XNOR_GATE_88 XNORING_8 ( .A(A[8]), .B(B[8]), .Y(L[8]) );
  XNOR_GATE_87 XNORING_9 ( .A(A[9]), .B(B[9]), .Y(L[9]) );
  XNOR_GATE_86 XNORING_10 ( .A(A[10]), .B(B[10]), .Y(L[10]) );
  XNOR_GATE_85 XNORING_11 ( .A(A[11]), .B(B[11]), .Y(L[11]) );
  XNOR_GATE_84 XNORING_12 ( .A(A[12]), .B(B[12]), .Y(L[12]) );
  XNOR_GATE_83 XNORING_13 ( .A(A[13]), .B(B[13]), .Y(L[13]) );
  XNOR_GATE_82 XNORING_14 ( .A(A[14]), .B(B[14]), .Y(L[14]) );
  XNOR_GATE_81 XNORING_15 ( .A(A[15]), .B(B[15]), .Y(L[15]) );
  XNOR_GATE_80 XNORING_16 ( .A(A[16]), .B(B[16]), .Y(L[16]) );
  XNOR_GATE_79 XNORING_17 ( .A(A[17]), .B(B[17]), .Y(L[17]) );
  XNOR_GATE_78 XNORING_18 ( .A(A[18]), .B(B[18]), .Y(L[18]) );
  XNOR_GATE_77 XNORING_19 ( .A(A[19]), .B(B[19]), .Y(L[19]) );
  XNOR_GATE_76 XNORING_20 ( .A(A[20]), .B(B[20]), .Y(L[20]) );
  XNOR_GATE_75 XNORING_21 ( .A(A[21]), .B(B[21]), .Y(L[21]) );
  XNOR_GATE_74 XNORING_22 ( .A(A[22]), .B(B[22]), .Y(L[22]) );
  XNOR_GATE_73 XNORING_23 ( .A(A[23]), .B(B[23]), .Y(L[23]) );
  XNOR_GATE_72 XNORING_24 ( .A(A[24]), .B(B[24]), .Y(L[24]) );
  XNOR_GATE_71 XNORING_25 ( .A(A[25]), .B(B[25]), .Y(L[25]) );
  XNOR_GATE_70 XNORING_26 ( .A(A[26]), .B(B[26]), .Y(L[26]) );
  XNOR_GATE_69 XNORING_27 ( .A(A[27]), .B(B[27]), .Y(L[27]) );
  XNOR_GATE_68 XNORING_28 ( .A(A[28]), .B(B[28]), .Y(L[28]) );
  XNOR_GATE_67 XNORING_29 ( .A(A[29]), .B(B[29]), .Y(L[29]) );
  XNOR_GATE_66 XNORING_30 ( .A(A[30]), .B(B[30]), .Y(L[30]) );
  XNOR_GATE_65 XNORING_31 ( .A(A[31]), .B(B[31]), .Y(L[31]) );
  N_AND_N32_3 ANDING ( .A(L), .Y(Y) );
endmodule


module EQU_COMPARATOR_N32_2 ( A, B, Y );
  input [31:0] A;
  input [31:0] B;
  output Y;

  wire   [31:0] L;

  XNOR_GATE_64 XNORING_0 ( .A(A[0]), .B(B[0]), .Y(L[0]) );
  XNOR_GATE_63 XNORING_1 ( .A(A[1]), .B(B[1]), .Y(L[1]) );
  XNOR_GATE_62 XNORING_2 ( .A(A[2]), .B(B[2]), .Y(L[2]) );
  XNOR_GATE_61 XNORING_3 ( .A(A[3]), .B(B[3]), .Y(L[3]) );
  XNOR_GATE_60 XNORING_4 ( .A(A[4]), .B(B[4]), .Y(L[4]) );
  XNOR_GATE_59 XNORING_5 ( .A(A[5]), .B(B[5]), .Y(L[5]) );
  XNOR_GATE_58 XNORING_6 ( .A(A[6]), .B(B[6]), .Y(L[6]) );
  XNOR_GATE_57 XNORING_7 ( .A(A[7]), .B(B[7]), .Y(L[7]) );
  XNOR_GATE_56 XNORING_8 ( .A(A[8]), .B(B[8]), .Y(L[8]) );
  XNOR_GATE_55 XNORING_9 ( .A(A[9]), .B(B[9]), .Y(L[9]) );
  XNOR_GATE_54 XNORING_10 ( .A(A[10]), .B(B[10]), .Y(L[10]) );
  XNOR_GATE_53 XNORING_11 ( .A(A[11]), .B(B[11]), .Y(L[11]) );
  XNOR_GATE_52 XNORING_12 ( .A(A[12]), .B(B[12]), .Y(L[12]) );
  XNOR_GATE_51 XNORING_13 ( .A(A[13]), .B(B[13]), .Y(L[13]) );
  XNOR_GATE_50 XNORING_14 ( .A(A[14]), .B(B[14]), .Y(L[14]) );
  XNOR_GATE_49 XNORING_15 ( .A(A[15]), .B(B[15]), .Y(L[15]) );
  XNOR_GATE_48 XNORING_16 ( .A(A[16]), .B(B[16]), .Y(L[16]) );
  XNOR_GATE_47 XNORING_17 ( .A(A[17]), .B(B[17]), .Y(L[17]) );
  XNOR_GATE_46 XNORING_18 ( .A(A[18]), .B(B[18]), .Y(L[18]) );
  XNOR_GATE_45 XNORING_19 ( .A(A[19]), .B(B[19]), .Y(L[19]) );
  XNOR_GATE_44 XNORING_20 ( .A(A[20]), .B(B[20]), .Y(L[20]) );
  XNOR_GATE_43 XNORING_21 ( .A(A[21]), .B(B[21]), .Y(L[21]) );
  XNOR_GATE_42 XNORING_22 ( .A(A[22]), .B(B[22]), .Y(L[22]) );
  XNOR_GATE_41 XNORING_23 ( .A(A[23]), .B(B[23]), .Y(L[23]) );
  XNOR_GATE_40 XNORING_24 ( .A(A[24]), .B(B[24]), .Y(L[24]) );
  XNOR_GATE_39 XNORING_25 ( .A(A[25]), .B(B[25]), .Y(L[25]) );
  XNOR_GATE_38 XNORING_26 ( .A(A[26]), .B(B[26]), .Y(L[26]) );
  XNOR_GATE_37 XNORING_27 ( .A(A[27]), .B(B[27]), .Y(L[27]) );
  XNOR_GATE_36 XNORING_28 ( .A(A[28]), .B(B[28]), .Y(L[28]) );
  XNOR_GATE_35 XNORING_29 ( .A(A[29]), .B(B[29]), .Y(L[29]) );
  XNOR_GATE_34 XNORING_30 ( .A(A[30]), .B(B[30]), .Y(L[30]) );
  XNOR_GATE_33 XNORING_31 ( .A(A[31]), .B(B[31]), .Y(L[31]) );
  N_AND_N32_2 ANDING ( .A(L), .Y(Y) );
endmodule


module EQU_COMPARATOR_N32_1 ( A, B, Y );
  input [31:0] A;
  input [31:0] B;
  output Y;

  wire   [31:0] L;

  XNOR_GATE_32 XNORING_0 ( .A(A[0]), .B(B[0]), .Y(L[0]) );
  XNOR_GATE_31 XNORING_1 ( .A(A[1]), .B(B[1]), .Y(L[1]) );
  XNOR_GATE_30 XNORING_2 ( .A(A[2]), .B(B[2]), .Y(L[2]) );
  XNOR_GATE_29 XNORING_3 ( .A(A[3]), .B(B[3]), .Y(L[3]) );
  XNOR_GATE_28 XNORING_4 ( .A(A[4]), .B(B[4]), .Y(L[4]) );
  XNOR_GATE_27 XNORING_5 ( .A(A[5]), .B(B[5]), .Y(L[5]) );
  XNOR_GATE_26 XNORING_6 ( .A(A[6]), .B(B[6]), .Y(L[6]) );
  XNOR_GATE_25 XNORING_7 ( .A(A[7]), .B(B[7]), .Y(L[7]) );
  XNOR_GATE_24 XNORING_8 ( .A(A[8]), .B(B[8]), .Y(L[8]) );
  XNOR_GATE_23 XNORING_9 ( .A(A[9]), .B(B[9]), .Y(L[9]) );
  XNOR_GATE_22 XNORING_10 ( .A(A[10]), .B(B[10]), .Y(L[10]) );
  XNOR_GATE_21 XNORING_11 ( .A(A[11]), .B(B[11]), .Y(L[11]) );
  XNOR_GATE_20 XNORING_12 ( .A(A[12]), .B(B[12]), .Y(L[12]) );
  XNOR_GATE_19 XNORING_13 ( .A(A[13]), .B(B[13]), .Y(L[13]) );
  XNOR_GATE_18 XNORING_14 ( .A(A[14]), .B(B[14]), .Y(L[14]) );
  XNOR_GATE_17 XNORING_15 ( .A(A[15]), .B(B[15]), .Y(L[15]) );
  XNOR_GATE_16 XNORING_16 ( .A(A[16]), .B(B[16]), .Y(L[16]) );
  XNOR_GATE_15 XNORING_17 ( .A(A[17]), .B(B[17]), .Y(L[17]) );
  XNOR_GATE_14 XNORING_18 ( .A(A[18]), .B(B[18]), .Y(L[18]) );
  XNOR_GATE_13 XNORING_19 ( .A(A[19]), .B(B[19]), .Y(L[19]) );
  XNOR_GATE_12 XNORING_20 ( .A(A[20]), .B(B[20]), .Y(L[20]) );
  XNOR_GATE_11 XNORING_21 ( .A(A[21]), .B(B[21]), .Y(L[21]) );
  XNOR_GATE_10 XNORING_22 ( .A(A[22]), .B(B[22]), .Y(L[22]) );
  XNOR_GATE_9 XNORING_23 ( .A(A[23]), .B(B[23]), .Y(L[23]) );
  XNOR_GATE_8 XNORING_24 ( .A(A[24]), .B(B[24]), .Y(L[24]) );
  XNOR_GATE_7 XNORING_25 ( .A(A[25]), .B(B[25]), .Y(L[25]) );
  XNOR_GATE_6 XNORING_26 ( .A(A[26]), .B(B[26]), .Y(L[26]) );
  XNOR_GATE_5 XNORING_27 ( .A(A[27]), .B(B[27]), .Y(L[27]) );
  XNOR_GATE_4 XNORING_28 ( .A(A[28]), .B(B[28]), .Y(L[28]) );
  XNOR_GATE_3 XNORING_29 ( .A(A[29]), .B(B[29]), .Y(L[29]) );
  XNOR_GATE_2 XNORING_30 ( .A(A[30]), .B(B[30]), .Y(L[30]) );
  XNOR_GATE_1 XNORING_31 ( .A(A[31]), .B(B[31]), .Y(L[31]) );
  N_AND_N32_1 ANDING ( .A(L), .Y(Y) );
endmodule


module NAND_GATE_1613 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1612 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1611 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1610 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1609 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1608 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1607 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1606 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1605 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1604 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1603 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1602 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1601 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1600 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1599 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1598 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1597 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1596 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1595 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1594 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1593 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1592 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1591 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1590 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1589 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1588 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1587 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1586 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1585 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1584 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1583 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1582 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1581 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1580 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1579 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1578 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1577 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1576 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1575 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1574 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1573 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1572 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1571 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1570 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1569 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1568 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1567 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1566 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1565 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1564 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1563 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1562 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1561 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1560 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1559 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1558 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1557 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1556 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1555 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1554 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1553 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1552 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1551 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1550 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1549 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1548 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1547 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1546 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1545 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1544 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1543 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1542 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1541 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1540 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1539 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1538 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1537 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1536 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1535 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1534 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1533 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1532 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1531 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1530 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1529 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1528 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1527 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1526 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module NAND_GATE_1525 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module NAND_GATE_1524 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1523 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module NAND_GATE_1522 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module NAND_GATE_1521 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1520 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module NAND_GATE_1519 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module NAND_GATE_1518 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1517 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1516 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1515 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1514 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1513 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1512 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1511 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1510 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1509 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1508 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1507 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1506 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1505 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1504 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1503 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1502 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1501 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1500 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1499 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1498 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1497 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1496 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1495 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1494 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1493 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1492 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1491 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1490 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1489 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1488 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1487 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1486 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1485 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1484 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1483 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1482 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1481 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1480 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1479 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1478 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1477 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1476 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1475 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1474 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1473 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1472 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1471 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1470 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1469 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1468 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1467 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1466 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1465 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1464 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1463 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1462 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1461 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1460 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1459 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1458 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1457 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1456 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1455 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1454 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1453 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1452 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1451 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1450 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1449 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1448 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1447 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1446 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1445 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1444 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1443 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1442 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1441 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1440 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1439 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1438 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1437 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1436 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1435 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1434 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1433 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1432 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1431 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1430 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module NAND_GATE_1429 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module NAND_GATE_1428 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1427 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module NAND_GATE_1426 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module NAND_GATE_1425 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1424 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module NAND_GATE_1423 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1422 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1421 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1420 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1419 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1418 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1417 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1416 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1415 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1414 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1413 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1412 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1411 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1410 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1409 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1408 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1407 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1406 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1405 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1404 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1403 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1402 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1401 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1400 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1399 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1398 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1397 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1396 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1395 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1394 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1393 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1392 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1391 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1390 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1389 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1388 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1387 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1386 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1385 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1384 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1383 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1382 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1381 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1380 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1379 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1378 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1377 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1376 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1375 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1374 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1373 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1372 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1371 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1370 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1369 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1368 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1367 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1366 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1365 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1364 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1363 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1362 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1361 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1360 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1359 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1358 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1357 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1356 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1355 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1354 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1353 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1352 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1351 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1350 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1349 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1348 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1347 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1346 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1345 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1344 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1343 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1342 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1341 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1340 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1339 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1338 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1337 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1336 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1335 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1334 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module NAND_GATE_1333 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module NAND_GATE_1332 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1331 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module NAND_GATE_1330 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module NAND_GATE_1329 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1328 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module NAND_GATE_1327 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1326 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1325 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1324 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1323 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1322 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1321 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1320 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1319 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1318 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1317 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1316 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1315 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1314 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1313 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1312 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1311 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1310 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1309 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1308 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1307 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1306 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1305 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1304 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1303 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1302 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1301 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1300 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1299 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1298 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1297 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1296 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1295 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1294 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1293 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1292 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1291 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1290 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1289 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1288 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1287 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1286 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1285 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1284 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1283 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1282 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1281 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1280 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1279 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1278 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1277 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1276 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1275 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1274 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1273 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1272 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1271 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1270 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1269 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1268 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1267 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1266 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1265 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1264 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1263 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1262 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1261 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1260 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1259 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1258 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1257 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1256 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1255 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1254 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1253 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1252 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1251 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1250 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1249 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1248 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1247 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1246 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1245 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1244 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1243 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1242 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1241 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1240 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1239 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1238 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1237 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1236 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1235 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1234 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1233 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1232 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1231 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1230 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1229 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1228 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1227 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1226 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1225 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1224 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1223 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1222 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1221 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1220 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1219 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1218 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1217 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1216 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1215 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1214 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1213 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1212 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1211 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1210 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1209 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1208 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1207 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1206 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1205 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1204 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1203 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1202 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1201 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1200 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1199 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1198 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1197 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1196 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1195 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1194 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1193 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1192 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1191 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1190 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1189 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1188 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1187 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1186 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1185 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1184 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1183 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1182 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1181 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1180 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1179 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1178 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1177 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1176 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1175 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1174 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1173 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1172 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1171 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1170 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1169 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1168 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1167 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1166 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1165 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1164 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1163 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1162 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1161 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1160 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1159 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1158 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1157 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1156 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1155 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1154 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1153 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1152 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1151 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1150 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1149 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1148 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1147 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1146 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1145 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1144 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1143 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1142 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1141 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1140 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1139 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1138 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1137 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1136 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1135 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1134 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1133 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1132 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1131 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1130 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1129 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1128 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1127 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1126 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1125 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1124 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1123 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1122 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1121 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1120 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1119 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1118 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1117 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1116 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1115 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1114 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1113 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1112 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1111 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1110 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1109 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1108 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1107 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1106 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1105 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1104 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1103 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1102 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1101 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1100 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1099 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1098 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1097 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1096 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1095 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1094 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1093 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1092 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1091 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1090 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1089 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1088 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1087 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1086 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1085 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1084 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1083 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1082 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1081 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1080 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1079 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1078 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1077 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1076 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1075 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1074 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1073 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1072 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1071 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1070 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1069 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1068 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1067 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1066 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1065 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1064 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1063 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1062 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1061 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1060 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1059 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1058 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1057 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1056 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1055 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1054 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1053 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1052 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1051 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1050 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1049 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1048 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1047 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1046 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1045 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1044 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1043 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1042 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1041 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1040 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1039 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1038 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1037 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1036 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1035 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1034 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1033 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1032 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1031 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1030 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1029 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1028 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1027 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1026 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1025 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1024 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1023 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1022 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1021 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1020 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1019 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1018 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1017 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1016 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1015 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1014 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1013 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1012 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1011 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1010 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1009 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1008 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1007 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1006 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1005 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1004 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1003 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1002 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1001 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1000 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_999 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_998 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_997 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_996 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_995 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_994 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_993 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_992 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_991 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_990 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_989 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_988 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_987 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_986 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_985 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_984 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_983 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_982 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_981 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_980 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_979 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_978 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_977 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_976 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_975 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_974 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_973 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_972 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_971 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_970 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_969 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_968 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_967 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_966 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_965 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_964 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_963 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_962 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_961 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_960 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_959 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_958 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_957 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_956 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_955 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_954 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_953 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_952 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_951 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_950 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_949 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_948 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_947 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_946 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_945 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_944 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_943 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_942 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_941 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_940 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_939 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_938 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_937 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_936 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_935 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_934 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_933 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_932 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_931 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_930 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_929 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_928 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_927 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_926 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_925 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_924 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_923 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_922 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_921 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_920 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_919 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_918 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_917 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_916 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_915 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_914 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_913 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_912 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_911 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_910 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_909 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_908 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_907 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_906 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_905 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_904 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_903 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_902 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_901 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_900 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_899 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_898 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_897 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_896 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_895 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_894 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_893 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_892 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_891 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_890 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_889 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_888 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_887 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_886 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_885 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_884 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_883 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_882 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_881 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_880 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_879 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_878 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_877 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_876 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_875 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_874 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_873 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_872 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_871 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_870 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_869 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_868 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_867 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_866 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_865 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_864 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_863 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_862 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_861 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_860 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_859 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_858 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_857 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_856 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_855 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_854 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_853 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_852 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_851 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_850 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_849 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_848 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_847 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_846 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_845 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_844 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_843 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_842 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_841 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_840 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_839 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_838 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_837 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_836 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_835 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_834 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_833 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_832 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_831 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_830 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_829 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_828 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_827 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_826 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_825 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_824 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_823 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_822 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_821 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_820 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_819 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_818 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_817 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_816 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_815 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_814 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_813 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_812 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_811 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_810 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_809 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_808 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_807 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_806 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_805 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_804 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_803 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_802 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_801 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_800 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_799 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_798 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_797 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_796 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_795 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_794 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_793 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_792 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_791 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_790 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_789 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_788 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_787 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_786 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_785 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_784 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_783 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_782 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_781 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_780 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_779 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_778 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_777 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_776 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_775 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_774 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_773 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_772 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_771 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_770 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_769 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_768 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_767 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_766 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_765 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_764 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_763 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_762 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_761 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_760 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_759 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_758 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_757 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_756 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_755 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_754 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_753 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_752 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_751 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_750 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_749 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_748 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_747 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_746 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_745 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_744 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_743 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_742 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_741 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_740 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_739 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_738 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_737 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_736 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_735 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_734 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_733 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_732 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_731 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_730 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_729 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_728 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_727 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_726 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_725 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_724 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_723 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_722 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_721 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_720 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_719 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_718 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_717 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_716 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_715 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_714 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_713 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_712 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_711 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_710 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_709 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_708 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_707 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_706 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_705 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_704 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_703 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_702 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_701 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_700 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_699 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_698 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_697 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_696 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_695 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_694 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_693 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_692 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_691 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_690 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_689 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_688 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_687 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_686 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_685 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_684 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_683 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_682 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_681 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_680 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_679 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_678 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_677 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_676 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_675 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_674 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_673 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_672 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_671 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_670 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_669 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_668 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_667 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_666 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_665 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_664 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_663 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_662 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_661 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_660 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_659 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_658 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_657 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_656 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_655 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_654 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_653 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_652 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_651 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_650 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_649 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_648 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_647 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_646 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_645 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_644 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_643 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_642 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_641 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_640 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_639 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_638 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_637 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_636 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_635 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_634 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_633 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_632 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_631 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_630 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_629 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_628 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_627 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_626 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_625 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_624 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_623 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_622 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_621 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_620 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_619 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_618 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_617 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_616 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_615 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_614 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_613 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_612 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_611 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_610 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_609 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_608 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_607 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_606 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_605 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_604 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_603 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_602 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_601 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_600 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_599 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_598 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_597 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_596 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_595 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_594 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_593 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_592 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_591 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_590 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_589 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_588 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_587 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_586 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_585 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_584 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_583 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_582 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_581 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_580 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_579 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_578 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_577 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_576 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_575 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_574 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_573 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_572 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_571 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_570 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_569 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_568 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_567 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_566 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_565 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_564 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_563 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_562 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_561 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_560 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_559 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_558 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_557 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_556 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_555 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_554 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_553 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_552 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_551 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_550 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_549 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_548 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_547 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_546 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_545 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_544 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_543 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_542 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_541 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_540 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_539 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_538 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_537 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_536 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_535 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_534 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_533 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_532 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_531 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_530 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_529 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_528 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_527 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_526 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_525 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_524 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_523 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_522 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_521 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_520 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_519 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_518 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_517 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_516 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_515 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_514 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_513 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_512 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_511 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_510 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_509 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_508 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_507 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_506 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_505 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_504 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_503 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_502 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_501 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_500 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_499 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_498 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_497 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_496 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_495 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_494 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_493 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_492 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_491 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_490 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_489 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_488 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_487 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_486 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_485 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_484 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_483 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_482 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_481 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_480 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_479 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_478 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_477 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_476 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_475 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_474 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_473 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_472 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_471 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_470 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_469 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_468 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_467 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_466 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_465 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_464 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_463 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_462 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_461 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_460 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_459 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_458 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_457 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_456 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_455 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_454 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_453 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_452 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_451 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_450 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_449 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_448 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_447 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_446 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_445 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_444 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_443 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_442 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_441 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_440 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_439 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_438 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_437 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_436 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_435 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_434 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_433 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_432 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_431 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_430 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_429 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_428 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_427 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_426 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_425 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_424 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_423 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_422 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_421 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_420 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_419 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_418 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_417 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_416 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_415 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_414 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_413 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_412 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_411 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_410 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_409 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_408 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_407 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_406 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_405 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_404 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_403 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_402 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_401 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_400 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_399 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_398 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_397 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_396 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_395 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_394 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_393 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_392 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_391 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_390 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_389 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_388 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_387 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_386 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_385 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_384 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_383 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_382 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_381 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_380 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_379 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_378 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_377 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_376 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_375 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_374 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_373 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_372 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_371 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_370 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_369 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_368 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_367 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_366 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_365 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_364 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_363 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_362 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_361 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_360 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_359 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_358 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_357 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_356 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_355 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_354 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_353 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_352 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_351 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_350 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_349 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_348 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_347 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_346 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_345 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_344 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_343 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_342 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_341 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_340 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_339 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_338 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_337 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_336 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_335 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_334 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_333 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_332 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_331 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_330 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_329 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_328 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_327 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_326 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_325 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_324 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_323 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_322 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_321 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_320 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_319 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_318 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_317 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_316 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_315 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_314 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_313 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_312 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_311 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_310 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_309 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_308 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_307 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_306 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_305 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_304 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_303 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_302 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_301 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_300 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_299 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_298 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_297 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_296 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_295 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_294 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_293 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_292 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_291 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_290 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_289 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_288 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_287 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_286 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_285 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_284 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_283 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_282 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_281 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_280 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_279 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_278 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_277 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_276 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_275 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_274 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_273 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_272 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_271 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_270 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_269 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_268 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_267 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_266 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_265 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_264 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_263 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_262 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_261 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_260 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_259 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_258 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_257 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_256 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_255 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_254 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_253 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_252 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_251 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_250 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_249 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_248 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_247 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_246 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_245 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_244 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_243 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_242 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_241 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_240 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_239 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_238 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_237 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_236 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_235 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_234 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_233 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_232 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_231 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_230 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_229 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_228 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_227 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_226 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_225 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_224 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_223 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_222 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_221 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_220 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_219 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_218 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_217 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_216 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_215 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_214 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_213 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_212 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_211 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_210 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_209 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_208 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_207 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_206 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_205 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_204 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_203 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_202 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_201 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_200 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_199 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_198 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_197 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_196 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_195 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_194 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_193 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_192 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_191 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_190 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_189 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_188 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_187 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_186 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_185 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_184 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_183 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_182 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_181 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_180 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_179 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_178 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_177 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_176 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_175 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_174 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_173 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_172 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_171 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_170 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_169 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_168 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_167 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_166 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_165 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_164 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_163 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_162 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_161 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_160 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_159 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_158 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_157 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_156 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_155 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_154 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_153 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_152 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_151 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_150 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_149 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_148 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_147 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_146 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_145 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_144 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_143 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_142 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_141 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_140 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_139 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_138 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_137 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_136 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_135 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_134 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_133 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_132 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_131 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_130 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_129 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_128 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_127 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_126 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_125 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_124 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_123 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_122 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_121 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_120 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_119 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_118 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_117 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_116 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_115 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_114 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_113 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_112 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_111 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_110 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_109 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_108 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_107 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_106 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_105 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_104 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_103 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_102 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_101 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_100 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_99 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_98 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_97 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_96 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_95 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_94 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_93 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_92 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_91 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_90 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_89 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_88 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_87 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_86 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_85 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_84 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_83 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_82 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_81 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_80 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_79 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_78 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_77 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_76 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_75 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_74 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_73 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_72 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_71 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_70 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_69 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_68 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_67 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_66 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_65 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_64 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_63 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_62 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_61 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_60 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_59 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_58 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_57 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_56 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_55 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_54 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_53 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_52 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_51 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_50 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_49 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_48 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_47 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_46 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_45 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_44 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_43 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_42 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_41 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_40 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_39 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_38 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_37 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_36 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_35 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_34 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_33 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_32 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_31 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_30 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_29 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_28 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_27 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_26 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_25 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_24 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_23 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_22 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_21 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_20 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_19 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_18 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_17 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_16 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_15 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_14 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_13 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_12 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_11 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_10 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_9 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_8 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_7 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_6 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_5 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_4 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_3 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_2 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module NAND_GATE_1 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module INV_1_127 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_126 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_125 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_124 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_123 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_122 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_121 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_120 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_119 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_118 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_117 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_116 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_115 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_114 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_113 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_112 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_111 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_110 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_109 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_108 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_107 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_106 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_105 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_104 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_103 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_102 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_101 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_100 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_99 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_98 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_97 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_96 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_95 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_94 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_93 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_92 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_91 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_90 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_89 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_88 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_87 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_86 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_85 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_84 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_83 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_82 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_81 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_80 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_79 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_78 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_77 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_76 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_75 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_74 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_73 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_72 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_71 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_70 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_69 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_68 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_67 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_66 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_65 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_64 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_63 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_62 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_61 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_60 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_59 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_58 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_57 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_56 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_55 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_54 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_53 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_52 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_51 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_50 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_49 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_48 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_47 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_46 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_45 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_44 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_43 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_42 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_41 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_40 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_39 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_38 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_37 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_36 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_35 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_34 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_33 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_32 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_31 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_30 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_29 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_28 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_27 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_26 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_25 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_24 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_23 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_22 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_21 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_20 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_19 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_18 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_17 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_16 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_15 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_14 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_13 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_12 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_11 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_10 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_9 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_8 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_7 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_6 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_5 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_4 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_3 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_2 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1_1 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module FA_297 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_635 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_634 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_700 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_699 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_337 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_296 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_633 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_632 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_698 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_697 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_336 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_295 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_631 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_630 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_696 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_695 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_335 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_294 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_629 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_628 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_694 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_693 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_334 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_293 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_627 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_626 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_692 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_691 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_333 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_292 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_625 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_624 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_690 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_689 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_332 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_291 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_623 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_622 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_688 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_687 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_331 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_290 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_621 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_620 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_686 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_685 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_330 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_289 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_619 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_618 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_684 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_683 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_329 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_288 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_617 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_616 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_682 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_681 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_328 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_287 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_615 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_614 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_680 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_679 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_327 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_286 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_613 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_612 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_678 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_677 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_326 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_285 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_611 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_610 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_676 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_675 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_325 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_284 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_609 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_608 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_674 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_673 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_324 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_283 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_607 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_606 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_672 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_671 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_323 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_282 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_605 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_604 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_670 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_669 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_322 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_281 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_603 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_602 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_668 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_667 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_321 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_280 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_601 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_600 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_666 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_665 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_320 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_279 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_599 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_598 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_664 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_663 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_319 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_278 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_597 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_596 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_662 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_661 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_318 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_277 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_595 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_594 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_660 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_659 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_317 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_276 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_593 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_592 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_658 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_657 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_316 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_275 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_591 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_590 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_656 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_655 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_315 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_274 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_589 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_588 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_654 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_653 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_314 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_273 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_587 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_586 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_652 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_651 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_313 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_272 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_585 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_584 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_650 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_649 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_312 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_271 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_583 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_582 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_648 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_647 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_311 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_270 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_581 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_580 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_646 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_645 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_310 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_269 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_579 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_578 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_642 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_641 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_306 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_268 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_577 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_576 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_640 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_639 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_305 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_267 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_575 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_574 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_638 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_637 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_304 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_266 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_573 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_572 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_636 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_635 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_303 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_265 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_571 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_570 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_634 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_633 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_302 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_264 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_569 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_568 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_632 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_631 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_301 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_263 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_567 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_566 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_630 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_629 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_300 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_262 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_565 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_564 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_628 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_627 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_299 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_261 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_563 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_562 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_626 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_625 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_298 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_260 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_561 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_560 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_624 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_623 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_297 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_259 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_559 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_558 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_622 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_621 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_296 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_258 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_557 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_556 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_620 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_619 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_295 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_257 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_555 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_554 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_618 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_617 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_294 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_256 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_553 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_552 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_616 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_615 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_293 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_255 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_551 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_550 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_614 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_613 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_292 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_254 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_549 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_548 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_612 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_611 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_291 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_253 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_547 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_546 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_610 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_609 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_290 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_252 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_545 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_544 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_608 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_607 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_289 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_251 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_543 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_542 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_606 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_605 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_288 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_250 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_541 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_540 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_604 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_603 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_287 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_249 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_539 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_538 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_602 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_601 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_286 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_248 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_537 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_536 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_600 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_599 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_285 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_247 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_535 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_534 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_598 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_597 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_284 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_246 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_533 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_532 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_596 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_595 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_283 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_245 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_531 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_530 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_594 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_593 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_282 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_244 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_529 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_528 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_592 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_591 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_281 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_243 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_527 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_526 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_590 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_589 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_280 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_242 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_525 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_524 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_588 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_587 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_279 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_241 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_523 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_522 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_586 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_585 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_278 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_240 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_521 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_520 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_584 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_583 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_277 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_239 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_519 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_518 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_582 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_581 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_276 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_238 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_517 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_516 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_580 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_579 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_275 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_237 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_515 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_514 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_578 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_577 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_274 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_236 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_513 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_512 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_576 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_575 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_273 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_235 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_511 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_510 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_574 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_573 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_272 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_234 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_509 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_508 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_572 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_571 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_271 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_233 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_507 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_506 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_570 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_569 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_270 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_232 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_505 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_504 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_568 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_567 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_269 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_231 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_503 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_502 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_566 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_565 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_268 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_230 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_501 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_500 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_564 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_563 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_267 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_229 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_499 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_498 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_562 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_561 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_266 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_228 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_497 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_496 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_560 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_559 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_265 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_227 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_495 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_494 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_558 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_557 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_264 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_226 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_493 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_492 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_556 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_555 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_263 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_225 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_491 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_490 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_554 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_553 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_262 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_224 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_489 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_488 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_552 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_551 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_261 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_223 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_487 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_486 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_550 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_549 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_260 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_222 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_485 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_484 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_548 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_547 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_259 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_221 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_483 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_482 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_546 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_545 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_258 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_220 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_481 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_480 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_544 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_543 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_257 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_219 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_479 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_478 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_542 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_541 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_256 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_218 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_477 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_476 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_540 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_539 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_255 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_217 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_475 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_474 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_538 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_537 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_254 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_216 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_473 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_472 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_536 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_535 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_253 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_215 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_471 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_470 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_534 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_533 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_252 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_214 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_469 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_468 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_532 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_531 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_251 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_213 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_467 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_466 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_530 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_529 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_250 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_212 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_465 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_464 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_528 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_527 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_249 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_211 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_463 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_462 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_526 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_525 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_248 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_210 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_461 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_460 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_524 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_523 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_247 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_209 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_459 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_458 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_522 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_521 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_246 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_208 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_457 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_456 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_520 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_519 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_245 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_207 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_455 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_454 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_518 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_517 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_244 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_206 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_453 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_452 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_516 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_515 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_243 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_205 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1, n2;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_417 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_416 XOR_GATE_2 ( .A(n2), .B(Ci), .Y(S) );
  AND_GATE_1_472 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_471 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_233 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  INV_X1 U1 ( .A(OUT_XOR), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(n2) );
endmodule


module FA_204 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_415 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_414 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_470 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_469 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_232 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_203 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_413 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_412 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_468 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_467 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_231 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_202 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_411 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_410 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_466 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_465 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_230 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_201 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_409 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_408 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_464 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_463 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_229 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_200 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_407 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_406 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_462 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_461 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_228 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_199 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_405 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_404 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_460 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_459 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_227 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_198 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_403 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_402 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_458 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_457 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_226 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_197 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_401 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_400 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_456 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_455 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_225 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_196 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_399 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_398 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_454 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_453 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_224 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_195 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_397 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_396 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_452 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_451 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_223 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_194 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_395 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_394 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_450 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_449 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_222 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_193 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_393 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_392 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_448 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_447 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_221 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_192 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_391 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_390 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_446 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_445 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_220 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_191 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_389 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_388 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_444 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_443 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_219 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_190 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_386 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_385 XOR_GATE_2 ( .A(n1), .B(Ci), .Y(S) );
  AND_GATE_1_386 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_385 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_190 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(OUT_XOR), .Z(n1) );
endmodule


module FA_189 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_384 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_383 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_384 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_383 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_189 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_188 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_382 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_381 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_382 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_381 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_188 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_187 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_380 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_379 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_380 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_379 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_187 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_186 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_378 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_377 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_378 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_377 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_186 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_185 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_376 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_375 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_376 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_375 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_185 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_184 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_374 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_373 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_374 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_373 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_184 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_183 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_372 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_371 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_372 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_371 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_183 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_182 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_370 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_369 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_370 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_369 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_182 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_181 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_368 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_367 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_368 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_367 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_181 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_180 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_366 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_365 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_366 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_365 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_180 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_179 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_364 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_363 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_364 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_363 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_179 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_178 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_362 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_361 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_362 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_361 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_178 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_177 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1, n2;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_360 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_359 XOR_GATE_2 ( .A(n2), .B(Ci), .Y(S) );
  AND_GATE_1_360 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_359 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_177 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  INV_X1 U1 ( .A(OUT_XOR), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(n2) );
endmodule


module FA_176 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_358 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_357 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_358 AND_GATE_1 ( .A(n1), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_357 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_176 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(A), .Z(n1) );
endmodule


module FA_175 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_356 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_355 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_356 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_355 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_175 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_174 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_354 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_353 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_354 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_353 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_174 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_173 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_352 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_351 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_352 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_351 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_173 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_172 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_349 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_348 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_349 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_348 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_172 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_171 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_347 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_346 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_347 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_346 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_171 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_170 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_345 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_344 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_345 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_344 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_170 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_169 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_343 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_342 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_343 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_342 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_169 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_168 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_341 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_340 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_341 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_340 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_168 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_167 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_339 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_338 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_339 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_338 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_167 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_166 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_337 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_336 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_337 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_336 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_166 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_165 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_335 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_334 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_335 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_334 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_165 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_164 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_333 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_332 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_333 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_332 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_164 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_163 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_331 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_330 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_331 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_330 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_163 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_162 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_329 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_328 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_329 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_328 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_162 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_161 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_327 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_326 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_327 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_326 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_161 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_160 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_325 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_324 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_325 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_324 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_160 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_159 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_323 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_322 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_323 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_322 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_159 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_158 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1, n2;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_321 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_320 XOR_GATE_2 ( .A(n1), .B(Ci), .Y(S) );
  AND_GATE_1_321 AND_GATE_1 ( .A(n2), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_320 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_158 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(OUT_XOR), .Z(n1) );
  CLKBUF_X1 U2 ( .A(A), .Z(n2) );
endmodule


module FA_157 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_319 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_318 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_319 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_318 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_157 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_156 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_317 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_316 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_317 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_316 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_156 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_155 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_315 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_314 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_315 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_314 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_155 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_154 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1, n2;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_312 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_311 XOR_GATE_2 ( .A(n2), .B(Ci), .Y(S) );
  AND_GATE_1_312 AND_GATE_1 ( .A(A), .B(n1), .Y(OUT_AND[0]) );
  AND_GATE_1_311 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_154 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(B), .Z(n1) );
  CLKBUF_X1 U2 ( .A(OUT_XOR), .Z(n2) );
endmodule


module FA_153 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1, n2;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_310 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_309 XOR_GATE_2 ( .A(OUT_XOR), .B(n2), .Y(S) );
  AND_GATE_1_310 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_309 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_153 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  INV_X1 U1 ( .A(Ci), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(n2) );
endmodule


module FA_152 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_308 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_307 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_308 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_307 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_152 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_151 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_306 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_305 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_306 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_305 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_151 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_150 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_304 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_303 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_304 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_303 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_150 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_149 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_302 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_301 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_302 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_301 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_149 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_148 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_300 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_299 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_300 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_299 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_148 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_147 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_298 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_297 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_298 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_297 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_147 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_146 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_296 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_295 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_296 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_295 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_146 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_145 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_294 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_293 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_294 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_293 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_145 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_144 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_292 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_291 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_292 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_291 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_144 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_143 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_290 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_289 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_290 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_289 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_143 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_142 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_288 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_287 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_288 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_287 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_142 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_141 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_286 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_285 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_286 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_285 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_141 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_140 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_284 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_283 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_284 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_283 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_140 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_139 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_282 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_281 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_282 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_281 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_139 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_138 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_280 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_279 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_280 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_279 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_138 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_137 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_278 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_277 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_278 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_277 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_137 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_136 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_275 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_274 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_275 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_274 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_136 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_135 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_273 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_272 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_273 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_272 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_135 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_134 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_271 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_270 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_271 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_270 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_134 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_133 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_269 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_268 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_269 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_268 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_133 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_132 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_267 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_266 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_267 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_266 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_132 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_131 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_265 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_264 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_265 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_264 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_131 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_130 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_263 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_262 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_263 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_262 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_130 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_129 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_261 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_260 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_261 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_260 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_129 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_128 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_259 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_258 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_259 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_258 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_128 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_127 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_257 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_256 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_257 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_256 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_127 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_126 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_255 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_254 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_255 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_254 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_126 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_125 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_253 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_252 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_253 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_252 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_125 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_124 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_251 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_250 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_251 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_250 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_124 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_123 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_249 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_248 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_249 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_248 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_123 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_122 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_247 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_246 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_247 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_246 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_122 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_121 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_245 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_244 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_245 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_244 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_121 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_120 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_243 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_242 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_243 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_242 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_120 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_119 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_241 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_240 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_241 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_240 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_119 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_118 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_238 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_237 XOR_GATE_2 ( .A(n1), .B(Ci), .Y(S) );
  AND_GATE_1_238 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_237 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_118 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(OUT_XOR), .Z(n1) );
endmodule


module FA_117 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_236 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_235 XOR_GATE_2 ( .A(n1), .B(Ci), .Y(S) );
  AND_GATE_1_236 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_235 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_117 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(OUT_XOR), .Z(n1) );
endmodule


module FA_116 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1, n2;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_234 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_233 XOR_GATE_2 ( .A(n2), .B(Ci), .Y(S) );
  AND_GATE_1_234 AND_GATE_1 ( .A(n1), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_233 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_116 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(A), .Z(n1) );
  CLKBUF_X1 U2 ( .A(OUT_XOR), .Z(n2) );
endmodule


module FA_115 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_232 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_231 XOR_GATE_2 ( .A(OUT_XOR), .B(n1), .Y(S) );
  AND_GATE_1_232 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_231 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_115 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n1) );
endmodule


module FA_114 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_230 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_229 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_230 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_229 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_114 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_113 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_228 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_227 XOR_GATE_2 ( .A(OUT_XOR), .B(n1), .Y(S) );
  AND_GATE_1_228 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_227 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_113 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n1) );
endmodule


module FA_112 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_226 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_225 XOR_GATE_2 ( .A(OUT_XOR), .B(n1), .Y(S) );
  AND_GATE_1_226 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_225 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_112 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n1) );
endmodule


module FA_111 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1, n2;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_224 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_223 XOR_GATE_2 ( .A(n1), .B(n2), .Y(S) );
  AND_GATE_1_224 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_223 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_111 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(OUT_XOR), .Z(n1) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n2) );
endmodule


module FA_110 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1, n2;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_222 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_221 XOR_GATE_2 ( .A(n1), .B(n2), .Y(S) );
  AND_GATE_1_222 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_221 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_110 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(OUT_XOR), .Z(n1) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n2) );
endmodule


module FA_109 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1, n2;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_220 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_219 XOR_GATE_2 ( .A(n1), .B(n2), .Y(S) );
  AND_GATE_1_220 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_219 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_109 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(OUT_XOR), .Z(n1) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n2) );
endmodule


module FA_108 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1, n2, n3;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_218 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_217 XOR_GATE_2 ( .A(n3), .B(n2), .Y(S) );
  AND_GATE_1_218 AND_GATE_1 ( .A(n1), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_217 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_108 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(A), .Z(n1) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n2) );
  CLKBUF_X1 U3 ( .A(OUT_XOR), .Z(n3) );
endmodule


module FA_107 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_216 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_215 XOR_GATE_2 ( .A(OUT_XOR), .B(n1), .Y(S) );
  AND_GATE_1_216 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_215 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_107 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n1) );
endmodule


module FA_106 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_214 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_213 XOR_GATE_2 ( .A(OUT_XOR), .B(n1), .Y(S) );
  AND_GATE_1_214 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_213 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_106 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(Ci), .Z(n1) );
endmodule


module FA_105 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1, n2, n3;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_212 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_211 XOR_GATE_2 ( .A(n2), .B(n3), .Y(S) );
  AND_GATE_1_212 AND_GATE_1 ( .A(n1), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_211 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_105 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(A), .Z(n1) );
  CLKBUF_X1 U2 ( .A(OUT_XOR), .Z(n2) );
  CLKBUF_X1 U3 ( .A(Ci), .Z(n3) );
endmodule


module FA_104 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1, n2, n3;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_210 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_209 XOR_GATE_2 ( .A(n1), .B(n3), .Y(S) );
  AND_GATE_1_210 AND_GATE_1 ( .A(n2), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_209 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_104 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(OUT_XOR), .Z(n1) );
  CLKBUF_X1 U2 ( .A(A), .Z(n2) );
  CLKBUF_X1 U3 ( .A(Ci), .Z(n3) );
endmodule


module FA_103 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1, n2, n3;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_208 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_207 XOR_GATE_2 ( .A(n2), .B(n3), .Y(S) );
  AND_GATE_1_208 AND_GATE_1 ( .A(n1), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_207 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_103 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(A), .Z(n1) );
  CLKBUF_X1 U2 ( .A(OUT_XOR), .Z(n2) );
  CLKBUF_X1 U3 ( .A(Ci), .Z(n3) );
endmodule


module FA_102 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_206 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_205 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_206 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_205 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_102 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_101 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_204 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_203 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_204 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_203 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_101 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_100 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_201 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_200 XOR_GATE_2 ( .A(n1), .B(Ci), .Y(S) );
  AND_GATE_1_201 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_200 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_100 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(OUT_XOR), .Z(n1) );
endmodule


module FA_99 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_199 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_198 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_199 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_198 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_99 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_98 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_197 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_196 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_197 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_196 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_98 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_97 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_195 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_194 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_195 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_194 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_97 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_96 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_193 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_192 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_193 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_192 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_96 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_95 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_191 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_190 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_191 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_190 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_95 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_94 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_189 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_188 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_189 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_188 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_94 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_93 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_187 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_186 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_187 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_186 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_93 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_92 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_185 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_184 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_185 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_184 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_92 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_91 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_183 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_182 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_183 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_182 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_91 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_90 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_181 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_180 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_181 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_180 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_90 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_89 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_179 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_178 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_179 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_178 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_89 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_88 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_177 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_176 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_177 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_176 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_88 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_87 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_175 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_174 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_175 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_174 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_87 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_86 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_173 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_172 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_173 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_172 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_86 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_85 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_171 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_170 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_171 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_170 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_85 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_84 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_169 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_168 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_169 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_168 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_84 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_83 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_167 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_166 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_167 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_166 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_83 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_82 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1, n2;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_164 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_163 XOR_GATE_2 ( .A(n2), .B(Ci), .Y(S) );
  AND_GATE_1_164 AND_GATE_1 ( .A(n1), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_163 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_82 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(A), .Z(n1) );
  CLKBUF_X1 U2 ( .A(OUT_XOR), .Z(n2) );
endmodule


module FA_81 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_162 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_161 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_162 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_161 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_81 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_80 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1, n2;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_160 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_159 XOR_GATE_2 ( .A(n2), .B(Ci), .Y(S) );
  AND_GATE_1_160 AND_GATE_1 ( .A(n1), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_159 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_80 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(A), .Z(n1) );
  CLKBUF_X1 U2 ( .A(OUT_XOR), .Z(n2) );
endmodule


module FA_79 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_158 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_157 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_158 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_157 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_79 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_78 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_156 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_155 XOR_GATE_2 ( .A(n1), .B(Ci), .Y(S) );
  AND_GATE_1_156 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_155 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_78 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(OUT_XOR), .Z(n1) );
endmodule


module FA_77 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_154 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_153 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_154 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_153 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_77 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_76 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_152 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_151 XOR_GATE_2 ( .A(n1), .B(Ci), .Y(S) );
  AND_GATE_1_152 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_151 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_76 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(OUT_XOR), .Z(n1) );
endmodule


module FA_75 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_150 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_149 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_150 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_149 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_75 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_74 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_148 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_147 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_148 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_147 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_74 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_73 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_146 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_145 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_146 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_145 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_73 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_72 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_144 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_143 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_144 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_143 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_72 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_71 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_142 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_141 XOR_GATE_2 ( .A(n1), .B(Ci), .Y(S) );
  AND_GATE_1_142 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_141 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_71 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(OUT_XOR), .Z(n1) );
endmodule


module FA_70 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_140 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_139 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_140 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_139 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_70 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_69 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_138 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_137 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_138 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_137 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_69 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_68 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_136 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_135 XOR_GATE_2 ( .A(n1), .B(Ci), .Y(S) );
  AND_GATE_1_136 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_135 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_68 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(OUT_XOR), .Z(n1) );
endmodule


module FA_67 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_134 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_133 XOR_GATE_2 ( .A(n1), .B(Ci), .Y(S) );
  AND_GATE_1_134 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_133 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_67 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(OUT_XOR), .Z(n1) );
endmodule


module FA_66 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_132 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_131 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_132 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_131 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_66 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_65 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_130 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_129 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_130 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_129 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_65 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_64 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_128 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_127 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_128 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_127 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_64 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_63 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_126 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_125 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_126 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_125 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_63 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_62 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_124 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_123 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_124 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_123 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_62 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_61 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_122 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_121 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_122 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_121 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_61 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_60 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_120 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_119 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_120 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_119 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_60 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_59 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_118 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_117 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_118 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_117 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_59 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_58 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_116 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_115 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_116 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_115 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_58 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_57 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_114 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_113 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_114 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_113 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_57 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_56 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_112 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_111 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_112 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_111 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_56 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_55 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_110 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_109 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_110 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_109 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_55 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_54 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_108 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_107 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_108 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_107 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_54 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_53 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_106 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_105 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_106 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_105 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_53 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_52 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_104 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_103 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_104 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_103 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_52 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_51 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_102 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_101 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_102 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_101 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_51 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_50 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_100 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_99 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_100 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_99 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_50 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_49 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_98 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_97 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_98 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_97 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_49 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_48 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_96 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_95 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_96 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_95 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_48 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_47 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_94 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_93 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_94 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_93 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_47 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_46 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_92 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_91 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_92 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_91 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_46 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_45 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_90 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_89 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_90 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_89 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_45 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_44 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_88 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_87 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_88 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_87 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_44 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_43 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_86 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_85 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_86 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_85 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_43 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_42 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_84 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_83 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_84 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_83 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_42 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_41 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_82 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_81 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_82 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_81 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_41 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_40 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_80 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_79 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_80 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_79 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_40 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_39 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_78 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_77 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_78 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_77 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_39 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_38 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_76 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_75 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_76 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_75 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_38 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_37 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_74 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_73 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_74 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_73 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_37 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_36 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_72 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_71 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_72 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_71 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_36 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_35 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_70 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_69 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_70 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_69 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_35 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_34 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_68 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_67 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_68 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_67 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_34 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_33 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_66 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_65 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_66 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_65 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_33 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_32 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_64 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_63 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_64 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_63 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_32 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_31 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_62 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_61 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_62 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_61 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_31 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_30 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_60 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_59 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_60 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_59 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_30 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_29 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_58 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_57 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_58 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_57 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_29 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_28 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_56 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_55 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_56 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_55 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_28 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_27 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_54 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_53 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_54 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_53 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_27 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_26 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_52 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_51 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_52 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_51 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_26 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_25 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_50 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_49 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_50 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_49 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_25 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_24 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_48 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_47 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_48 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_47 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_24 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_23 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_46 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_45 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_46 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_45 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_23 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_22 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_44 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_43 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_44 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_43 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_22 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_21 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_42 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_41 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_42 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_41 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_21 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_20 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_40 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_39 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_40 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_39 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_20 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_19 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_38 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_37 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_38 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_37 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_19 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_18 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_36 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_35 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_36 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_35 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_18 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_17 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_34 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_33 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_34 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_33 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_17 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_16 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_32 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_31 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_32 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_31 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_16 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_15 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_30 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_29 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_30 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_29 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_15 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_14 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_28 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_27 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_28 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_27 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_14 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_13 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_26 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_25 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_26 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_25 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_13 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_12 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_24 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_23 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_24 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_23 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_12 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_11 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_22 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_21 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_22 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_21 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_11 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_10 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_20 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_19 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_20 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_19 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_10 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_9 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_18 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_17 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_18 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_17 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_9 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_8 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_16 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_15 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_16 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_15 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_8 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_7 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_14 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_13 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_14 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_13 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_7 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_6 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_12 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_11 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_12 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_11 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_6 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_5 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_10 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_9 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_10 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_9 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_5 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_4 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_8 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_7 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_8 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_7 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_4 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_3 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_6 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_5 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_6 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_5 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_3 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_2 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_4 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_3 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_4 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_3 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_2 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module FA_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_2 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_1 XOR_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(S) );
  AND_GATE_1_2 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_1 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_1 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
endmodule


module HA_8 ( A, B, S, Co );
  input A, B;
  output S, Co;


  XOR_GATE_1_418 XOR_GATE_INST ( .A(A), .B(B), .Y(S) );
  AND_GATE_1_473 AND_GATE_INST ( .A(A), .B(B), .Y(Co) );
endmodule


module HA_7 ( A, B, S, Co );
  input A, B;
  output S, Co;


  XOR_GATE_1_387 XOR_GATE_INST ( .A(A), .B(B), .Y(S) );
  AND_GATE_1_387 AND_GATE_INST ( .A(A), .B(B), .Y(Co) );
endmodule


module HA_6 ( A, B, S, Co );
  input A, B;
  output S, Co;


  XOR_GATE_1_350 XOR_GATE_INST ( .A(A), .B(B), .Y(S) );
  AND_GATE_1_350 AND_GATE_INST ( .A(A), .B(B), .Y(Co) );
endmodule


module HA_5 ( A, B, S, Co );
  input A, B;
  output S, Co;
  wire   n1;

  XOR_GATE_1_313 XOR_GATE_INST ( .A(A), .B(n1), .Y(S) );
  AND_GATE_1_313 AND_GATE_INST ( .A(A), .B(B), .Y(Co) );
  CLKBUF_X1 U1 ( .A(B), .Z(n1) );
endmodule


module HA_4 ( A, B, S, Co );
  input A, B;
  output S, Co;


  XOR_GATE_1_276 XOR_GATE_INST ( .A(A), .B(B), .Y(S) );
  AND_GATE_1_276 AND_GATE_INST ( .A(A), .B(B), .Y(Co) );
endmodule


module HA_3 ( A, B, S, Co );
  input A, B;
  output S, Co;


  XOR_GATE_1_239 XOR_GATE_INST ( .A(A), .B(B), .Y(S) );
  AND_GATE_1_239 AND_GATE_INST ( .A(A), .B(B), .Y(Co) );
endmodule


module HA_2 ( A, B, S, Co );
  input A, B;
  output S, Co;


  XOR_GATE_1_202 XOR_GATE_INST ( .A(A), .B(B), .Y(S) );
  AND_GATE_1_202 AND_GATE_INST ( .A(A), .B(B), .Y(Co) );
endmodule


module HA_1 ( A, B, S, Co );
  input A, B;
  output S, Co;


  XOR_GATE_1_165 XOR_GATE_INST ( .A(A), .B(B), .Y(S) );
  AND_GATE_1_165 AND_GATE_INST ( .A(A), .B(B), .Y(Co) );
endmodule


module REG_N6_2 ( D, Q, EN, RST, CLK );
  input [5:0] D;
  output [5:0] Q;
  input EN, RST, CLK;
  wire   n1;

  FD_1_109 FF_0 ( .D(D[0]), .CLK(CLK), .EN(n1), .RST(RST), .Q(Q[0]) );
  FD_1_108 FF_1 ( .D(D[1]), .CLK(CLK), .EN(n1), .RST(RST), .Q(Q[1]) );
  FD_1_107 FF_2 ( .D(D[2]), .CLK(CLK), .EN(n1), .RST(RST), .Q(Q[2]) );
  FD_1_106 FF_3 ( .D(D[3]), .CLK(CLK), .EN(n1), .RST(RST), .Q(Q[3]) );
  FD_1_105 FF_4 ( .D(D[4]), .CLK(CLK), .EN(n1), .RST(RST), .Q(Q[4]) );
  FD_1_104 FF_5 ( .D(D[5]), .CLK(CLK), .EN(n1), .RST(RST), .Q(Q[5]) );
  BUF_X1 U1 ( .A(EN), .Z(n1) );
endmodule


module REG_N6_1 ( D, Q, EN, RST, CLK );
  input [5:0] D;
  output [5:0] Q;
  input EN, RST, CLK;


  FD_1_103 FF_0 ( .D(D[0]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[0]) );
  FD_1_102 FF_1 ( .D(D[1]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[1]) );
  FD_1_101 FF_2 ( .D(D[2]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[2]) );
  FD_1_100 FF_3 ( .D(D[3]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[3]) );
  FD_1_99 FF_4 ( .D(D[4]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[4]) );
  FD_1_98 FF_5 ( .D(D[5]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[5]) );
endmodule


module EQU_COMPARATOR_N5_6 ( A, B, Y );
  input [4:0] A;
  input [4:0] B;
  output Y;

  wire   [4:0] L;

  XNOR_GATE_213 XNORING_0 ( .A(A[0]), .B(B[0]), .Y(L[0]) );
  XNOR_GATE_212 XNORING_1 ( .A(A[1]), .B(B[1]), .Y(L[1]) );
  XNOR_GATE_211 XNORING_2 ( .A(A[2]), .B(B[2]), .Y(L[2]) );
  XNOR_GATE_210 XNORING_3 ( .A(A[3]), .B(B[3]), .Y(L[3]) );
  XNOR_GATE_209 XNORING_4 ( .A(A[4]), .B(B[4]), .Y(L[4]) );
  N_AND_N5_6 ANDING ( .A(L), .Y(Y) );
endmodule


module EQU_COMPARATOR_N5_5 ( A, B, Y );
  input [4:0] A;
  input [4:0] B;
  output Y;

  wire   [4:0] L;

  XNOR_GATE_208 XNORING_0 ( .A(A[0]), .B(B[0]), .Y(L[0]) );
  XNOR_GATE_207 XNORING_1 ( .A(A[1]), .B(B[1]), .Y(L[1]) );
  XNOR_GATE_206 XNORING_2 ( .A(A[2]), .B(B[2]), .Y(L[2]) );
  XNOR_GATE_205 XNORING_3 ( .A(A[3]), .B(B[3]), .Y(L[3]) );
  XNOR_GATE_204 XNORING_4 ( .A(A[4]), .B(B[4]), .Y(L[4]) );
  N_AND_N5_5 ANDING ( .A(L), .Y(Y) );
endmodule


module EQU_COMPARATOR_N5_4 ( A, B, Y );
  input [4:0] A;
  input [4:0] B;
  output Y;

  wire   [4:0] L;

  XNOR_GATE_203 XNORING_0 ( .A(A[0]), .B(B[0]), .Y(L[0]) );
  XNOR_GATE_202 XNORING_1 ( .A(A[1]), .B(B[1]), .Y(L[1]) );
  XNOR_GATE_201 XNORING_2 ( .A(A[2]), .B(B[2]), .Y(L[2]) );
  XNOR_GATE_200 XNORING_3 ( .A(A[3]), .B(B[3]), .Y(L[3]) );
  XNOR_GATE_199 XNORING_4 ( .A(A[4]), .B(B[4]), .Y(L[4]) );
  N_AND_N5_4 ANDING ( .A(L), .Y(Y) );
endmodule


module EQU_COMPARATOR_N5_3 ( A, B, Y );
  input [4:0] A;
  input [4:0] B;
  output Y;

  wire   [4:0] L;

  XNOR_GATE_198 XNORING_0 ( .A(A[0]), .B(B[0]), .Y(L[0]) );
  XNOR_GATE_197 XNORING_1 ( .A(A[1]), .B(B[1]), .Y(L[1]) );
  XNOR_GATE_196 XNORING_2 ( .A(A[2]), .B(B[2]), .Y(L[2]) );
  XNOR_GATE_195 XNORING_3 ( .A(A[3]), .B(B[3]), .Y(L[3]) );
  XNOR_GATE_194 XNORING_4 ( .A(A[4]), .B(B[4]), .Y(L[4]) );
  N_AND_N5_3 ANDING ( .A(L), .Y(Y) );
endmodule


module EQU_COMPARATOR_N5_2 ( A, B, Y );
  input [4:0] A;
  input [4:0] B;
  output Y;

  wire   [4:0] L;

  XNOR_GATE_193 XNORING_0 ( .A(A[0]), .B(B[0]), .Y(L[0]) );
  XNOR_GATE_192 XNORING_1 ( .A(A[1]), .B(B[1]), .Y(L[1]) );
  XNOR_GATE_191 XNORING_2 ( .A(A[2]), .B(B[2]), .Y(L[2]) );
  XNOR_GATE_190 XNORING_3 ( .A(A[3]), .B(B[3]), .Y(L[3]) );
  XNOR_GATE_189 XNORING_4 ( .A(A[4]), .B(B[4]), .Y(L[4]) );
  N_AND_N5_2 ANDING ( .A(L), .Y(Y) );
endmodule


module EQU_COMPARATOR_N5_1 ( A, B, Y );
  input [4:0] A;
  input [4:0] B;
  output Y;

  wire   [4:0] L;

  XNOR_GATE_188 XNORING_0 ( .A(A[0]), .B(B[0]), .Y(L[0]) );
  XNOR_GATE_187 XNORING_1 ( .A(A[1]), .B(B[1]), .Y(L[1]) );
  XNOR_GATE_186 XNORING_2 ( .A(A[2]), .B(B[2]), .Y(L[2]) );
  XNOR_GATE_185 XNORING_3 ( .A(A[3]), .B(B[3]), .Y(L[3]) );
  XNOR_GATE_184 XNORING_4 ( .A(A[4]), .B(B[4]), .Y(L[4]) );
  N_AND_N5_1 ANDING ( .A(L), .Y(Y) );
endmodule


module MUX51_GEN_N32_1 ( A, B, C, D, E, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [2:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n3, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157;

  NAND2_X1 U72 ( .A1(n157), .A2(n156), .ZN(Y[9]) );
  NAND2_X1 U73 ( .A1(n150), .A2(n149), .ZN(Y[8]) );
  NAND2_X1 U74 ( .A1(n148), .A2(n147), .ZN(Y[7]) );
  NAND2_X1 U75 ( .A1(n146), .A2(n145), .ZN(Y[6]) );
  NAND2_X1 U76 ( .A1(n144), .A2(n143), .ZN(Y[5]) );
  NAND2_X1 U77 ( .A1(n142), .A2(n141), .ZN(Y[4]) );
  NAND2_X1 U78 ( .A1(n140), .A2(n139), .ZN(Y[3]) );
  NAND2_X1 U79 ( .A1(n138), .A2(n137), .ZN(Y[31]) );
  NAND2_X1 U80 ( .A1(n136), .A2(n135), .ZN(Y[30]) );
  NAND2_X1 U81 ( .A1(n134), .A2(n133), .ZN(Y[2]) );
  NAND2_X1 U82 ( .A1(n132), .A2(n131), .ZN(Y[29]) );
  NAND2_X1 U83 ( .A1(n130), .A2(n129), .ZN(Y[28]) );
  NAND2_X1 U84 ( .A1(n128), .A2(n127), .ZN(Y[27]) );
  NAND2_X1 U85 ( .A1(n126), .A2(n125), .ZN(Y[26]) );
  NAND2_X1 U86 ( .A1(n124), .A2(n123), .ZN(Y[25]) );
  NAND2_X1 U87 ( .A1(n122), .A2(n121), .ZN(Y[24]) );
  NAND2_X1 U88 ( .A1(n120), .A2(n119), .ZN(Y[23]) );
  NAND2_X1 U89 ( .A1(n118), .A2(n117), .ZN(Y[22]) );
  NAND2_X1 U90 ( .A1(n116), .A2(n115), .ZN(Y[21]) );
  NAND2_X1 U91 ( .A1(n114), .A2(n113), .ZN(Y[20]) );
  NAND2_X1 U92 ( .A1(n112), .A2(n111), .ZN(Y[1]) );
  NAND2_X1 U93 ( .A1(n110), .A2(n109), .ZN(Y[19]) );
  NAND2_X1 U94 ( .A1(n108), .A2(n107), .ZN(Y[18]) );
  NAND2_X1 U95 ( .A1(n106), .A2(n105), .ZN(Y[17]) );
  NAND2_X1 U96 ( .A1(n104), .A2(n103), .ZN(Y[16]) );
  NAND2_X1 U97 ( .A1(n102), .A2(n101), .ZN(Y[15]) );
  NAND2_X1 U98 ( .A1(n100), .A2(n99), .ZN(Y[14]) );
  NAND2_X1 U99 ( .A1(n98), .A2(n97), .ZN(Y[13]) );
  NAND2_X1 U100 ( .A1(n96), .A2(n95), .ZN(Y[12]) );
  NAND2_X1 U101 ( .A1(n94), .A2(n93), .ZN(Y[11]) );
  NAND2_X1 U102 ( .A1(n92), .A2(n91), .ZN(Y[10]) );
  NAND2_X1 U103 ( .A1(n90), .A2(n89), .ZN(Y[0]) );
  BUF_X1 U1 ( .A(n155), .Z(n84) );
  BUF_X1 U2 ( .A(n155), .Z(n85) );
  BUF_X1 U3 ( .A(n155), .Z(n86) );
  NOR4_X1 U4 ( .A1(n78), .A2(n81), .A3(n75), .A4(n1), .ZN(n155) );
  AOI222_X1 U5 ( .A1(E[7]), .A2(n86), .B1(B[7]), .B2(n83), .C1(D[7]), .C2(n80), 
        .ZN(n147) );
  BUF_X1 U6 ( .A(n152), .Z(n77) );
  BUF_X1 U7 ( .A(n151), .Z(n3) );
  BUF_X1 U8 ( .A(n154), .Z(n83) );
  BUF_X1 U9 ( .A(n153), .Z(n80) );
  AOI22_X1 U10 ( .A1(C[7]), .A2(n77), .B1(A[7]), .B2(n3), .ZN(n148) );
  BUF_X1 U11 ( .A(n152), .Z(n75) );
  BUF_X1 U12 ( .A(n152), .Z(n76) );
  BUF_X1 U13 ( .A(n151), .Z(n1) );
  BUF_X1 U14 ( .A(n151), .Z(n2) );
  BUF_X1 U15 ( .A(n154), .Z(n81) );
  BUF_X1 U16 ( .A(n154), .Z(n82) );
  BUF_X1 U17 ( .A(n153), .Z(n78) );
  BUF_X1 U18 ( .A(n153), .Z(n79) );
  AOI222_X1 U19 ( .A1(E[0]), .A2(n84), .B1(B[0]), .B2(n81), .C1(D[0]), .C2(n78), .ZN(n89) );
  AOI222_X1 U20 ( .A1(E[1]), .A2(n84), .B1(B[1]), .B2(n81), .C1(D[1]), .C2(n78), .ZN(n111) );
  AOI222_X1 U21 ( .A1(E[2]), .A2(n85), .B1(B[2]), .B2(n82), .C1(D[2]), .C2(n79), .ZN(n133) );
  AOI222_X1 U22 ( .A1(E[3]), .A2(n85), .B1(B[3]), .B2(n83), .C1(D[3]), .C2(n80), .ZN(n139) );
  AOI222_X1 U23 ( .A1(E[4]), .A2(n86), .B1(B[4]), .B2(n83), .C1(D[4]), .C2(n80), .ZN(n141) );
  AOI222_X1 U24 ( .A1(E[5]), .A2(n86), .B1(B[5]), .B2(n83), .C1(D[5]), .C2(n80), .ZN(n143) );
  AOI222_X1 U25 ( .A1(E[6]), .A2(n86), .B1(B[6]), .B2(n83), .C1(D[6]), .C2(n80), .ZN(n145) );
  AOI222_X1 U26 ( .A1(E[8]), .A2(n86), .B1(B[8]), .B2(n83), .C1(D[8]), .C2(n80), .ZN(n149) );
  AOI222_X1 U27 ( .A1(E[9]), .A2(n86), .B1(B[9]), .B2(n83), .C1(D[9]), .C2(n80), .ZN(n156) );
  AOI222_X1 U28 ( .A1(E[10]), .A2(n84), .B1(B[10]), .B2(n81), .C1(D[10]), .C2(
        n78), .ZN(n91) );
  AOI222_X1 U29 ( .A1(E[11]), .A2(n84), .B1(B[11]), .B2(n81), .C1(D[11]), .C2(
        n78), .ZN(n93) );
  AOI222_X1 U30 ( .A1(E[12]), .A2(n84), .B1(B[12]), .B2(n81), .C1(D[12]), .C2(
        n78), .ZN(n95) );
  AOI222_X1 U31 ( .A1(E[13]), .A2(n84), .B1(B[13]), .B2(n81), .C1(D[13]), .C2(
        n78), .ZN(n97) );
  AOI222_X1 U32 ( .A1(E[14]), .A2(n84), .B1(B[14]), .B2(n81), .C1(D[14]), .C2(
        n78), .ZN(n99) );
  AOI222_X1 U33 ( .A1(E[15]), .A2(n84), .B1(B[15]), .B2(n81), .C1(D[15]), .C2(
        n78), .ZN(n101) );
  AOI222_X1 U34 ( .A1(E[16]), .A2(n84), .B1(B[16]), .B2(n81), .C1(D[16]), .C2(
        n78), .ZN(n103) );
  AOI222_X1 U35 ( .A1(E[17]), .A2(n84), .B1(B[17]), .B2(n81), .C1(D[17]), .C2(
        n78), .ZN(n105) );
  AOI222_X1 U36 ( .A1(E[18]), .A2(n84), .B1(B[18]), .B2(n81), .C1(D[18]), .C2(
        n78), .ZN(n107) );
  AOI222_X1 U37 ( .A1(E[19]), .A2(n84), .B1(B[19]), .B2(n81), .C1(D[19]), .C2(
        n78), .ZN(n109) );
  AOI222_X1 U38 ( .A1(E[20]), .A2(n84), .B1(B[20]), .B2(n82), .C1(D[20]), .C2(
        n79), .ZN(n113) );
  AOI222_X1 U39 ( .A1(E[21]), .A2(n85), .B1(B[21]), .B2(n82), .C1(D[21]), .C2(
        n79), .ZN(n115) );
  AOI222_X1 U40 ( .A1(E[22]), .A2(n85), .B1(B[22]), .B2(n82), .C1(D[22]), .C2(
        n79), .ZN(n117) );
  AOI222_X1 U41 ( .A1(E[23]), .A2(n85), .B1(B[23]), .B2(n82), .C1(D[23]), .C2(
        n79), .ZN(n119) );
  AOI222_X1 U42 ( .A1(E[24]), .A2(n85), .B1(B[24]), .B2(n82), .C1(D[24]), .C2(
        n79), .ZN(n121) );
  AOI222_X1 U43 ( .A1(E[25]), .A2(n85), .B1(B[25]), .B2(n82), .C1(D[25]), .C2(
        n79), .ZN(n123) );
  AOI222_X1 U44 ( .A1(E[26]), .A2(n85), .B1(B[26]), .B2(n82), .C1(D[26]), .C2(
        n79), .ZN(n125) );
  AOI222_X1 U45 ( .A1(E[27]), .A2(n85), .B1(B[27]), .B2(n82), .C1(D[27]), .C2(
        n79), .ZN(n127) );
  AOI222_X1 U46 ( .A1(E[28]), .A2(n85), .B1(B[28]), .B2(n82), .C1(D[28]), .C2(
        n79), .ZN(n129) );
  AOI222_X1 U47 ( .A1(E[29]), .A2(n85), .B1(B[29]), .B2(n82), .C1(D[29]), .C2(
        n79), .ZN(n131) );
  AOI222_X1 U48 ( .A1(E[30]), .A2(n85), .B1(B[30]), .B2(n82), .C1(D[30]), .C2(
        n79), .ZN(n135) );
  AOI222_X1 U49 ( .A1(E[31]), .A2(n85), .B1(B[31]), .B2(n82), .C1(D[31]), .C2(
        n79), .ZN(n137) );
  AND3_X1 U50 ( .A1(SEL[2]), .A2(n87), .A3(SEL[0]), .ZN(n152) );
  AND3_X1 U51 ( .A1(SEL[2]), .A2(SEL[1]), .A3(SEL[0]), .ZN(n151) );
  AND3_X1 U52 ( .A1(SEL[1]), .A2(n88), .A3(SEL[2]), .ZN(n154) );
  AND3_X1 U53 ( .A1(n88), .A2(n87), .A3(SEL[2]), .ZN(n153) );
  AOI22_X1 U54 ( .A1(C[3]), .A2(n77), .B1(A[3]), .B2(n3), .ZN(n140) );
  AOI22_X1 U55 ( .A1(C[4]), .A2(n77), .B1(A[4]), .B2(n3), .ZN(n142) );
  AOI22_X1 U56 ( .A1(C[5]), .A2(n77), .B1(A[5]), .B2(n3), .ZN(n144) );
  AOI22_X1 U57 ( .A1(C[6]), .A2(n77), .B1(A[6]), .B2(n3), .ZN(n146) );
  AOI22_X1 U58 ( .A1(C[8]), .A2(n77), .B1(A[8]), .B2(n3), .ZN(n150) );
  AOI22_X1 U59 ( .A1(C[31]), .A2(n77), .B1(A[31]), .B2(n3), .ZN(n138) );
  AOI22_X1 U60 ( .A1(C[0]), .A2(n76), .B1(A[0]), .B2(n2), .ZN(n90) );
  AOI22_X1 U61 ( .A1(C[1]), .A2(n75), .B1(A[1]), .B2(n1), .ZN(n112) );
  AOI22_X1 U62 ( .A1(C[2]), .A2(n76), .B1(A[2]), .B2(n2), .ZN(n134) );
  AOI22_X1 U63 ( .A1(C[9]), .A2(n75), .B1(A[9]), .B2(n1), .ZN(n157) );
  AOI22_X1 U64 ( .A1(C[10]), .A2(n75), .B1(A[10]), .B2(n1), .ZN(n92) );
  AOI22_X1 U65 ( .A1(C[11]), .A2(n75), .B1(A[11]), .B2(n1), .ZN(n94) );
  AOI22_X1 U66 ( .A1(C[12]), .A2(n75), .B1(A[12]), .B2(n1), .ZN(n96) );
  AOI22_X1 U67 ( .A1(C[13]), .A2(n75), .B1(A[13]), .B2(n1), .ZN(n98) );
  AOI22_X1 U68 ( .A1(C[14]), .A2(n75), .B1(A[14]), .B2(n1), .ZN(n100) );
  AOI22_X1 U69 ( .A1(C[15]), .A2(n75), .B1(A[15]), .B2(n1), .ZN(n102) );
  AOI22_X1 U70 ( .A1(C[16]), .A2(n75), .B1(A[16]), .B2(n1), .ZN(n104) );
  AOI22_X1 U71 ( .A1(C[17]), .A2(n75), .B1(A[17]), .B2(n1), .ZN(n106) );
  AOI22_X1 U104 ( .A1(C[18]), .A2(n75), .B1(A[18]), .B2(n1), .ZN(n108) );
  AOI22_X1 U105 ( .A1(C[19]), .A2(n75), .B1(A[19]), .B2(n1), .ZN(n110) );
  AOI22_X1 U106 ( .A1(C[20]), .A2(n76), .B1(A[20]), .B2(n2), .ZN(n114) );
  AOI22_X1 U107 ( .A1(C[21]), .A2(n76), .B1(A[21]), .B2(n2), .ZN(n116) );
  AOI22_X1 U108 ( .A1(C[22]), .A2(n76), .B1(A[22]), .B2(n2), .ZN(n118) );
  AOI22_X1 U109 ( .A1(C[23]), .A2(n76), .B1(A[23]), .B2(n2), .ZN(n120) );
  AOI22_X1 U110 ( .A1(C[24]), .A2(n76), .B1(A[24]), .B2(n2), .ZN(n122) );
  AOI22_X1 U111 ( .A1(C[25]), .A2(n76), .B1(A[25]), .B2(n2), .ZN(n124) );
  AOI22_X1 U112 ( .A1(C[26]), .A2(n76), .B1(A[26]), .B2(n2), .ZN(n126) );
  AOI22_X1 U113 ( .A1(C[27]), .A2(n76), .B1(A[27]), .B2(n2), .ZN(n128) );
  AOI22_X1 U114 ( .A1(C[28]), .A2(n76), .B1(A[28]), .B2(n2), .ZN(n130) );
  AOI22_X1 U115 ( .A1(C[29]), .A2(n76), .B1(A[29]), .B2(n2), .ZN(n132) );
  AOI22_X1 U116 ( .A1(C[30]), .A2(n76), .B1(A[30]), .B2(n2), .ZN(n136) );
  INV_X1 U117 ( .A(SEL[1]), .ZN(n87) );
  INV_X1 U118 ( .A(SEL[0]), .ZN(n88) );
endmodule


module MUX41_GEN_N32_3 ( A, B, C, D, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] SEL;
  output [31:0] Y;
  wire   n250, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249;

  OAI221_X4 U1 ( .B1(n19), .B2(n42), .C1(n16), .C2(n41), .A(n40), .ZN(Y[2]) );
  OAI221_X4 U2 ( .B1(n19), .B2(n49), .C1(n16), .C2(n48), .A(n47), .ZN(Y[3]) );
  OAI221_X4 U3 ( .B1(n19), .B2(n56), .C1(n16), .C2(n55), .A(n54), .ZN(Y[4]) );
  OAI221_X4 U4 ( .B1(n19), .B2(n63), .C1(n16), .C2(n62), .A(n61), .ZN(Y[5]) );
  NOR2_X1 U5 ( .A1(n16), .A2(n27), .ZN(n4) );
  NOR2_X2 U6 ( .A1(n16), .A2(n34), .ZN(n6) );
  OAI221_X2 U7 ( .B1(n18), .B2(n70), .C1(n15), .C2(n69), .A(n68), .ZN(Y[6]) );
  OAI221_X2 U8 ( .B1(n18), .B2(n77), .C1(n15), .C2(n76), .A(n75), .ZN(Y[7]) );
  OAI221_X2 U9 ( .B1(n18), .B2(n84), .C1(n15), .C2(n83), .A(n82), .ZN(Y[8]) );
  OAI221_X2 U10 ( .B1(n18), .B2(n91), .C1(n15), .C2(n90), .A(n89), .ZN(Y[9])
         );
  OAI221_X2 U11 ( .B1(n18), .B2(n98), .C1(n15), .C2(n97), .A(n96), .ZN(Y[10])
         );
  OAI221_X2 U12 ( .B1(n18), .B2(n105), .C1(n15), .C2(n104), .A(n103), .ZN(
        Y[11]) );
  OR2_X1 U13 ( .A1(n26), .A2(n25), .ZN(n1) );
  BUF_X2 U14 ( .A(n247), .Z(n16) );
  BUF_X4 U15 ( .A(n249), .Z(n19) );
  BUF_X4 U16 ( .A(n240), .Z(n10) );
  OR3_X4 U17 ( .A1(n3), .A2(n4), .A3(n1), .ZN(Y[0]) );
  OR2_X1 U18 ( .A1(n5), .A2(n7), .ZN(n2) );
  OR2_X4 U19 ( .A1(n2), .A2(n6), .ZN(Y[1]) );
  OAI221_X2 U20 ( .B1(n18), .B2(n112), .C1(n15), .C2(n111), .A(n110), .ZN(
        Y[12]) );
  OAI221_X2 U21 ( .B1(n18), .B2(n119), .C1(n15), .C2(n118), .A(n117), .ZN(
        Y[13]) );
  OAI221_X2 U22 ( .B1(n18), .B2(n126), .C1(n15), .C2(n125), .A(n124), .ZN(
        Y[14]) );
  CLKBUF_X1 U23 ( .A(n247), .Z(n15) );
  NOR2_X1 U24 ( .A1(n19), .A2(n28), .ZN(n3) );
  NOR2_X1 U25 ( .A1(n19), .A2(n35), .ZN(n5) );
  INV_X1 U26 ( .A(n33), .ZN(n7) );
  CLKBUF_X1 U27 ( .A(n247), .Z(n14) );
  CLKBUF_X1 U28 ( .A(n249), .Z(n17) );
  BUF_X2 U29 ( .A(n242), .Z(n13) );
  NAND3_X1 U30 ( .A1(n19), .A2(n13), .A3(n10), .ZN(n247) );
  BUF_X1 U31 ( .A(n240), .Z(n9) );
  BUF_X1 U32 ( .A(n240), .Z(n8) );
  BUF_X1 U33 ( .A(n242), .Z(n11) );
  BUF_X1 U34 ( .A(n249), .Z(n18) );
  NOR2_X1 U35 ( .A1(n116), .A2(n115), .ZN(n117) );
  NOR2_X1 U36 ( .A1(n109), .A2(n108), .ZN(n110) );
  NOR2_X1 U37 ( .A1(n123), .A2(n122), .ZN(n124) );
  NOR2_X1 U38 ( .A1(n67), .A2(n66), .ZN(n68) );
  NOR2_X1 U39 ( .A1(n74), .A2(n73), .ZN(n75) );
  NOR2_X1 U40 ( .A1(n81), .A2(n80), .ZN(n82) );
  NOR2_X1 U41 ( .A1(n88), .A2(n87), .ZN(n89) );
  NOR2_X1 U42 ( .A1(n95), .A2(n94), .ZN(n96) );
  NOR2_X1 U43 ( .A1(n102), .A2(n101), .ZN(n103) );
  NOR2_X1 U44 ( .A1(n60), .A2(n59), .ZN(n61) );
  NOR2_X1 U45 ( .A1(n53), .A2(n52), .ZN(n54) );
  NOR2_X1 U46 ( .A1(n39), .A2(n38), .ZN(n40) );
  NOR2_X1 U47 ( .A1(n32), .A2(n31), .ZN(n33) );
  NOR2_X1 U48 ( .A1(n46), .A2(n45), .ZN(n47) );
  NOR2_X1 U49 ( .A1(n244), .A2(n243), .ZN(n245) );
  NOR2_X1 U50 ( .A1(n235), .A2(n234), .ZN(n236) );
  NOR2_X1 U51 ( .A1(n214), .A2(n213), .ZN(n215) );
  NOR2_X1 U52 ( .A1(n200), .A2(n199), .ZN(n201) );
  NOR2_X1 U53 ( .A1(n221), .A2(n220), .ZN(n222) );
  NOR2_X1 U54 ( .A1(n207), .A2(n206), .ZN(n208) );
  NOR2_X1 U55 ( .A1(n228), .A2(n227), .ZN(n229) );
  NOR2_X1 U56 ( .A1(n193), .A2(n192), .ZN(n194) );
  NOR2_X1 U57 ( .A1(n144), .A2(n143), .ZN(n145) );
  NOR2_X1 U58 ( .A1(n151), .A2(n150), .ZN(n152) );
  NOR2_X1 U59 ( .A1(n158), .A2(n157), .ZN(n159) );
  NOR2_X1 U60 ( .A1(n165), .A2(n164), .ZN(n166) );
  NOR2_X1 U61 ( .A1(n172), .A2(n171), .ZN(n173) );
  NOR2_X1 U62 ( .A1(n179), .A2(n178), .ZN(n180) );
  NOR2_X1 U63 ( .A1(n186), .A2(n185), .ZN(n187) );
  NOR2_X1 U64 ( .A1(n12), .A2(n114), .ZN(n115) );
  NOR2_X1 U65 ( .A1(n12), .A2(n107), .ZN(n108) );
  NOR2_X1 U66 ( .A1(n12), .A2(n121), .ZN(n122) );
  NOR2_X1 U67 ( .A1(n12), .A2(n142), .ZN(n143) );
  NOR2_X1 U68 ( .A1(n12), .A2(n149), .ZN(n150) );
  NOR2_X1 U69 ( .A1(n12), .A2(n135), .ZN(n136) );
  NOR2_X1 U70 ( .A1(n12), .A2(n65), .ZN(n66) );
  NOR2_X1 U71 ( .A1(n12), .A2(n72), .ZN(n73) );
  NOR2_X1 U72 ( .A1(n12), .A2(n79), .ZN(n80) );
  NOR2_X1 U73 ( .A1(n12), .A2(n86), .ZN(n87) );
  NOR2_X1 U74 ( .A1(n12), .A2(n93), .ZN(n94) );
  NOR2_X1 U75 ( .A1(n12), .A2(n100), .ZN(n101) );
  NOR2_X1 U76 ( .A1(n13), .A2(n44), .ZN(n45) );
  NOR2_X1 U77 ( .A1(n13), .A2(n24), .ZN(n25) );
  NOR2_X1 U78 ( .A1(n13), .A2(n37), .ZN(n38) );
  NOR2_X1 U79 ( .A1(n13), .A2(n30), .ZN(n31) );
  NOR2_X1 U80 ( .A1(n13), .A2(n51), .ZN(n52) );
  NOR2_X1 U81 ( .A1(n13), .A2(n58), .ZN(n59) );
  NOR2_X1 U82 ( .A1(n11), .A2(n156), .ZN(n157) );
  NOR2_X1 U83 ( .A1(n11), .A2(n163), .ZN(n164) );
  NOR2_X1 U84 ( .A1(n11), .A2(n170), .ZN(n171) );
  NOR2_X1 U85 ( .A1(n11), .A2(n177), .ZN(n178) );
  NOR2_X1 U86 ( .A1(n11), .A2(n184), .ZN(n185) );
  NOR2_X1 U87 ( .A1(n11), .A2(n233), .ZN(n234) );
  NOR2_X1 U88 ( .A1(n11), .A2(n241), .ZN(n243) );
  NOR2_X1 U89 ( .A1(n11), .A2(n191), .ZN(n192) );
  NOR2_X1 U90 ( .A1(n11), .A2(n212), .ZN(n213) );
  NOR2_X1 U91 ( .A1(n11), .A2(n198), .ZN(n199) );
  NOR2_X1 U92 ( .A1(n11), .A2(n219), .ZN(n220) );
  NOR2_X1 U93 ( .A1(n11), .A2(n205), .ZN(n206) );
  NOR2_X1 U94 ( .A1(n11), .A2(n226), .ZN(n227) );
  NOR2_X1 U95 ( .A1(n10), .A2(n43), .ZN(n46) );
  NOR2_X1 U96 ( .A1(n10), .A2(n23), .ZN(n26) );
  NOR2_X1 U97 ( .A1(n10), .A2(n36), .ZN(n39) );
  NOR2_X1 U98 ( .A1(n10), .A2(n29), .ZN(n32) );
  NOR2_X1 U99 ( .A1(n10), .A2(n50), .ZN(n53) );
  NOR2_X1 U100 ( .A1(n10), .A2(n57), .ZN(n60) );
  NOR2_X1 U101 ( .A1(n9), .A2(n113), .ZN(n116) );
  NOR2_X1 U102 ( .A1(n9), .A2(n106), .ZN(n109) );
  NOR2_X1 U103 ( .A1(n9), .A2(n120), .ZN(n123) );
  NOR2_X1 U104 ( .A1(n9), .A2(n141), .ZN(n144) );
  NOR2_X1 U105 ( .A1(n9), .A2(n148), .ZN(n151) );
  NOR2_X1 U106 ( .A1(n8), .A2(n155), .ZN(n158) );
  NOR2_X1 U107 ( .A1(n8), .A2(n162), .ZN(n165) );
  NOR2_X1 U108 ( .A1(n8), .A2(n169), .ZN(n172) );
  NOR2_X1 U109 ( .A1(n8), .A2(n176), .ZN(n179) );
  NOR2_X1 U110 ( .A1(n8), .A2(n183), .ZN(n186) );
  NOR2_X1 U111 ( .A1(n8), .A2(n232), .ZN(n235) );
  NOR2_X1 U112 ( .A1(n8), .A2(n239), .ZN(n244) );
  NOR2_X1 U113 ( .A1(n8), .A2(n190), .ZN(n193) );
  NOR2_X1 U114 ( .A1(n9), .A2(n134), .ZN(n137) );
  NOR2_X1 U115 ( .A1(n8), .A2(n211), .ZN(n214) );
  NOR2_X1 U116 ( .A1(n8), .A2(n197), .ZN(n200) );
  NOR2_X1 U117 ( .A1(n8), .A2(n218), .ZN(n221) );
  NOR2_X1 U118 ( .A1(n8), .A2(n204), .ZN(n207) );
  NOR2_X1 U119 ( .A1(n8), .A2(n225), .ZN(n228) );
  NOR2_X1 U120 ( .A1(n9), .A2(n64), .ZN(n67) );
  NOR2_X1 U121 ( .A1(n9), .A2(n71), .ZN(n74) );
  NOR2_X1 U122 ( .A1(n9), .A2(n78), .ZN(n81) );
  NOR2_X1 U123 ( .A1(n9), .A2(n85), .ZN(n88) );
  NOR2_X1 U124 ( .A1(n9), .A2(n92), .ZN(n95) );
  NOR2_X1 U125 ( .A1(n9), .A2(n99), .ZN(n102) );
  NOR2_X1 U126 ( .A1(n130), .A2(n129), .ZN(n131) );
  NOR2_X1 U127 ( .A1(n9), .A2(n127), .ZN(n130) );
  NOR2_X1 U128 ( .A1(n12), .A2(n128), .ZN(n129) );
  NOR2_X1 U129 ( .A1(n137), .A2(n136), .ZN(n138) );
  BUF_X1 U130 ( .A(n242), .Z(n12) );
  CLKBUF_X1 U131 ( .A(n250), .Z(Y[15]) );
  INV_X1 U132 ( .A(SEL[0]), .ZN(n21) );
  NAND2_X1 U133 ( .A1(SEL[1]), .A2(n21), .ZN(n249) );
  INV_X1 U134 ( .A(B[0]), .ZN(n28) );
  NAND2_X1 U135 ( .A1(SEL[1]), .A2(SEL[0]), .ZN(n242) );
  INV_X1 U136 ( .A(SEL[1]), .ZN(n22) );
  NAND2_X1 U137 ( .A1(n22), .A2(SEL[0]), .ZN(n240) );
  INV_X1 U138 ( .A(D[0]), .ZN(n27) );
  INV_X1 U139 ( .A(C[0]), .ZN(n23) );
  INV_X1 U140 ( .A(A[0]), .ZN(n24) );
  INV_X1 U141 ( .A(B[1]), .ZN(n35) );
  INV_X1 U142 ( .A(D[1]), .ZN(n34) );
  INV_X1 U143 ( .A(C[1]), .ZN(n29) );
  INV_X1 U144 ( .A(A[1]), .ZN(n30) );
  INV_X1 U145 ( .A(B[2]), .ZN(n42) );
  INV_X1 U146 ( .A(D[2]), .ZN(n41) );
  INV_X1 U147 ( .A(C[2]), .ZN(n36) );
  INV_X1 U148 ( .A(A[2]), .ZN(n37) );
  INV_X1 U149 ( .A(B[3]), .ZN(n49) );
  INV_X1 U150 ( .A(D[3]), .ZN(n48) );
  INV_X1 U151 ( .A(C[3]), .ZN(n43) );
  INV_X1 U152 ( .A(A[3]), .ZN(n44) );
  INV_X1 U153 ( .A(B[4]), .ZN(n56) );
  INV_X1 U154 ( .A(D[4]), .ZN(n55) );
  INV_X1 U155 ( .A(C[4]), .ZN(n50) );
  INV_X1 U156 ( .A(A[4]), .ZN(n51) );
  INV_X1 U157 ( .A(B[5]), .ZN(n63) );
  INV_X1 U158 ( .A(D[5]), .ZN(n62) );
  INV_X1 U159 ( .A(C[5]), .ZN(n57) );
  INV_X1 U160 ( .A(A[5]), .ZN(n58) );
  INV_X1 U161 ( .A(B[6]), .ZN(n70) );
  INV_X1 U162 ( .A(D[6]), .ZN(n69) );
  INV_X1 U163 ( .A(C[6]), .ZN(n64) );
  INV_X1 U164 ( .A(A[6]), .ZN(n65) );
  INV_X1 U165 ( .A(B[7]), .ZN(n77) );
  INV_X1 U166 ( .A(D[7]), .ZN(n76) );
  INV_X1 U167 ( .A(C[7]), .ZN(n71) );
  INV_X1 U168 ( .A(A[7]), .ZN(n72) );
  INV_X1 U169 ( .A(B[8]), .ZN(n84) );
  INV_X1 U170 ( .A(D[8]), .ZN(n83) );
  INV_X1 U171 ( .A(C[8]), .ZN(n78) );
  INV_X1 U172 ( .A(A[8]), .ZN(n79) );
  INV_X1 U173 ( .A(B[9]), .ZN(n91) );
  INV_X1 U174 ( .A(D[9]), .ZN(n90) );
  INV_X1 U175 ( .A(C[9]), .ZN(n85) );
  INV_X1 U176 ( .A(A[9]), .ZN(n86) );
  INV_X1 U177 ( .A(B[10]), .ZN(n98) );
  INV_X1 U178 ( .A(D[10]), .ZN(n97) );
  INV_X1 U179 ( .A(C[10]), .ZN(n92) );
  INV_X1 U180 ( .A(A[10]), .ZN(n93) );
  INV_X1 U181 ( .A(B[11]), .ZN(n105) );
  INV_X1 U182 ( .A(D[11]), .ZN(n104) );
  INV_X1 U183 ( .A(C[11]), .ZN(n99) );
  INV_X1 U184 ( .A(A[11]), .ZN(n100) );
  INV_X1 U185 ( .A(B[12]), .ZN(n112) );
  INV_X1 U186 ( .A(D[12]), .ZN(n111) );
  INV_X1 U187 ( .A(C[12]), .ZN(n106) );
  INV_X1 U188 ( .A(A[12]), .ZN(n107) );
  INV_X1 U189 ( .A(B[13]), .ZN(n119) );
  INV_X1 U190 ( .A(D[13]), .ZN(n118) );
  INV_X1 U191 ( .A(C[13]), .ZN(n113) );
  INV_X1 U192 ( .A(A[13]), .ZN(n114) );
  INV_X1 U193 ( .A(B[14]), .ZN(n126) );
  INV_X1 U194 ( .A(D[14]), .ZN(n125) );
  INV_X1 U195 ( .A(C[14]), .ZN(n120) );
  INV_X1 U196 ( .A(A[14]), .ZN(n121) );
  INV_X1 U197 ( .A(B[15]), .ZN(n133) );
  INV_X1 U198 ( .A(D[15]), .ZN(n132) );
  INV_X1 U199 ( .A(C[15]), .ZN(n127) );
  INV_X1 U200 ( .A(A[15]), .ZN(n128) );
  OAI221_X1 U201 ( .B1(n18), .B2(n133), .C1(n15), .C2(n132), .A(n131), .ZN(
        n250) );
  INV_X1 U202 ( .A(B[16]), .ZN(n140) );
  INV_X1 U203 ( .A(D[16]), .ZN(n139) );
  INV_X1 U204 ( .A(C[16]), .ZN(n134) );
  INV_X1 U205 ( .A(A[16]), .ZN(n135) );
  OAI221_X1 U206 ( .B1(n18), .B2(n140), .C1(n15), .C2(n139), .A(n138), .ZN(
        Y[16]) );
  INV_X1 U207 ( .A(B[17]), .ZN(n147) );
  INV_X1 U208 ( .A(D[17]), .ZN(n146) );
  INV_X1 U209 ( .A(C[17]), .ZN(n141) );
  INV_X1 U210 ( .A(A[17]), .ZN(n142) );
  OAI221_X1 U211 ( .B1(n18), .B2(n147), .C1(n15), .C2(n146), .A(n145), .ZN(
        Y[17]) );
  INV_X1 U212 ( .A(B[18]), .ZN(n154) );
  INV_X1 U213 ( .A(D[18]), .ZN(n153) );
  INV_X1 U214 ( .A(C[18]), .ZN(n148) );
  INV_X1 U215 ( .A(A[18]), .ZN(n149) );
  OAI221_X1 U216 ( .B1(n18), .B2(n154), .C1(n15), .C2(n153), .A(n152), .ZN(
        Y[18]) );
  INV_X1 U217 ( .A(B[19]), .ZN(n161) );
  INV_X1 U218 ( .A(D[19]), .ZN(n160) );
  INV_X1 U219 ( .A(C[19]), .ZN(n155) );
  INV_X1 U220 ( .A(A[19]), .ZN(n156) );
  OAI221_X1 U221 ( .B1(n17), .B2(n161), .C1(n14), .C2(n160), .A(n159), .ZN(
        Y[19]) );
  INV_X1 U222 ( .A(B[20]), .ZN(n168) );
  INV_X1 U223 ( .A(D[20]), .ZN(n167) );
  INV_X1 U224 ( .A(C[20]), .ZN(n162) );
  INV_X1 U225 ( .A(A[20]), .ZN(n163) );
  OAI221_X1 U226 ( .B1(n17), .B2(n168), .C1(n14), .C2(n167), .A(n166), .ZN(
        Y[20]) );
  INV_X1 U227 ( .A(B[21]), .ZN(n175) );
  INV_X1 U228 ( .A(D[21]), .ZN(n174) );
  INV_X1 U229 ( .A(C[21]), .ZN(n169) );
  INV_X1 U230 ( .A(A[21]), .ZN(n170) );
  OAI221_X1 U231 ( .B1(n17), .B2(n175), .C1(n14), .C2(n174), .A(n173), .ZN(
        Y[21]) );
  INV_X1 U232 ( .A(B[22]), .ZN(n182) );
  INV_X1 U233 ( .A(D[22]), .ZN(n181) );
  INV_X1 U234 ( .A(C[22]), .ZN(n176) );
  INV_X1 U235 ( .A(A[22]), .ZN(n177) );
  OAI221_X1 U236 ( .B1(n17), .B2(n182), .C1(n14), .C2(n181), .A(n180), .ZN(
        Y[22]) );
  INV_X1 U237 ( .A(B[23]), .ZN(n189) );
  INV_X1 U238 ( .A(D[23]), .ZN(n188) );
  INV_X1 U239 ( .A(C[23]), .ZN(n183) );
  INV_X1 U240 ( .A(A[23]), .ZN(n184) );
  OAI221_X1 U241 ( .B1(n17), .B2(n189), .C1(n14), .C2(n188), .A(n187), .ZN(
        Y[23]) );
  INV_X1 U242 ( .A(B[24]), .ZN(n196) );
  INV_X1 U243 ( .A(D[24]), .ZN(n195) );
  INV_X1 U244 ( .A(C[24]), .ZN(n190) );
  INV_X1 U245 ( .A(A[24]), .ZN(n191) );
  OAI221_X1 U246 ( .B1(n17), .B2(n196), .C1(n14), .C2(n195), .A(n194), .ZN(
        Y[24]) );
  INV_X1 U247 ( .A(B[25]), .ZN(n203) );
  INV_X1 U248 ( .A(D[25]), .ZN(n202) );
  INV_X1 U249 ( .A(C[25]), .ZN(n197) );
  INV_X1 U250 ( .A(A[25]), .ZN(n198) );
  OAI221_X1 U251 ( .B1(n17), .B2(n203), .C1(n14), .C2(n202), .A(n201), .ZN(
        Y[25]) );
  INV_X1 U252 ( .A(B[26]), .ZN(n210) );
  INV_X1 U253 ( .A(D[26]), .ZN(n209) );
  INV_X1 U254 ( .A(C[26]), .ZN(n204) );
  INV_X1 U255 ( .A(A[26]), .ZN(n205) );
  OAI221_X1 U256 ( .B1(n17), .B2(n210), .C1(n14), .C2(n209), .A(n208), .ZN(
        Y[26]) );
  INV_X1 U257 ( .A(B[27]), .ZN(n217) );
  INV_X1 U258 ( .A(D[27]), .ZN(n216) );
  INV_X1 U259 ( .A(C[27]), .ZN(n211) );
  INV_X1 U260 ( .A(A[27]), .ZN(n212) );
  OAI221_X1 U261 ( .B1(n17), .B2(n217), .C1(n14), .C2(n216), .A(n215), .ZN(
        Y[27]) );
  INV_X1 U262 ( .A(B[28]), .ZN(n224) );
  INV_X1 U263 ( .A(D[28]), .ZN(n223) );
  INV_X1 U264 ( .A(C[28]), .ZN(n218) );
  INV_X1 U265 ( .A(A[28]), .ZN(n219) );
  OAI221_X1 U266 ( .B1(n17), .B2(n224), .C1(n14), .C2(n223), .A(n222), .ZN(
        Y[28]) );
  INV_X1 U267 ( .A(B[29]), .ZN(n231) );
  INV_X1 U268 ( .A(D[29]), .ZN(n230) );
  INV_X1 U269 ( .A(C[29]), .ZN(n225) );
  INV_X1 U270 ( .A(A[29]), .ZN(n226) );
  OAI221_X1 U271 ( .B1(n17), .B2(n231), .C1(n14), .C2(n230), .A(n229), .ZN(
        Y[29]) );
  INV_X1 U272 ( .A(B[30]), .ZN(n238) );
  INV_X1 U273 ( .A(D[30]), .ZN(n237) );
  INV_X1 U274 ( .A(C[30]), .ZN(n232) );
  INV_X1 U275 ( .A(A[30]), .ZN(n233) );
  OAI221_X1 U276 ( .B1(n17), .B2(n238), .C1(n14), .C2(n237), .A(n236), .ZN(
        Y[30]) );
  INV_X1 U277 ( .A(B[31]), .ZN(n248) );
  INV_X1 U278 ( .A(D[31]), .ZN(n246) );
  INV_X1 U279 ( .A(C[31]), .ZN(n239) );
  INV_X1 U280 ( .A(A[31]), .ZN(n241) );
  OAI221_X1 U281 ( .B1(n17), .B2(n248), .C1(n14), .C2(n246), .A(n245), .ZN(
        Y[31]) );
endmodule


module MUX41_GEN_N32_2 ( A, B, C, D, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150;

  NAND2_X1 U70 ( .A1(n150), .A2(n149), .ZN(Y[9]) );
  NAND2_X1 U71 ( .A1(n144), .A2(n143), .ZN(Y[8]) );
  NAND2_X1 U72 ( .A1(n142), .A2(n141), .ZN(Y[7]) );
  NAND2_X1 U73 ( .A1(n140), .A2(n139), .ZN(Y[6]) );
  NAND2_X1 U74 ( .A1(n138), .A2(n137), .ZN(Y[5]) );
  NAND2_X1 U75 ( .A1(n136), .A2(n135), .ZN(Y[4]) );
  NAND2_X1 U76 ( .A1(n134), .A2(n133), .ZN(Y[3]) );
  NAND2_X1 U77 ( .A1(n132), .A2(n131), .ZN(Y[31]) );
  NAND2_X1 U78 ( .A1(n130), .A2(n129), .ZN(Y[30]) );
  NAND2_X1 U79 ( .A1(n128), .A2(n127), .ZN(Y[2]) );
  NAND2_X1 U80 ( .A1(n126), .A2(n125), .ZN(Y[29]) );
  NAND2_X1 U81 ( .A1(n124), .A2(n123), .ZN(Y[28]) );
  NAND2_X1 U82 ( .A1(n122), .A2(n121), .ZN(Y[27]) );
  NAND2_X1 U83 ( .A1(n120), .A2(n119), .ZN(Y[26]) );
  NAND2_X1 U84 ( .A1(n118), .A2(n117), .ZN(Y[25]) );
  NAND2_X1 U85 ( .A1(n116), .A2(n115), .ZN(Y[24]) );
  NAND2_X1 U86 ( .A1(n114), .A2(n113), .ZN(Y[23]) );
  NAND2_X1 U87 ( .A1(n112), .A2(n111), .ZN(Y[22]) );
  NAND2_X1 U88 ( .A1(n110), .A2(n109), .ZN(Y[21]) );
  NAND2_X1 U89 ( .A1(n108), .A2(n107), .ZN(Y[20]) );
  NAND2_X1 U90 ( .A1(n106), .A2(n105), .ZN(Y[1]) );
  NAND2_X1 U91 ( .A1(n104), .A2(n103), .ZN(Y[19]) );
  NAND2_X1 U92 ( .A1(n102), .A2(n101), .ZN(Y[18]) );
  NAND2_X1 U93 ( .A1(n100), .A2(n99), .ZN(Y[17]) );
  NAND2_X1 U94 ( .A1(n98), .A2(n97), .ZN(Y[16]) );
  NAND2_X1 U95 ( .A1(n96), .A2(n95), .ZN(Y[15]) );
  NAND2_X1 U96 ( .A1(n94), .A2(n93), .ZN(Y[14]) );
  NAND2_X1 U97 ( .A1(n92), .A2(n91), .ZN(Y[13]) );
  NAND2_X1 U98 ( .A1(n90), .A2(n89), .ZN(Y[12]) );
  NAND2_X1 U99 ( .A1(n88), .A2(n87), .ZN(Y[11]) );
  NAND2_X1 U100 ( .A1(n86), .A2(n85), .ZN(Y[10]) );
  NAND2_X1 U101 ( .A1(n84), .A2(n83), .ZN(Y[0]) );
  BUF_X1 U1 ( .A(n146), .Z(n73) );
  BUF_X1 U2 ( .A(n146), .Z(n74) );
  BUF_X1 U3 ( .A(n146), .Z(n75) );
  NOR3_X1 U4 ( .A1(n78), .A2(n72), .A3(n81), .ZN(n146) );
  BUF_X1 U5 ( .A(n147), .Z(n78) );
  BUF_X1 U6 ( .A(n148), .Z(n81) );
  BUF_X1 U7 ( .A(n145), .Z(n72) );
  BUF_X1 U8 ( .A(n147), .Z(n77) );
  BUF_X1 U9 ( .A(n147), .Z(n76) );
  BUF_X1 U10 ( .A(n148), .Z(n80) );
  BUF_X1 U11 ( .A(n148), .Z(n79) );
  BUF_X1 U12 ( .A(n145), .Z(n2) );
  BUF_X1 U13 ( .A(n145), .Z(n1) );
  NOR2_X1 U14 ( .A1(n82), .A2(SEL[1]), .ZN(n147) );
  AND2_X1 U15 ( .A1(SEL[1]), .A2(n82), .ZN(n148) );
  AND2_X1 U16 ( .A1(SEL[0]), .A2(SEL[1]), .ZN(n145) );
  INV_X1 U17 ( .A(SEL[0]), .ZN(n82) );
  AOI22_X1 U18 ( .A1(D[0]), .A2(n73), .B1(A[0]), .B2(n72), .ZN(n84) );
  AOI22_X1 U19 ( .A1(B[0]), .A2(n81), .B1(C[0]), .B2(n78), .ZN(n83) );
  AOI22_X1 U20 ( .A1(D[1]), .A2(n73), .B1(A[1]), .B2(n2), .ZN(n106) );
  AOI22_X1 U21 ( .A1(B[1]), .A2(n80), .B1(C[1]), .B2(n77), .ZN(n105) );
  AOI22_X1 U22 ( .A1(D[2]), .A2(n74), .B1(A[2]), .B2(n1), .ZN(n128) );
  AOI22_X1 U23 ( .A1(B[2]), .A2(n79), .B1(C[2]), .B2(n76), .ZN(n127) );
  AOI22_X1 U24 ( .A1(D[3]), .A2(n74), .B1(A[3]), .B2(n1), .ZN(n134) );
  AOI22_X1 U25 ( .A1(B[3]), .A2(n79), .B1(C[3]), .B2(n76), .ZN(n133) );
  AOI22_X1 U26 ( .A1(D[4]), .A2(n75), .B1(A[4]), .B2(n1), .ZN(n136) );
  AOI22_X1 U27 ( .A1(B[4]), .A2(n79), .B1(C[4]), .B2(n76), .ZN(n135) );
  AOI22_X1 U28 ( .A1(D[5]), .A2(n75), .B1(A[5]), .B2(n1), .ZN(n138) );
  AOI22_X1 U29 ( .A1(B[5]), .A2(n79), .B1(C[5]), .B2(n76), .ZN(n137) );
  AOI22_X1 U30 ( .A1(D[6]), .A2(n75), .B1(A[6]), .B2(n1), .ZN(n140) );
  AOI22_X1 U31 ( .A1(B[6]), .A2(n79), .B1(C[6]), .B2(n76), .ZN(n139) );
  AOI22_X1 U32 ( .A1(D[7]), .A2(n75), .B1(A[7]), .B2(n1), .ZN(n142) );
  AOI22_X1 U33 ( .A1(B[7]), .A2(n79), .B1(C[7]), .B2(n76), .ZN(n141) );
  AOI22_X1 U34 ( .A1(D[16]), .A2(n73), .B1(A[16]), .B2(n2), .ZN(n98) );
  AOI22_X1 U35 ( .A1(B[16]), .A2(n80), .B1(C[16]), .B2(n77), .ZN(n97) );
  AOI22_X1 U36 ( .A1(D[17]), .A2(n73), .B1(A[17]), .B2(n2), .ZN(n100) );
  AOI22_X1 U37 ( .A1(B[17]), .A2(n80), .B1(C[17]), .B2(n77), .ZN(n99) );
  AOI22_X1 U38 ( .A1(D[18]), .A2(n73), .B1(A[18]), .B2(n2), .ZN(n102) );
  AOI22_X1 U39 ( .A1(B[18]), .A2(n80), .B1(C[18]), .B2(n77), .ZN(n101) );
  AOI22_X1 U40 ( .A1(D[19]), .A2(n73), .B1(A[19]), .B2(n2), .ZN(n104) );
  AOI22_X1 U41 ( .A1(B[19]), .A2(n80), .B1(C[19]), .B2(n77), .ZN(n103) );
  AOI22_X1 U42 ( .A1(D[20]), .A2(n73), .B1(A[20]), .B2(n2), .ZN(n108) );
  AOI22_X1 U43 ( .A1(B[20]), .A2(n80), .B1(C[20]), .B2(n77), .ZN(n107) );
  AOI22_X1 U44 ( .A1(D[21]), .A2(n74), .B1(A[21]), .B2(n2), .ZN(n110) );
  AOI22_X1 U45 ( .A1(B[21]), .A2(n80), .B1(C[21]), .B2(n77), .ZN(n109) );
  AOI22_X1 U46 ( .A1(D[22]), .A2(n74), .B1(A[22]), .B2(n2), .ZN(n112) );
  AOI22_X1 U47 ( .A1(B[22]), .A2(n80), .B1(C[22]), .B2(n77), .ZN(n111) );
  AOI22_X1 U48 ( .A1(D[23]), .A2(n74), .B1(A[23]), .B2(n2), .ZN(n114) );
  AOI22_X1 U49 ( .A1(B[23]), .A2(n80), .B1(C[23]), .B2(n77), .ZN(n113) );
  AOI22_X1 U50 ( .A1(D[24]), .A2(n74), .B1(A[24]), .B2(n2), .ZN(n116) );
  AOI22_X1 U51 ( .A1(B[24]), .A2(n80), .B1(C[24]), .B2(n77), .ZN(n115) );
  AOI22_X1 U52 ( .A1(D[25]), .A2(n74), .B1(A[25]), .B2(n2), .ZN(n118) );
  AOI22_X1 U53 ( .A1(B[25]), .A2(n80), .B1(C[25]), .B2(n77), .ZN(n117) );
  AOI22_X1 U54 ( .A1(D[26]), .A2(n74), .B1(A[26]), .B2(n2), .ZN(n120) );
  AOI22_X1 U55 ( .A1(B[26]), .A2(n80), .B1(C[26]), .B2(n77), .ZN(n119) );
  AOI22_X1 U56 ( .A1(D[27]), .A2(n74), .B1(A[27]), .B2(n1), .ZN(n122) );
  AOI22_X1 U57 ( .A1(B[27]), .A2(n79), .B1(C[27]), .B2(n76), .ZN(n121) );
  AOI22_X1 U58 ( .A1(D[28]), .A2(n74), .B1(A[28]), .B2(n1), .ZN(n124) );
  AOI22_X1 U59 ( .A1(B[28]), .A2(n79), .B1(C[28]), .B2(n76), .ZN(n123) );
  AOI22_X1 U60 ( .A1(D[29]), .A2(n74), .B1(A[29]), .B2(n1), .ZN(n126) );
  AOI22_X1 U61 ( .A1(B[29]), .A2(n79), .B1(C[29]), .B2(n76), .ZN(n125) );
  AOI22_X1 U62 ( .A1(D[30]), .A2(n74), .B1(A[30]), .B2(n1), .ZN(n130) );
  AOI22_X1 U63 ( .A1(B[30]), .A2(n79), .B1(C[30]), .B2(n76), .ZN(n129) );
  AOI22_X1 U64 ( .A1(D[31]), .A2(n74), .B1(A[31]), .B2(n1), .ZN(n132) );
  AOI22_X1 U65 ( .A1(B[31]), .A2(n79), .B1(C[31]), .B2(n76), .ZN(n131) );
  AOI22_X1 U66 ( .A1(D[8]), .A2(n75), .B1(A[8]), .B2(n1), .ZN(n144) );
  AOI22_X1 U67 ( .A1(B[8]), .A2(n79), .B1(C[8]), .B2(n76), .ZN(n143) );
  AOI22_X1 U68 ( .A1(D[9]), .A2(n75), .B1(A[9]), .B2(n1), .ZN(n150) );
  AOI22_X1 U69 ( .A1(B[9]), .A2(n79), .B1(C[9]), .B2(n76), .ZN(n149) );
  AOI22_X1 U102 ( .A1(D[10]), .A2(n73), .B1(A[10]), .B2(n72), .ZN(n86) );
  AOI22_X1 U103 ( .A1(B[10]), .A2(n81), .B1(C[10]), .B2(n78), .ZN(n85) );
  AOI22_X1 U104 ( .A1(D[11]), .A2(n73), .B1(A[11]), .B2(n72), .ZN(n88) );
  AOI22_X1 U105 ( .A1(B[11]), .A2(n81), .B1(C[11]), .B2(n78), .ZN(n87) );
  AOI22_X1 U106 ( .A1(D[12]), .A2(n73), .B1(A[12]), .B2(n72), .ZN(n90) );
  AOI22_X1 U107 ( .A1(B[12]), .A2(n81), .B1(C[12]), .B2(n78), .ZN(n89) );
  AOI22_X1 U108 ( .A1(D[13]), .A2(n73), .B1(A[13]), .B2(n72), .ZN(n92) );
  AOI22_X1 U109 ( .A1(B[13]), .A2(n81), .B1(C[13]), .B2(n78), .ZN(n91) );
  AOI22_X1 U110 ( .A1(D[14]), .A2(n73), .B1(A[14]), .B2(n72), .ZN(n94) );
  AOI22_X1 U111 ( .A1(B[14]), .A2(n81), .B1(C[14]), .B2(n78), .ZN(n93) );
  AOI22_X1 U112 ( .A1(D[15]), .A2(n73), .B1(A[15]), .B2(n2), .ZN(n96) );
  AOI22_X1 U113 ( .A1(B[15]), .A2(n80), .B1(C[15]), .B2(n77), .ZN(n95) );
endmodule


module MUX41_GEN_N32_1 ( A, B, C, D, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150;

  NAND2_X1 U70 ( .A1(n150), .A2(n149), .ZN(Y[9]) );
  NAND2_X1 U71 ( .A1(n144), .A2(n143), .ZN(Y[8]) );
  NAND2_X1 U72 ( .A1(n142), .A2(n141), .ZN(Y[7]) );
  NAND2_X1 U73 ( .A1(n140), .A2(n139), .ZN(Y[6]) );
  NAND2_X1 U74 ( .A1(n138), .A2(n137), .ZN(Y[5]) );
  NAND2_X1 U75 ( .A1(n136), .A2(n135), .ZN(Y[4]) );
  NAND2_X1 U76 ( .A1(n134), .A2(n133), .ZN(Y[3]) );
  NAND2_X1 U77 ( .A1(n132), .A2(n131), .ZN(Y[31]) );
  NAND2_X1 U78 ( .A1(n130), .A2(n129), .ZN(Y[30]) );
  NAND2_X1 U79 ( .A1(n128), .A2(n127), .ZN(Y[2]) );
  NAND2_X1 U80 ( .A1(n126), .A2(n125), .ZN(Y[29]) );
  NAND2_X1 U81 ( .A1(n124), .A2(n123), .ZN(Y[28]) );
  NAND2_X1 U82 ( .A1(n122), .A2(n121), .ZN(Y[27]) );
  NAND2_X1 U83 ( .A1(n120), .A2(n119), .ZN(Y[26]) );
  NAND2_X1 U84 ( .A1(n118), .A2(n117), .ZN(Y[25]) );
  NAND2_X1 U85 ( .A1(n116), .A2(n115), .ZN(Y[24]) );
  NAND2_X1 U86 ( .A1(n114), .A2(n113), .ZN(Y[23]) );
  NAND2_X1 U87 ( .A1(n112), .A2(n111), .ZN(Y[22]) );
  NAND2_X1 U88 ( .A1(n110), .A2(n109), .ZN(Y[21]) );
  NAND2_X1 U89 ( .A1(n108), .A2(n107), .ZN(Y[20]) );
  NAND2_X1 U90 ( .A1(n106), .A2(n105), .ZN(Y[1]) );
  NAND2_X1 U91 ( .A1(n104), .A2(n103), .ZN(Y[19]) );
  NAND2_X1 U92 ( .A1(n102), .A2(n101), .ZN(Y[18]) );
  NAND2_X1 U93 ( .A1(n100), .A2(n99), .ZN(Y[17]) );
  NAND2_X1 U94 ( .A1(n98), .A2(n97), .ZN(Y[16]) );
  NAND2_X1 U95 ( .A1(n96), .A2(n95), .ZN(Y[15]) );
  NAND2_X1 U96 ( .A1(n94), .A2(n93), .ZN(Y[14]) );
  NAND2_X1 U97 ( .A1(n92), .A2(n91), .ZN(Y[13]) );
  NAND2_X1 U98 ( .A1(n90), .A2(n89), .ZN(Y[12]) );
  NAND2_X1 U99 ( .A1(n88), .A2(n87), .ZN(Y[11]) );
  NAND2_X1 U100 ( .A1(n86), .A2(n85), .ZN(Y[10]) );
  NAND2_X1 U101 ( .A1(n84), .A2(n83), .ZN(Y[0]) );
  BUF_X1 U1 ( .A(n146), .Z(n73) );
  BUF_X1 U2 ( .A(n146), .Z(n74) );
  BUF_X1 U3 ( .A(n146), .Z(n75) );
  NOR3_X1 U4 ( .A1(n78), .A2(n72), .A3(n81), .ZN(n146) );
  BUF_X1 U5 ( .A(n147), .Z(n78) );
  BUF_X1 U6 ( .A(n148), .Z(n81) );
  BUF_X1 U7 ( .A(n145), .Z(n72) );
  BUF_X1 U8 ( .A(n147), .Z(n77) );
  BUF_X1 U9 ( .A(n147), .Z(n76) );
  BUF_X1 U10 ( .A(n148), .Z(n80) );
  BUF_X1 U11 ( .A(n148), .Z(n79) );
  BUF_X1 U12 ( .A(n145), .Z(n2) );
  BUF_X1 U13 ( .A(n145), .Z(n1) );
  NOR2_X1 U14 ( .A1(n82), .A2(SEL[1]), .ZN(n147) );
  AOI22_X1 U15 ( .A1(B[0]), .A2(n81), .B1(C[0]), .B2(n78), .ZN(n83) );
  AOI22_X1 U16 ( .A1(D[0]), .A2(n73), .B1(A[0]), .B2(n72), .ZN(n84) );
  AOI22_X1 U17 ( .A1(B[1]), .A2(n80), .B1(C[1]), .B2(n77), .ZN(n105) );
  AOI22_X1 U18 ( .A1(D[1]), .A2(n73), .B1(A[1]), .B2(n2), .ZN(n106) );
  AOI22_X1 U19 ( .A1(B[2]), .A2(n79), .B1(C[2]), .B2(n76), .ZN(n127) );
  AOI22_X1 U20 ( .A1(D[2]), .A2(n74), .B1(A[2]), .B2(n1), .ZN(n128) );
  AOI22_X1 U21 ( .A1(B[3]), .A2(n79), .B1(C[3]), .B2(n76), .ZN(n133) );
  AOI22_X1 U22 ( .A1(D[3]), .A2(n74), .B1(A[3]), .B2(n1), .ZN(n134) );
  AOI22_X1 U23 ( .A1(B[4]), .A2(n79), .B1(C[4]), .B2(n76), .ZN(n135) );
  AOI22_X1 U24 ( .A1(D[4]), .A2(n75), .B1(A[4]), .B2(n1), .ZN(n136) );
  AOI22_X1 U25 ( .A1(B[5]), .A2(n79), .B1(C[5]), .B2(n76), .ZN(n137) );
  AOI22_X1 U26 ( .A1(D[5]), .A2(n75), .B1(A[5]), .B2(n1), .ZN(n138) );
  AOI22_X1 U27 ( .A1(B[6]), .A2(n79), .B1(C[6]), .B2(n76), .ZN(n139) );
  AOI22_X1 U28 ( .A1(D[6]), .A2(n75), .B1(A[6]), .B2(n1), .ZN(n140) );
  AOI22_X1 U29 ( .A1(B[7]), .A2(n79), .B1(C[7]), .B2(n76), .ZN(n141) );
  AOI22_X1 U30 ( .A1(D[7]), .A2(n75), .B1(A[7]), .B2(n1), .ZN(n142) );
  AOI22_X1 U31 ( .A1(B[8]), .A2(n79), .B1(C[8]), .B2(n76), .ZN(n143) );
  AOI22_X1 U32 ( .A1(D[8]), .A2(n75), .B1(A[8]), .B2(n1), .ZN(n144) );
  AOI22_X1 U33 ( .A1(B[9]), .A2(n79), .B1(C[9]), .B2(n76), .ZN(n149) );
  AOI22_X1 U34 ( .A1(D[9]), .A2(n75), .B1(A[9]), .B2(n1), .ZN(n150) );
  AOI22_X1 U35 ( .A1(B[10]), .A2(n81), .B1(C[10]), .B2(n78), .ZN(n85) );
  AOI22_X1 U36 ( .A1(D[10]), .A2(n73), .B1(A[10]), .B2(n72), .ZN(n86) );
  AOI22_X1 U37 ( .A1(B[11]), .A2(n81), .B1(C[11]), .B2(n78), .ZN(n87) );
  AOI22_X1 U38 ( .A1(D[11]), .A2(n73), .B1(A[11]), .B2(n72), .ZN(n88) );
  AOI22_X1 U39 ( .A1(B[12]), .A2(n81), .B1(C[12]), .B2(n78), .ZN(n89) );
  AOI22_X1 U40 ( .A1(D[12]), .A2(n73), .B1(A[12]), .B2(n72), .ZN(n90) );
  AOI22_X1 U41 ( .A1(B[13]), .A2(n81), .B1(C[13]), .B2(n78), .ZN(n91) );
  AOI22_X1 U42 ( .A1(D[13]), .A2(n73), .B1(A[13]), .B2(n72), .ZN(n92) );
  AOI22_X1 U43 ( .A1(B[14]), .A2(n81), .B1(C[14]), .B2(n78), .ZN(n93) );
  AOI22_X1 U44 ( .A1(D[14]), .A2(n73), .B1(A[14]), .B2(n72), .ZN(n94) );
  AOI22_X1 U45 ( .A1(B[15]), .A2(n80), .B1(C[15]), .B2(n77), .ZN(n95) );
  AOI22_X1 U46 ( .A1(D[15]), .A2(n73), .B1(A[15]), .B2(n2), .ZN(n96) );
  AOI22_X1 U47 ( .A1(B[16]), .A2(n80), .B1(C[16]), .B2(n77), .ZN(n97) );
  AOI22_X1 U48 ( .A1(D[16]), .A2(n73), .B1(A[16]), .B2(n2), .ZN(n98) );
  AOI22_X1 U49 ( .A1(B[17]), .A2(n80), .B1(C[17]), .B2(n77), .ZN(n99) );
  AOI22_X1 U50 ( .A1(D[17]), .A2(n73), .B1(A[17]), .B2(n2), .ZN(n100) );
  AOI22_X1 U51 ( .A1(B[18]), .A2(n80), .B1(C[18]), .B2(n77), .ZN(n101) );
  AOI22_X1 U52 ( .A1(D[18]), .A2(n73), .B1(A[18]), .B2(n2), .ZN(n102) );
  AOI22_X1 U53 ( .A1(B[19]), .A2(n80), .B1(C[19]), .B2(n77), .ZN(n103) );
  AOI22_X1 U54 ( .A1(D[19]), .A2(n73), .B1(A[19]), .B2(n2), .ZN(n104) );
  AOI22_X1 U55 ( .A1(B[20]), .A2(n80), .B1(C[20]), .B2(n77), .ZN(n107) );
  AOI22_X1 U56 ( .A1(D[20]), .A2(n73), .B1(A[20]), .B2(n2), .ZN(n108) );
  AOI22_X1 U57 ( .A1(B[21]), .A2(n80), .B1(C[21]), .B2(n77), .ZN(n109) );
  AOI22_X1 U58 ( .A1(D[21]), .A2(n74), .B1(A[21]), .B2(n2), .ZN(n110) );
  AOI22_X1 U59 ( .A1(B[22]), .A2(n80), .B1(C[22]), .B2(n77), .ZN(n111) );
  AOI22_X1 U60 ( .A1(D[22]), .A2(n74), .B1(A[22]), .B2(n2), .ZN(n112) );
  AOI22_X1 U61 ( .A1(B[23]), .A2(n80), .B1(C[23]), .B2(n77), .ZN(n113) );
  AOI22_X1 U62 ( .A1(D[23]), .A2(n74), .B1(A[23]), .B2(n2), .ZN(n114) );
  AOI22_X1 U63 ( .A1(B[24]), .A2(n80), .B1(C[24]), .B2(n77), .ZN(n115) );
  AOI22_X1 U64 ( .A1(D[24]), .A2(n74), .B1(A[24]), .B2(n2), .ZN(n116) );
  AOI22_X1 U65 ( .A1(B[25]), .A2(n80), .B1(C[25]), .B2(n77), .ZN(n117) );
  AOI22_X1 U66 ( .A1(D[25]), .A2(n74), .B1(A[25]), .B2(n2), .ZN(n118) );
  AOI22_X1 U67 ( .A1(B[26]), .A2(n80), .B1(C[26]), .B2(n77), .ZN(n119) );
  AOI22_X1 U68 ( .A1(D[26]), .A2(n74), .B1(A[26]), .B2(n2), .ZN(n120) );
  AOI22_X1 U69 ( .A1(B[27]), .A2(n79), .B1(C[27]), .B2(n76), .ZN(n121) );
  AOI22_X1 U102 ( .A1(D[27]), .A2(n74), .B1(A[27]), .B2(n1), .ZN(n122) );
  AOI22_X1 U103 ( .A1(B[28]), .A2(n79), .B1(C[28]), .B2(n76), .ZN(n123) );
  AOI22_X1 U104 ( .A1(D[28]), .A2(n74), .B1(A[28]), .B2(n1), .ZN(n124) );
  AOI22_X1 U105 ( .A1(B[29]), .A2(n79), .B1(C[29]), .B2(n76), .ZN(n125) );
  AOI22_X1 U106 ( .A1(D[29]), .A2(n74), .B1(A[29]), .B2(n1), .ZN(n126) );
  AOI22_X1 U107 ( .A1(B[30]), .A2(n79), .B1(C[30]), .B2(n76), .ZN(n129) );
  AOI22_X1 U108 ( .A1(D[30]), .A2(n74), .B1(A[30]), .B2(n1), .ZN(n130) );
  AOI22_X1 U109 ( .A1(B[31]), .A2(n79), .B1(C[31]), .B2(n76), .ZN(n131) );
  AOI22_X1 U110 ( .A1(D[31]), .A2(n74), .B1(A[31]), .B2(n1), .ZN(n132) );
  AND2_X1 U111 ( .A1(SEL[1]), .A2(n82), .ZN(n148) );
  AND2_X1 U112 ( .A1(SEL[0]), .A2(SEL[1]), .ZN(n145) );
  INV_X1 U113 ( .A(SEL[0]), .ZN(n82) );
endmodule


module CSA_N4_15 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_RCA_1;
  wire   [3:0] S_RCA_2;

  RCA_GEN_N4_30 RCA_1 ( .A(A), .B(B), .Ci(1'b0), .S(S_RCA_1) );
  RCA_GEN_N4_29 RCA_2 ( .A(A), .B(B), .Ci(1'b1), .S(S_RCA_2) );
  MUX21_GEN_N4_15 MUX_SUM ( .A(S_RCA_2), .B(S_RCA_1), .SEL(Ci), .Y(S) );
endmodule


module CSA_N4_14 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_RCA_1;
  wire   [3:0] S_RCA_2;

  RCA_GEN_N4_28 RCA_1 ( .A(A), .B(B), .Ci(1'b0), .S(S_RCA_1) );
  RCA_GEN_N4_27 RCA_2 ( .A(A), .B(B), .Ci(1'b1), .S(S_RCA_2) );
  MUX21_GEN_N4_14 MUX_SUM ( .A(S_RCA_2), .B(S_RCA_1), .SEL(Ci), .Y(S) );
endmodule


module CSA_N4_13 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_RCA_1;
  wire   [3:0] S_RCA_2;

  RCA_GEN_N4_26 RCA_1 ( .A(A), .B(B), .Ci(1'b0), .S(S_RCA_1) );
  RCA_GEN_N4_25 RCA_2 ( .A(A), .B(B), .Ci(1'b1), .S(S_RCA_2) );
  MUX21_GEN_N4_13 MUX_SUM ( .A(S_RCA_2), .B(S_RCA_1), .SEL(Ci), .Y(S) );
endmodule


module CSA_N4_12 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_RCA_1;
  wire   [3:0] S_RCA_2;

  RCA_GEN_N4_24 RCA_1 ( .A(A), .B(B), .Ci(1'b0), .S(S_RCA_1) );
  RCA_GEN_N4_23 RCA_2 ( .A(A), .B(B), .Ci(1'b1), .S(S_RCA_2) );
  MUX21_GEN_N4_12 MUX_SUM ( .A(S_RCA_2), .B(S_RCA_1), .SEL(Ci), .Y(S) );
endmodule


module CSA_N4_11 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_RCA_1;
  wire   [3:0] S_RCA_2;

  RCA_GEN_N4_22 RCA_1 ( .A(A), .B(B), .Ci(1'b0), .S(S_RCA_1) );
  RCA_GEN_N4_21 RCA_2 ( .A(A), .B(B), .Ci(1'b1), .S(S_RCA_2) );
  MUX21_GEN_N4_11 MUX_SUM ( .A(S_RCA_2), .B(S_RCA_1), .SEL(Ci), .Y(S) );
endmodule


module CSA_N4_10 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_RCA_1;
  wire   [3:0] S_RCA_2;

  RCA_GEN_N4_20 RCA_1 ( .A(A), .B(B), .Ci(1'b0), .S(S_RCA_1) );
  RCA_GEN_N4_19 RCA_2 ( .A(A), .B(B), .Ci(1'b1), .S(S_RCA_2) );
  MUX21_GEN_N4_10 MUX_SUM ( .A(S_RCA_2), .B(S_RCA_1), .SEL(Ci), .Y(S) );
endmodule


module CSA_N4_9 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_RCA_1;
  wire   [3:0] S_RCA_2;

  RCA_GEN_N4_18 RCA_1 ( .A(A), .B(B), .Ci(1'b0), .S(S_RCA_1) );
  RCA_GEN_N4_17 RCA_2 ( .A(A), .B(B), .Ci(1'b1), .S(S_RCA_2) );
  MUX21_GEN_N4_9 MUX_SUM ( .A(S_RCA_2), .B(S_RCA_1), .SEL(Ci), .Y(S) );
endmodule


module CSA_N4_8 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_RCA_1;
  wire   [3:0] S_RCA_2;

  RCA_GEN_N4_16 RCA_1 ( .A(A), .B(B), .Ci(1'b0), .S(S_RCA_1) );
  RCA_GEN_N4_15 RCA_2 ( .A(A), .B(B), .Ci(1'b1), .S(S_RCA_2) );
  MUX21_GEN_N4_8 MUX_SUM ( .A(S_RCA_2), .B(S_RCA_1), .SEL(Ci), .Y(S) );
endmodule


module CSA_N4_7 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_RCA_1;
  wire   [3:0] S_RCA_2;

  RCA_GEN_N4_14 RCA_1 ( .A(A), .B(B), .Ci(1'b0), .S(S_RCA_1) );
  RCA_GEN_N4_13 RCA_2 ( .A(A), .B(B), .Ci(1'b1), .S(S_RCA_2) );
  MUX21_GEN_N4_7 MUX_SUM ( .A(S_RCA_2), .B(S_RCA_1), .SEL(Ci), .Y(S) );
endmodule


module CSA_N4_6 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_RCA_1;
  wire   [3:0] S_RCA_2;

  RCA_GEN_N4_12 RCA_1 ( .A(A), .B(B), .Ci(1'b0), .S(S_RCA_1) );
  RCA_GEN_N4_11 RCA_2 ( .A(A), .B(B), .Ci(1'b1), .S(S_RCA_2) );
  MUX21_GEN_N4_6 MUX_SUM ( .A(S_RCA_2), .B(S_RCA_1), .SEL(Ci), .Y(S) );
endmodule


module CSA_N4_5 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_RCA_1;
  wire   [3:0] S_RCA_2;

  RCA_GEN_N4_10 RCA_1 ( .A(A), .B(B), .Ci(1'b0), .S(S_RCA_1) );
  RCA_GEN_N4_9 RCA_2 ( .A(A), .B(B), .Ci(1'b1), .S(S_RCA_2) );
  MUX21_GEN_N4_5 MUX_SUM ( .A(S_RCA_2), .B(S_RCA_1), .SEL(Ci), .Y(S) );
endmodule


module CSA_N4_4 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_RCA_1;
  wire   [3:0] S_RCA_2;

  RCA_GEN_N4_8 RCA_1 ( .A(A), .B(B), .Ci(1'b0), .S(S_RCA_1) );
  RCA_GEN_N4_7 RCA_2 ( .A(A), .B(B), .Ci(1'b1), .S(S_RCA_2) );
  MUX21_GEN_N4_4 MUX_SUM ( .A(S_RCA_2), .B(S_RCA_1), .SEL(Ci), .Y(S) );
endmodule


module CSA_N4_3 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_RCA_1;
  wire   [3:0] S_RCA_2;

  RCA_GEN_N4_6 RCA_1 ( .A(A), .B(B), .Ci(1'b0), .S(S_RCA_1) );
  RCA_GEN_N4_5 RCA_2 ( .A(A), .B(B), .Ci(1'b1), .S(S_RCA_2) );
  MUX21_GEN_N4_3 MUX_SUM ( .A(S_RCA_2), .B(S_RCA_1), .SEL(Ci), .Y(S) );
endmodule


module CSA_N4_2 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_RCA_1;
  wire   [3:0] S_RCA_2;

  RCA_GEN_N4_4 RCA_1 ( .A(A), .B(B), .Ci(1'b0), .S(S_RCA_1) );
  RCA_GEN_N4_3 RCA_2 ( .A(A), .B(B), .Ci(1'b1), .S(S_RCA_2) );
  MUX21_GEN_N4_2 MUX_SUM ( .A(S_RCA_2), .B(S_RCA_1), .SEL(Ci), .Y(S) );
endmodule


module CSA_N4_1 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_RCA_1;
  wire   [3:0] S_RCA_2;

  RCA_GEN_N4_2 RCA_1 ( .A(A), .B(B), .Ci(1'b0), .S(S_RCA_1) );
  RCA_GEN_N4_1 RCA_2 ( .A(A), .B(B), .Ci(1'b1), .S(S_RCA_2) );
  MUX21_GEN_N4_1 MUX_SUM ( .A(S_RCA_2), .B(S_RCA_1), .SEL(Ci), .Y(S) );
endmodule


module AND_GATE_1_737 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_736 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_735 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_734 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_733 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_732 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_731 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_730 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_729 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_728 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_727 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_726 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_725 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_724 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_723 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_722 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_721 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_720 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_719 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_718 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_717 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_716 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_715 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_714 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_713 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_712 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_711 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_710 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_709 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_708 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_707 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_706 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_705 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_704 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_703 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_702 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_701 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_700 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_699 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_698 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_697 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_696 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_695 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_694 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_693 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_692 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_691 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_690 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_689 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_688 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_687 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_686 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_685 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_684 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_683 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_682 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_681 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_680 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_679 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_678 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_677 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_676 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_675 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_674 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_673 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_672 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_671 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_670 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_669 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_668 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_667 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_666 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_665 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_664 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_663 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_662 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_661 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_660 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_659 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_658 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_657 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_656 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_655 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_654 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_653 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_652 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_651 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_650 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_649 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_648 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_647 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_646 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_645 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_644 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_643 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_642 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_641 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_640 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_639 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_638 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_637 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_636 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_635 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_634 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_633 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_632 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_631 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_630 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_629 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_628 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_627 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_626 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_625 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_624 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_623 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_622 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_621 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_620 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_619 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_618 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_617 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_616 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_615 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_614 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_613 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_612 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_611 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_610 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_609 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_608 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_607 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_606 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_605 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_604 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_603 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_602 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_601 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_600 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_599 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_598 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_597 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_596 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_595 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_594 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_593 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_592 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_591 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_590 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_589 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_588 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_587 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_586 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_585 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_584 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_583 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_582 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_581 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_580 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_579 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_578 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_577 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_576 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_575 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_574 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_573 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_572 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_571 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_570 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_569 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_568 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_567 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_566 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_565 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_564 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_563 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_562 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_561 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_560 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_559 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_558 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_557 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_556 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_555 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_554 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_553 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_552 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_551 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_550 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_549 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_548 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_547 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_546 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_545 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_544 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_543 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_542 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_541 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_540 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_539 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_538 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_537 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_536 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_535 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_534 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_533 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_532 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_531 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_530 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_529 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_528 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_527 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_526 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_525 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_524 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_523 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_522 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_521 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_520 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_519 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_518 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_517 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_516 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_515 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_514 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_513 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_512 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_511 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_510 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_509 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_508 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_507 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_506 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_505 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_504 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_503 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_502 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_501 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_500 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_499 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_498 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_497 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_496 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_495 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_494 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_493 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_492 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_491 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_490 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_489 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_488 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_487 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_486 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_485 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_484 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_483 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_482 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_481 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_480 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_479 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_478 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_477 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_476 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_475 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_474 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_473 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_472 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_471 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_470 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_469 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_468 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_467 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_466 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_465 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_464 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_463 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_462 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_461 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_460 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_459 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_458 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_457 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_456 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_455 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_454 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_453 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_452 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_451 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_450 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_449 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_448 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_447 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_446 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_445 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_444 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_443 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_442 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_441 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_440 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_439 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_438 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_437 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_436 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_435 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_434 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_433 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_432 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_431 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_430 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_429 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_428 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_427 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_426 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_425 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_424 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_423 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_422 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_421 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_420 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_419 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_418 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_417 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_416 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_415 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_414 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_413 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_412 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_411 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_410 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_409 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_408 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_407 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_406 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_405 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_404 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_403 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_402 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_401 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_400 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_399 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_398 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_397 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_396 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_395 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_394 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_393 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_392 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_391 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_390 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_389 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_388 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_387 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_386 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_385 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_384 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_383 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_382 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_381 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_380 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_379 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_378 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_377 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_376 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_375 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_374 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_373 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_372 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_371 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_370 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_369 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_368 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_367 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_366 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_365 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_364 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_363 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_362 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_361 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_360 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_359 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_358 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_357 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_356 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_355 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_354 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_353 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_352 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_351 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_350 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_349 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_348 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_347 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_346 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_345 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_344 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_343 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_342 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_341 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_340 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_339 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1;

  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Y) );
endmodule


module AND_GATE_1_338 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_337 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_336 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_335 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_334 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_333 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_332 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_331 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_330 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_329 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_328 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_327 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_326 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_325 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_324 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_323 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_322 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_321 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_320 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_319 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_318 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_317 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_316 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_315 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_314 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_313 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_312 ( A, B, Y );
  input A, B;
  output Y;
  wire   n1;

  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Y) );
endmodule


module AND_GATE_1_311 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_310 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_309 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_308 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_307 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_306 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_305 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_304 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_303 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_302 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_301 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_300 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_299 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_298 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_297 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_296 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_295 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_294 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_293 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_292 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_291 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_290 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_289 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_288 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_287 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_286 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_285 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_284 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_283 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_282 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_281 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_280 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_279 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_278 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_277 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_276 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_275 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_274 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_273 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_272 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_271 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_270 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_269 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_268 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_267 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_266 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_265 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_264 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_263 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_262 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_261 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_260 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_259 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_258 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_257 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_256 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_255 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_254 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_253 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_252 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_251 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_250 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_249 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_248 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_247 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_246 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_245 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_244 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_243 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_242 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_241 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_240 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_239 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_238 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_237 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_236 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_235 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_234 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_233 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_232 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_231 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_230 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_229 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_228 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_227 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_226 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_225 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_224 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_223 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_222 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_221 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_220 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_219 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_218 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_217 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_216 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_215 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_214 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_213 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_212 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_211 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_210 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_209 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_208 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_207 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_206 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_205 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_204 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_203 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_202 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_201 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_200 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_199 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_198 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_197 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_196 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_195 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_194 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_193 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_192 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_191 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_190 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_189 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_188 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_187 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_186 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_185 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_184 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_183 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_182 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_181 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_180 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_179 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_178 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_177 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_176 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_175 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_174 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_173 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_172 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_171 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_170 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_169 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_168 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_167 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_166 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_165 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_164 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_163 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_162 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_161 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module AND_GATE_1_160 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_159 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_158 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_157 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_156 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_155 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_154 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_153 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_152 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_151 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_150 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_149 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_148 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_147 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_146 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_145 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_144 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_143 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_142 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_141 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_140 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_139 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_138 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_137 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_136 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_135 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_134 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_133 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_132 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_131 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X4 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_130 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_129 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_128 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_127 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_126 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_125 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_124 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_123 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_122 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_121 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_120 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_119 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_118 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_117 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_116 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_115 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_114 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_113 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_112 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_111 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_110 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_109 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_108 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_107 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_106 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_105 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_104 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_103 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_102 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_101 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_100 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_99 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_98 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_97 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_96 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_95 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_94 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_93 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_92 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_91 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_90 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_89 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_88 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_87 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_86 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_85 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_84 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_83 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_82 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_81 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_80 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_79 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_78 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_77 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_76 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_75 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_74 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_73 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_72 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_71 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_70 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_69 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_68 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_67 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_66 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_65 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_64 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_63 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_62 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_61 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_60 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_59 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_58 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_57 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_56 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_55 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_54 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_53 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_52 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_51 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_50 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_49 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_48 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_47 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_46 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_45 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_44 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_43 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_42 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_41 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_40 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_39 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_38 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_37 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_36 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_35 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_34 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_33 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_32 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_31 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_30 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_29 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_28 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_27 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_26 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_25 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_24 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_23 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_22 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_21 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_20 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_19 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_18 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_17 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_16 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_15 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_14 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_13 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_12 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_11 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_10 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_9 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_8 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_7 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_6 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_5 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_4 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_3 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_2 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1_1 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module FD_1_581 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_580 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_579 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_578 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_577 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_576 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_575 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_574 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_573 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_572 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_571 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_570 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_569 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_568 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_567 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_566 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_565 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_564 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_563 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_562 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_561 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_560 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_559 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_558 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_557 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_556 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_555 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_554 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_553 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_552 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_551 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_550 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_549 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n2, n3;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  AND2_X1 U3 ( .A1(n2), .A2(n3), .ZN(n1) );
  INV_X1 U4 ( .A(RST), .ZN(n2) );
  MUX2_X1 U5 ( .A(Q), .B(D), .S(EN), .Z(n3) );
endmodule


module FD_1_548 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_547 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_546 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_545 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_544 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_543 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_542 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_541 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_540 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_539 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_538 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_537 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_536 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_535 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_534 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_533 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_532 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_531 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_530 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_529 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_528 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_527 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_526 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_525 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_524 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_523 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_522 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_521 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_520 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_519 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_518 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_517 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_516 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_515 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_514 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_513 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_512 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_511 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_510 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_509 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_508 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_507 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_506 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_505 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_504 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_503 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_502 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_501 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_500 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_499 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_498 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_497 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_496 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_495 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_494 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_493 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_492 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_491 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_490 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_489 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_488 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_487 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_486 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_485 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_484 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_483 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_482 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_481 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_480 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_479 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_478 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_477 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_476 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_475 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_474 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_473 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_472 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_471 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_470 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_469 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_468 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_467 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_466 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_465 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_464 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_463 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_462 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_461 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_460 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_459 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_458 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_457 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_456 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_455 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_454 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_453 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_452 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_451 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_450 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_449 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_448 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_447 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_446 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_445 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_444 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_443 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_442 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_441 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_440 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_439 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_438 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_437 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_436 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_435 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_434 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_433 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_432 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_431 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_430 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_429 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_428 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_427 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_426 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_425 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_424 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_423 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_422 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_421 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_420 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_419 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_418 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_417 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_416 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_415 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_414 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_413 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_412 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_411 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_410 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_409 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_408 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_407 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_406 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_405 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_404 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_403 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_402 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_401 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_400 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_399 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_398 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_397 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_396 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_395 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_394 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_393 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_392 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_391 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_390 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_389 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_388 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_387 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_386 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_385 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_384 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_383 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_382 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_381 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_380 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_379 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_378 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  AOI22_X1 U3 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  NOR2_X1 U4 ( .A1(RST), .A2(n4), .ZN(n3) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_377 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_376 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_375 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_374 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_373 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_372 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_371 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_370 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_369 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_368 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_367 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_366 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_365 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_364 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_363 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_362 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_361 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_360 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_359 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_358 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_357 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_356 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_355 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_354 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_353 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_352 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_351 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_350 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_349 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_348 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  AOI22_X2 U3 ( .A1(D), .A2(EN), .B1(Q), .B2(n1), .ZN(n4) );
  NOR2_X1 U4 ( .A1(n4), .A2(RST), .ZN(n3) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_347 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  AOI22_X2 U3 ( .A1(D), .A2(EN), .B1(Q), .B2(n1), .ZN(n4) );
  NOR2_X1 U4 ( .A1(n4), .A2(RST), .ZN(n3) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_346 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_345 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_344 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_343 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_342 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_341 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_340 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_339 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_338 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_337 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_336 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_335 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_334 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_333 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_332 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_331 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_330 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_329 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_328 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_327 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_326 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_325 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_324 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_323 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_322 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_321 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_320 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_319 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_318 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_317 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_316 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_315 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_314 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_313 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_312 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_311 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_310 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_309 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_308 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_307 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_306 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_305 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_304 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_303 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_302 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_301 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_300 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_299 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_298 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_297 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_296 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_295 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_294 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_293 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_292 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_291 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_290 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_289 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_288 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_287 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_286 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_285 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_284 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_283 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_282 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_281 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_280 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_279 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_278 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_277 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_276 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_275 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_274 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_273 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_272 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_271 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_270 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_269 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_268 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_267 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_266 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_265 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_264 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_263 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_262 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_261 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_260 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_259 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_258 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_257 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_256 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_255 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_254 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_253 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_252 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_251 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_250 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_249 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_248 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_247 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_246 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_245 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_244 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_243 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_242 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_241 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_240 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_239 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_238 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_237 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_236 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_235 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_234 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_233 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_232 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_231 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_230 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_229 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_228 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_227 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_226 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_225 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_224 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_223 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_222 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_221 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_220 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_219 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_218 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_217 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_216 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_215 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_214 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_213 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_212 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_211 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_210 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_209 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_208 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_207 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_206 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_205 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_204 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_203 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_202 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_201 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_200 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_199 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_198 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_197 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_196 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_195 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_194 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_193 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_192 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_191 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_190 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_189 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_188 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_187 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_186 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_185 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_184 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_183 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_182 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_181 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_180 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_179 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_178 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_177 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_176 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_175 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_174 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_173 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_172 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_171 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_170 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_169 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_168 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_167 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_166 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_165 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_164 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_163 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_162 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_161 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_160 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_159 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_158 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_157 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_156 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_155 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_154 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_153 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_152 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_151 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_150 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_149 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_148 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_147 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_146 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_145 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n8, n1, n4, n6, n7;

  DFF_X1 Q_reg ( .D(n6), .CK(CLK), .Q(n8), .QN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(Q) );
  NOR2_X1 U4 ( .A1(RST), .A2(n7), .ZN(n6) );
  AOI22_X1 U5 ( .A1(EN), .A2(D), .B1(n8), .B2(n4), .ZN(n7) );
  INV_X1 U6 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_144 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n8, n1, n4, n6, n7;

  DFF_X1 Q_reg ( .D(n6), .CK(CLK), .Q(n8), .QN(n1) );
  INV_X2 U3 ( .A(n1), .ZN(Q) );
  NOR2_X1 U4 ( .A1(RST), .A2(n7), .ZN(n6) );
  AOI22_X1 U5 ( .A1(EN), .A2(D), .B1(n8), .B2(n4), .ZN(n7) );
  INV_X1 U6 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_143 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_142 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_141 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_140 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_139 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n6, n1, n4, n5;

  DFF_X1 Q_reg ( .D(n4), .CK(CLK), .Q(n6) );
  BUF_X1 U3 ( .A(n6), .Z(Q) );
  NOR2_X1 U4 ( .A1(RST), .A2(n5), .ZN(n4) );
  AOI22_X1 U5 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n5) );
  INV_X1 U6 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_138 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_137 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_136 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_135 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_134 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_133 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_132 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_131 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_130 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_129 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_128 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_127 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_126 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_125 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_124 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_123 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_122 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_121 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_120 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_119 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_118 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n2, n3;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  AND2_X1 U3 ( .A1(n2), .A2(n3), .ZN(n1) );
  INV_X1 U4 ( .A(RST), .ZN(n2) );
  MUX2_X1 U5 ( .A(Q), .B(D), .S(EN), .Z(n3) );
endmodule


module FD_1_117 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n2, n3;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  AND2_X1 U3 ( .A1(n2), .A2(n3), .ZN(n1) );
  INV_X1 U4 ( .A(RST), .ZN(n2) );
  MUX2_X1 U5 ( .A(Q), .B(D), .S(EN), .Z(n3) );
endmodule


module FD_1_116 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n2, n3, n4, n5, n6;

  DFF_X1 Q_reg ( .D(n4), .CK(CLK), .Q(Q) );
  NAND2_X1 U3 ( .A1(Q), .A2(n1), .ZN(n2) );
  NAND2_X1 U4 ( .A1(D), .A2(EN), .ZN(n3) );
  NAND2_X1 U5 ( .A1(n2), .A2(n3), .ZN(n6) );
  INV_X1 U6 ( .A(EN), .ZN(n1) );
  AND2_X2 U7 ( .A1(n5), .A2(n6), .ZN(n4) );
  INV_X1 U8 ( .A(RST), .ZN(n5) );
endmodule


module FD_1_115 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_114 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_113 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_112 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_111 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_110 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_109 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_108 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_107 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_106 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_105 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_104 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_103 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_102 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_101 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_100 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_99 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_98 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_97 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_96 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_95 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_94 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_93 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_92 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_91 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_90 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_89 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_88 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_87 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_86 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_85 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_84 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_83 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_82 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_81 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_80 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_79 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_78 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_77 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_76 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_75 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_74 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_73 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_72 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_71 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_70 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_69 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_68 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_67 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_66 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1_65 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_64 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_63 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_62 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_61 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_60 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_59 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_58 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_57 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_56 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_55 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_54 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_53 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_52 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_51 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_50 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_49 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_48 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_47 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_46 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_45 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_44 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_43 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_42 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_41 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_40 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_39 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_38 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_37 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_36 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_35 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_34 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_33 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_32 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_31 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_30 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_29 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_28 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_27 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_26 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_25 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_24 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_23 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_22 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_21 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_20 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_19 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_18 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_17 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_16 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_15 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_14 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_13 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_12 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_11 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_10 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_9 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_8 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_7 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_6 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_5 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_4 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_3 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_2 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_1_1 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module MUX21_GEN_N32_7 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  INV_1_127 UIV ( .A(n1), .Y(SB) );
  NAND_GATE_1518 UND1_0 ( .A(A[0]), .B(n3), .Y(Y1[0]) );
  NAND_GATE_1517 UND2_0 ( .A(B[0]), .B(n6), .Y(Y2[0]) );
  NAND_GATE_1516 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_1515 UND1_1 ( .A(A[1]), .B(n3), .Y(Y1[1]) );
  NAND_GATE_1514 UND2_1 ( .A(B[1]), .B(n6), .Y(Y2[1]) );
  NAND_GATE_1513 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_1512 UND1_2 ( .A(A[2]), .B(n3), .Y(Y1[2]) );
  NAND_GATE_1511 UND2_2 ( .A(B[2]), .B(n6), .Y(Y2[2]) );
  NAND_GATE_1510 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_1509 UND1_3 ( .A(A[3]), .B(n3), .Y(Y1[3]) );
  NAND_GATE_1508 UND2_3 ( .A(B[3]), .B(n6), .Y(Y2[3]) );
  NAND_GATE_1507 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_1506 UND1_4 ( .A(A[4]), .B(n3), .Y(Y1[4]) );
  NAND_GATE_1505 UND2_4 ( .A(B[4]), .B(n6), .Y(Y2[4]) );
  NAND_GATE_1504 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_1503 UND1_5 ( .A(A[5]), .B(n3), .Y(Y1[5]) );
  NAND_GATE_1502 UND2_5 ( .A(B[5]), .B(n6), .Y(Y2[5]) );
  NAND_GATE_1501 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_1500 UND1_6 ( .A(A[6]), .B(n3), .Y(Y1[6]) );
  NAND_GATE_1499 UND2_6 ( .A(B[6]), .B(n5), .Y(Y2[6]) );
  NAND_GATE_1498 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_1497 UND1_7 ( .A(A[7]), .B(n2), .Y(Y1[7]) );
  NAND_GATE_1496 UND2_7 ( .A(B[7]), .B(n5), .Y(Y2[7]) );
  NAND_GATE_1495 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  NAND_GATE_1494 UND1_8 ( .A(A[8]), .B(n2), .Y(Y1[8]) );
  NAND_GATE_1493 UND2_8 ( .A(B[8]), .B(n5), .Y(Y2[8]) );
  NAND_GATE_1492 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  NAND_GATE_1491 UND1_9 ( .A(A[9]), .B(n2), .Y(Y1[9]) );
  NAND_GATE_1490 UND2_9 ( .A(B[9]), .B(n5), .Y(Y2[9]) );
  NAND_GATE_1489 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  NAND_GATE_1488 UND1_10 ( .A(A[10]), .B(n2), .Y(Y1[10]) );
  NAND_GATE_1487 UND2_10 ( .A(B[10]), .B(n5), .Y(Y2[10]) );
  NAND_GATE_1486 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  NAND_GATE_1485 UND1_11 ( .A(A[11]), .B(n2), .Y(Y1[11]) );
  NAND_GATE_1484 UND2_11 ( .A(B[11]), .B(n5), .Y(Y2[11]) );
  NAND_GATE_1483 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  NAND_GATE_1482 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  NAND_GATE_1481 UND2_12 ( .A(B[12]), .B(n5), .Y(Y2[12]) );
  NAND_GATE_1480 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  NAND_GATE_1479 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  NAND_GATE_1478 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  NAND_GATE_1477 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  NAND_GATE_1476 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  NAND_GATE_1475 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  NAND_GATE_1474 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  NAND_GATE_1473 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  NAND_GATE_1472 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  NAND_GATE_1471 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  NAND_GATE_1470 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  NAND_GATE_1469 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  NAND_GATE_1468 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  NAND_GATE_1467 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  NAND_GATE_1466 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  NAND_GATE_1465 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  NAND_GATE_1464 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  NAND_GATE_1463 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  NAND_GATE_1462 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  NAND_GATE_1461 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  NAND_GATE_1460 UND2_19 ( .A(B[19]), .B(n4), .Y(Y2[19]) );
  NAND_GATE_1459 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  NAND_GATE_1458 UND1_20 ( .A(A[20]), .B(n1), .Y(Y1[20]) );
  NAND_GATE_1457 UND2_20 ( .A(B[20]), .B(n4), .Y(Y2[20]) );
  NAND_GATE_1456 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  NAND_GATE_1455 UND1_21 ( .A(A[21]), .B(n1), .Y(Y1[21]) );
  NAND_GATE_1454 UND2_21 ( .A(B[21]), .B(n4), .Y(Y2[21]) );
  NAND_GATE_1453 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  NAND_GATE_1452 UND1_22 ( .A(A[22]), .B(n1), .Y(Y1[22]) );
  NAND_GATE_1451 UND2_22 ( .A(B[22]), .B(n4), .Y(Y2[22]) );
  NAND_GATE_1450 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  NAND_GATE_1449 UND1_23 ( .A(A[23]), .B(n1), .Y(Y1[23]) );
  NAND_GATE_1448 UND2_23 ( .A(B[23]), .B(n4), .Y(Y2[23]) );
  NAND_GATE_1447 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  NAND_GATE_1446 UND1_24 ( .A(A[24]), .B(n1), .Y(Y1[24]) );
  NAND_GATE_1445 UND2_24 ( .A(B[24]), .B(n4), .Y(Y2[24]) );
  NAND_GATE_1444 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  NAND_GATE_1443 UND1_25 ( .A(A[25]), .B(n1), .Y(Y1[25]) );
  NAND_GATE_1442 UND2_25 ( .A(B[25]), .B(n4), .Y(Y2[25]) );
  NAND_GATE_1441 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  NAND_GATE_1440 UND1_26 ( .A(A[26]), .B(n1), .Y(Y1[26]) );
  NAND_GATE_1439 UND2_26 ( .A(B[26]), .B(n4), .Y(Y2[26]) );
  NAND_GATE_1438 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  NAND_GATE_1437 UND1_27 ( .A(A[27]), .B(n1), .Y(Y1[27]) );
  NAND_GATE_1436 UND2_27 ( .A(B[27]), .B(n4), .Y(Y2[27]) );
  NAND_GATE_1435 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  NAND_GATE_1434 UND1_28 ( .A(A[28]), .B(n1), .Y(Y1[28]) );
  NAND_GATE_1433 UND2_28 ( .A(B[28]), .B(n4), .Y(Y2[28]) );
  NAND_GATE_1432 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  NAND_GATE_1431 UND1_29 ( .A(A[29]), .B(n1), .Y(Y1[29]) );
  NAND_GATE_1430 UND2_29 ( .A(B[29]), .B(n4), .Y(Y2[29]) );
  NAND_GATE_1429 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  NAND_GATE_1428 UND1_30 ( .A(A[30]), .B(n1), .Y(Y1[30]) );
  NAND_GATE_1427 UND2_30 ( .A(B[30]), .B(n4), .Y(Y2[30]) );
  NAND_GATE_1426 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  NAND_GATE_1425 UND1_31 ( .A(A[31]), .B(n1), .Y(Y1[31]) );
  NAND_GATE_1424 UND2_31 ( .A(B[31]), .B(n4), .Y(Y2[31]) );
  NAND_GATE_1423 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  BUF_X1 U1 ( .A(SB), .Z(n4) );
  BUF_X1 U2 ( .A(SB), .Z(n5) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GEN_N32_6 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  INV_1_126 UIV ( .A(n1), .Y(SB) );
  NAND_GATE_1422 UND1_0 ( .A(A[0]), .B(n3), .Y(Y1[0]) );
  NAND_GATE_1421 UND2_0 ( .A(B[0]), .B(n6), .Y(Y2[0]) );
  NAND_GATE_1420 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_1419 UND1_1 ( .A(A[1]), .B(n3), .Y(Y1[1]) );
  NAND_GATE_1418 UND2_1 ( .A(B[1]), .B(n6), .Y(Y2[1]) );
  NAND_GATE_1417 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_1416 UND1_2 ( .A(A[2]), .B(n3), .Y(Y1[2]) );
  NAND_GATE_1415 UND2_2 ( .A(B[2]), .B(n6), .Y(Y2[2]) );
  NAND_GATE_1414 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_1413 UND1_3 ( .A(A[3]), .B(n3), .Y(Y1[3]) );
  NAND_GATE_1412 UND2_3 ( .A(B[3]), .B(n6), .Y(Y2[3]) );
  NAND_GATE_1411 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_1410 UND1_4 ( .A(A[4]), .B(n3), .Y(Y1[4]) );
  NAND_GATE_1409 UND2_4 ( .A(B[4]), .B(n6), .Y(Y2[4]) );
  NAND_GATE_1408 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_1407 UND1_5 ( .A(A[5]), .B(n3), .Y(Y1[5]) );
  NAND_GATE_1406 UND2_5 ( .A(B[5]), .B(n6), .Y(Y2[5]) );
  NAND_GATE_1405 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_1404 UND1_6 ( .A(A[6]), .B(n3), .Y(Y1[6]) );
  NAND_GATE_1403 UND2_6 ( .A(B[6]), .B(n5), .Y(Y2[6]) );
  NAND_GATE_1402 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_1401 UND1_7 ( .A(A[7]), .B(n2), .Y(Y1[7]) );
  NAND_GATE_1400 UND2_7 ( .A(B[7]), .B(n5), .Y(Y2[7]) );
  NAND_GATE_1399 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  NAND_GATE_1398 UND1_8 ( .A(A[8]), .B(n2), .Y(Y1[8]) );
  NAND_GATE_1397 UND2_8 ( .A(B[8]), .B(n5), .Y(Y2[8]) );
  NAND_GATE_1396 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  NAND_GATE_1395 UND1_9 ( .A(A[9]), .B(n2), .Y(Y1[9]) );
  NAND_GATE_1394 UND2_9 ( .A(B[9]), .B(n5), .Y(Y2[9]) );
  NAND_GATE_1393 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  NAND_GATE_1392 UND1_10 ( .A(A[10]), .B(n2), .Y(Y1[10]) );
  NAND_GATE_1391 UND2_10 ( .A(B[10]), .B(n5), .Y(Y2[10]) );
  NAND_GATE_1390 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  NAND_GATE_1389 UND1_11 ( .A(A[11]), .B(n2), .Y(Y1[11]) );
  NAND_GATE_1388 UND2_11 ( .A(B[11]), .B(n5), .Y(Y2[11]) );
  NAND_GATE_1387 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  NAND_GATE_1386 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  NAND_GATE_1385 UND2_12 ( .A(B[12]), .B(n5), .Y(Y2[12]) );
  NAND_GATE_1384 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  NAND_GATE_1383 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  NAND_GATE_1382 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  NAND_GATE_1381 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  NAND_GATE_1380 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  NAND_GATE_1379 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  NAND_GATE_1378 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  NAND_GATE_1377 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  NAND_GATE_1376 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  NAND_GATE_1375 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  NAND_GATE_1374 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  NAND_GATE_1373 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  NAND_GATE_1372 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  NAND_GATE_1371 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  NAND_GATE_1370 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  NAND_GATE_1369 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  NAND_GATE_1368 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  NAND_GATE_1367 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  NAND_GATE_1366 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  NAND_GATE_1365 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  NAND_GATE_1364 UND2_19 ( .A(B[19]), .B(n4), .Y(Y2[19]) );
  NAND_GATE_1363 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  NAND_GATE_1362 UND1_20 ( .A(A[20]), .B(n1), .Y(Y1[20]) );
  NAND_GATE_1361 UND2_20 ( .A(B[20]), .B(n4), .Y(Y2[20]) );
  NAND_GATE_1360 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  NAND_GATE_1359 UND1_21 ( .A(A[21]), .B(n1), .Y(Y1[21]) );
  NAND_GATE_1358 UND2_21 ( .A(B[21]), .B(n4), .Y(Y2[21]) );
  NAND_GATE_1357 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  NAND_GATE_1356 UND1_22 ( .A(A[22]), .B(n1), .Y(Y1[22]) );
  NAND_GATE_1355 UND2_22 ( .A(B[22]), .B(n4), .Y(Y2[22]) );
  NAND_GATE_1354 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  NAND_GATE_1353 UND1_23 ( .A(A[23]), .B(n1), .Y(Y1[23]) );
  NAND_GATE_1352 UND2_23 ( .A(B[23]), .B(n4), .Y(Y2[23]) );
  NAND_GATE_1351 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  NAND_GATE_1350 UND1_24 ( .A(A[24]), .B(n1), .Y(Y1[24]) );
  NAND_GATE_1349 UND2_24 ( .A(B[24]), .B(n4), .Y(Y2[24]) );
  NAND_GATE_1348 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  NAND_GATE_1347 UND1_25 ( .A(A[25]), .B(n1), .Y(Y1[25]) );
  NAND_GATE_1346 UND2_25 ( .A(B[25]), .B(n4), .Y(Y2[25]) );
  NAND_GATE_1345 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  NAND_GATE_1344 UND1_26 ( .A(A[26]), .B(n1), .Y(Y1[26]) );
  NAND_GATE_1343 UND2_26 ( .A(B[26]), .B(n4), .Y(Y2[26]) );
  NAND_GATE_1342 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  NAND_GATE_1341 UND1_27 ( .A(A[27]), .B(n1), .Y(Y1[27]) );
  NAND_GATE_1340 UND2_27 ( .A(B[27]), .B(n4), .Y(Y2[27]) );
  NAND_GATE_1339 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  NAND_GATE_1338 UND1_28 ( .A(A[28]), .B(n1), .Y(Y1[28]) );
  NAND_GATE_1337 UND2_28 ( .A(B[28]), .B(n4), .Y(Y2[28]) );
  NAND_GATE_1336 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  NAND_GATE_1335 UND1_29 ( .A(A[29]), .B(n1), .Y(Y1[29]) );
  NAND_GATE_1334 UND2_29 ( .A(B[29]), .B(n4), .Y(Y2[29]) );
  NAND_GATE_1333 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  NAND_GATE_1332 UND1_30 ( .A(A[30]), .B(n1), .Y(Y1[30]) );
  NAND_GATE_1331 UND2_30 ( .A(B[30]), .B(n4), .Y(Y2[30]) );
  NAND_GATE_1330 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  NAND_GATE_1329 UND1_31 ( .A(A[31]), .B(n1), .Y(Y1[31]) );
  NAND_GATE_1328 UND2_31 ( .A(B[31]), .B(n4), .Y(Y2[31]) );
  NAND_GATE_1327 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  BUF_X1 U1 ( .A(SB), .Z(n4) );
  BUF_X1 U2 ( .A(SB), .Z(n5) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n3) );
  BUF_X1 U5 ( .A(SEL), .Z(n1) );
  BUF_X1 U6 ( .A(SEL), .Z(n2) );
endmodule


module MUX21_GEN_N32_5 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  INV_1_125 UIV ( .A(n1), .Y(SB) );
  NAND_GATE_1326 UND1_0 ( .A(A[0]), .B(n3), .Y(Y1[0]) );
  NAND_GATE_1325 UND2_0 ( .A(B[0]), .B(n6), .Y(Y2[0]) );
  NAND_GATE_1324 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_1323 UND1_1 ( .A(A[1]), .B(n3), .Y(Y1[1]) );
  NAND_GATE_1322 UND2_1 ( .A(B[1]), .B(n6), .Y(Y2[1]) );
  NAND_GATE_1321 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_1320 UND1_2 ( .A(A[2]), .B(n3), .Y(Y1[2]) );
  NAND_GATE_1319 UND2_2 ( .A(B[2]), .B(n6), .Y(Y2[2]) );
  NAND_GATE_1318 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_1317 UND1_3 ( .A(A[3]), .B(n3), .Y(Y1[3]) );
  NAND_GATE_1316 UND2_3 ( .A(B[3]), .B(n6), .Y(Y2[3]) );
  NAND_GATE_1315 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_1314 UND1_4 ( .A(A[4]), .B(n3), .Y(Y1[4]) );
  NAND_GATE_1313 UND2_4 ( .A(B[4]), .B(n6), .Y(Y2[4]) );
  NAND_GATE_1312 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_1311 UND1_5 ( .A(A[5]), .B(n3), .Y(Y1[5]) );
  NAND_GATE_1310 UND2_5 ( .A(B[5]), .B(n6), .Y(Y2[5]) );
  NAND_GATE_1309 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_1308 UND1_6 ( .A(A[6]), .B(n3), .Y(Y1[6]) );
  NAND_GATE_1307 UND2_6 ( .A(B[6]), .B(n5), .Y(Y2[6]) );
  NAND_GATE_1306 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_1305 UND1_7 ( .A(A[7]), .B(n2), .Y(Y1[7]) );
  NAND_GATE_1304 UND2_7 ( .A(B[7]), .B(n5), .Y(Y2[7]) );
  NAND_GATE_1303 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  NAND_GATE_1302 UND1_8 ( .A(A[8]), .B(n2), .Y(Y1[8]) );
  NAND_GATE_1301 UND2_8 ( .A(B[8]), .B(n5), .Y(Y2[8]) );
  NAND_GATE_1300 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  NAND_GATE_1299 UND1_9 ( .A(A[9]), .B(n2), .Y(Y1[9]) );
  NAND_GATE_1298 UND2_9 ( .A(B[9]), .B(n5), .Y(Y2[9]) );
  NAND_GATE_1297 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  NAND_GATE_1296 UND1_10 ( .A(A[10]), .B(n2), .Y(Y1[10]) );
  NAND_GATE_1295 UND2_10 ( .A(B[10]), .B(n5), .Y(Y2[10]) );
  NAND_GATE_1294 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  NAND_GATE_1293 UND1_11 ( .A(A[11]), .B(n2), .Y(Y1[11]) );
  NAND_GATE_1292 UND2_11 ( .A(B[11]), .B(n5), .Y(Y2[11]) );
  NAND_GATE_1291 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  NAND_GATE_1290 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  NAND_GATE_1289 UND2_12 ( .A(B[12]), .B(n5), .Y(Y2[12]) );
  NAND_GATE_1288 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  NAND_GATE_1287 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  NAND_GATE_1286 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  NAND_GATE_1285 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  NAND_GATE_1284 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  NAND_GATE_1283 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  NAND_GATE_1282 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  NAND_GATE_1281 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  NAND_GATE_1280 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  NAND_GATE_1279 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  NAND_GATE_1278 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  NAND_GATE_1277 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  NAND_GATE_1276 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  NAND_GATE_1275 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  NAND_GATE_1274 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  NAND_GATE_1273 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  NAND_GATE_1272 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  NAND_GATE_1271 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  NAND_GATE_1270 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  NAND_GATE_1269 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  NAND_GATE_1268 UND2_19 ( .A(B[19]), .B(n4), .Y(Y2[19]) );
  NAND_GATE_1267 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  NAND_GATE_1266 UND1_20 ( .A(A[20]), .B(n1), .Y(Y1[20]) );
  NAND_GATE_1265 UND2_20 ( .A(B[20]), .B(n4), .Y(Y2[20]) );
  NAND_GATE_1264 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  NAND_GATE_1263 UND1_21 ( .A(A[21]), .B(n1), .Y(Y1[21]) );
  NAND_GATE_1262 UND2_21 ( .A(B[21]), .B(n4), .Y(Y2[21]) );
  NAND_GATE_1261 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  NAND_GATE_1260 UND1_22 ( .A(A[22]), .B(n1), .Y(Y1[22]) );
  NAND_GATE_1259 UND2_22 ( .A(B[22]), .B(n4), .Y(Y2[22]) );
  NAND_GATE_1258 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  NAND_GATE_1257 UND1_23 ( .A(A[23]), .B(n1), .Y(Y1[23]) );
  NAND_GATE_1256 UND2_23 ( .A(B[23]), .B(n4), .Y(Y2[23]) );
  NAND_GATE_1255 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  NAND_GATE_1254 UND1_24 ( .A(A[24]), .B(n1), .Y(Y1[24]) );
  NAND_GATE_1253 UND2_24 ( .A(B[24]), .B(n4), .Y(Y2[24]) );
  NAND_GATE_1252 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  NAND_GATE_1251 UND1_25 ( .A(A[25]), .B(n1), .Y(Y1[25]) );
  NAND_GATE_1250 UND2_25 ( .A(B[25]), .B(n4), .Y(Y2[25]) );
  NAND_GATE_1249 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  NAND_GATE_1248 UND1_26 ( .A(A[26]), .B(n1), .Y(Y1[26]) );
  NAND_GATE_1247 UND2_26 ( .A(B[26]), .B(n4), .Y(Y2[26]) );
  NAND_GATE_1246 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  NAND_GATE_1245 UND1_27 ( .A(A[27]), .B(n1), .Y(Y1[27]) );
  NAND_GATE_1244 UND2_27 ( .A(B[27]), .B(n4), .Y(Y2[27]) );
  NAND_GATE_1243 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  NAND_GATE_1242 UND1_28 ( .A(A[28]), .B(n1), .Y(Y1[28]) );
  NAND_GATE_1241 UND2_28 ( .A(B[28]), .B(n4), .Y(Y2[28]) );
  NAND_GATE_1240 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  NAND_GATE_1239 UND1_29 ( .A(A[29]), .B(n1), .Y(Y1[29]) );
  NAND_GATE_1238 UND2_29 ( .A(B[29]), .B(n4), .Y(Y2[29]) );
  NAND_GATE_1237 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  NAND_GATE_1236 UND1_30 ( .A(A[30]), .B(n1), .Y(Y1[30]) );
  NAND_GATE_1235 UND2_30 ( .A(B[30]), .B(n4), .Y(Y2[30]) );
  NAND_GATE_1234 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  NAND_GATE_1233 UND1_31 ( .A(A[31]), .B(n1), .Y(Y1[31]) );
  NAND_GATE_1232 UND2_31 ( .A(B[31]), .B(n4), .Y(Y2[31]) );
  NAND_GATE_1231 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  BUF_X1 U1 ( .A(SB), .Z(n5) );
  BUF_X1 U2 ( .A(SB), .Z(n4) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GEN_N32_4 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  INV_1_124 UIV ( .A(n1), .Y(SB) );
  NAND_GATE_1230 UND1_0 ( .A(A[0]), .B(n3), .Y(Y1[0]) );
  NAND_GATE_1229 UND2_0 ( .A(B[0]), .B(n6), .Y(Y2[0]) );
  NAND_GATE_1228 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_1227 UND1_1 ( .A(A[1]), .B(n3), .Y(Y1[1]) );
  NAND_GATE_1226 UND2_1 ( .A(B[1]), .B(n6), .Y(Y2[1]) );
  NAND_GATE_1225 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_1224 UND1_2 ( .A(A[2]), .B(n3), .Y(Y1[2]) );
  NAND_GATE_1223 UND2_2 ( .A(B[2]), .B(n6), .Y(Y2[2]) );
  NAND_GATE_1222 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_1221 UND1_3 ( .A(A[3]), .B(n3), .Y(Y1[3]) );
  NAND_GATE_1220 UND2_3 ( .A(B[3]), .B(n6), .Y(Y2[3]) );
  NAND_GATE_1219 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_1218 UND1_4 ( .A(A[4]), .B(n3), .Y(Y1[4]) );
  NAND_GATE_1217 UND2_4 ( .A(B[4]), .B(n6), .Y(Y2[4]) );
  NAND_GATE_1216 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_1215 UND1_5 ( .A(A[5]), .B(n3), .Y(Y1[5]) );
  NAND_GATE_1214 UND2_5 ( .A(B[5]), .B(n6), .Y(Y2[5]) );
  NAND_GATE_1213 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_1212 UND1_6 ( .A(A[6]), .B(n3), .Y(Y1[6]) );
  NAND_GATE_1211 UND2_6 ( .A(B[6]), .B(n5), .Y(Y2[6]) );
  NAND_GATE_1210 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_1209 UND1_7 ( .A(A[7]), .B(n2), .Y(Y1[7]) );
  NAND_GATE_1208 UND2_7 ( .A(B[7]), .B(n5), .Y(Y2[7]) );
  NAND_GATE_1207 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  NAND_GATE_1206 UND1_8 ( .A(A[8]), .B(n2), .Y(Y1[8]) );
  NAND_GATE_1205 UND2_8 ( .A(B[8]), .B(n5), .Y(Y2[8]) );
  NAND_GATE_1204 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  NAND_GATE_1203 UND1_9 ( .A(A[9]), .B(n2), .Y(Y1[9]) );
  NAND_GATE_1202 UND2_9 ( .A(B[9]), .B(n5), .Y(Y2[9]) );
  NAND_GATE_1201 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  NAND_GATE_1200 UND1_10 ( .A(A[10]), .B(n2), .Y(Y1[10]) );
  NAND_GATE_1199 UND2_10 ( .A(B[10]), .B(n5), .Y(Y2[10]) );
  NAND_GATE_1198 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  NAND_GATE_1197 UND1_11 ( .A(A[11]), .B(n2), .Y(Y1[11]) );
  NAND_GATE_1196 UND2_11 ( .A(B[11]), .B(n5), .Y(Y2[11]) );
  NAND_GATE_1195 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  NAND_GATE_1194 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  NAND_GATE_1193 UND2_12 ( .A(B[12]), .B(n5), .Y(Y2[12]) );
  NAND_GATE_1192 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  NAND_GATE_1191 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  NAND_GATE_1190 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  NAND_GATE_1189 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  NAND_GATE_1188 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  NAND_GATE_1187 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  NAND_GATE_1186 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  NAND_GATE_1185 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  NAND_GATE_1184 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  NAND_GATE_1183 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  NAND_GATE_1182 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  NAND_GATE_1181 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  NAND_GATE_1180 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  NAND_GATE_1179 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  NAND_GATE_1178 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  NAND_GATE_1177 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  NAND_GATE_1176 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  NAND_GATE_1175 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  NAND_GATE_1174 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  NAND_GATE_1173 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  NAND_GATE_1172 UND2_19 ( .A(B[19]), .B(n4), .Y(Y2[19]) );
  NAND_GATE_1171 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  NAND_GATE_1170 UND1_20 ( .A(A[20]), .B(n1), .Y(Y1[20]) );
  NAND_GATE_1169 UND2_20 ( .A(B[20]), .B(n4), .Y(Y2[20]) );
  NAND_GATE_1168 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  NAND_GATE_1167 UND1_21 ( .A(A[21]), .B(n1), .Y(Y1[21]) );
  NAND_GATE_1166 UND2_21 ( .A(B[21]), .B(n4), .Y(Y2[21]) );
  NAND_GATE_1165 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  NAND_GATE_1164 UND1_22 ( .A(A[22]), .B(n1), .Y(Y1[22]) );
  NAND_GATE_1163 UND2_22 ( .A(B[22]), .B(n4), .Y(Y2[22]) );
  NAND_GATE_1162 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  NAND_GATE_1161 UND1_23 ( .A(A[23]), .B(n1), .Y(Y1[23]) );
  NAND_GATE_1160 UND2_23 ( .A(B[23]), .B(n4), .Y(Y2[23]) );
  NAND_GATE_1159 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  NAND_GATE_1158 UND1_24 ( .A(A[24]), .B(n1), .Y(Y1[24]) );
  NAND_GATE_1157 UND2_24 ( .A(B[24]), .B(n4), .Y(Y2[24]) );
  NAND_GATE_1156 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  NAND_GATE_1155 UND1_25 ( .A(A[25]), .B(n1), .Y(Y1[25]) );
  NAND_GATE_1154 UND2_25 ( .A(B[25]), .B(n4), .Y(Y2[25]) );
  NAND_GATE_1153 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  NAND_GATE_1152 UND1_26 ( .A(A[26]), .B(n1), .Y(Y1[26]) );
  NAND_GATE_1151 UND2_26 ( .A(B[26]), .B(n4), .Y(Y2[26]) );
  NAND_GATE_1150 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  NAND_GATE_1149 UND1_27 ( .A(A[27]), .B(n1), .Y(Y1[27]) );
  NAND_GATE_1148 UND2_27 ( .A(B[27]), .B(n4), .Y(Y2[27]) );
  NAND_GATE_1147 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  NAND_GATE_1146 UND1_28 ( .A(A[28]), .B(n1), .Y(Y1[28]) );
  NAND_GATE_1145 UND2_28 ( .A(B[28]), .B(n4), .Y(Y2[28]) );
  NAND_GATE_1144 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  NAND_GATE_1143 UND1_29 ( .A(A[29]), .B(n1), .Y(Y1[29]) );
  NAND_GATE_1142 UND2_29 ( .A(B[29]), .B(n4), .Y(Y2[29]) );
  NAND_GATE_1141 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  NAND_GATE_1140 UND1_30 ( .A(A[30]), .B(n1), .Y(Y1[30]) );
  NAND_GATE_1139 UND2_30 ( .A(B[30]), .B(n4), .Y(Y2[30]) );
  NAND_GATE_1138 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  NAND_GATE_1137 UND1_31 ( .A(A[31]), .B(n1), .Y(Y1[31]) );
  NAND_GATE_1136 UND2_31 ( .A(B[31]), .B(n4), .Y(Y2[31]) );
  NAND_GATE_1135 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  BUF_X1 U1 ( .A(SB), .Z(n5) );
  BUF_X1 U2 ( .A(SB), .Z(n4) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GEN_N32_3 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  INV_1_121 UIV ( .A(n1), .Y(SB) );
  NAND_GATE_1119 UND1_0 ( .A(A[0]), .B(n3), .Y(Y1[0]) );
  NAND_GATE_1118 UND2_0 ( .A(B[0]), .B(n6), .Y(Y2[0]) );
  NAND_GATE_1117 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_1116 UND1_1 ( .A(A[1]), .B(n3), .Y(Y1[1]) );
  NAND_GATE_1115 UND2_1 ( .A(B[1]), .B(n6), .Y(Y2[1]) );
  NAND_GATE_1114 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_1113 UND1_2 ( .A(A[2]), .B(n3), .Y(Y1[2]) );
  NAND_GATE_1112 UND2_2 ( .A(B[2]), .B(n6), .Y(Y2[2]) );
  NAND_GATE_1111 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_1110 UND1_3 ( .A(A[3]), .B(n3), .Y(Y1[3]) );
  NAND_GATE_1109 UND2_3 ( .A(B[3]), .B(n6), .Y(Y2[3]) );
  NAND_GATE_1108 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_1107 UND1_4 ( .A(A[4]), .B(n3), .Y(Y1[4]) );
  NAND_GATE_1106 UND2_4 ( .A(B[4]), .B(n6), .Y(Y2[4]) );
  NAND_GATE_1105 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_1104 UND1_5 ( .A(A[5]), .B(n3), .Y(Y1[5]) );
  NAND_GATE_1103 UND2_5 ( .A(B[5]), .B(n6), .Y(Y2[5]) );
  NAND_GATE_1102 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_1101 UND1_6 ( .A(A[6]), .B(n3), .Y(Y1[6]) );
  NAND_GATE_1100 UND2_6 ( .A(B[6]), .B(n5), .Y(Y2[6]) );
  NAND_GATE_1099 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_1098 UND1_7 ( .A(A[7]), .B(n2), .Y(Y1[7]) );
  NAND_GATE_1097 UND2_7 ( .A(B[7]), .B(n5), .Y(Y2[7]) );
  NAND_GATE_1096 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  NAND_GATE_1095 UND1_8 ( .A(A[8]), .B(n2), .Y(Y1[8]) );
  NAND_GATE_1094 UND2_8 ( .A(B[8]), .B(n5), .Y(Y2[8]) );
  NAND_GATE_1093 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  NAND_GATE_1092 UND1_9 ( .A(A[9]), .B(n2), .Y(Y1[9]) );
  NAND_GATE_1091 UND2_9 ( .A(B[9]), .B(n5), .Y(Y2[9]) );
  NAND_GATE_1090 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  NAND_GATE_1089 UND1_10 ( .A(A[10]), .B(n2), .Y(Y1[10]) );
  NAND_GATE_1088 UND2_10 ( .A(B[10]), .B(n5), .Y(Y2[10]) );
  NAND_GATE_1087 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  NAND_GATE_1086 UND1_11 ( .A(A[11]), .B(n2), .Y(Y1[11]) );
  NAND_GATE_1085 UND2_11 ( .A(B[11]), .B(n5), .Y(Y2[11]) );
  NAND_GATE_1084 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  NAND_GATE_1083 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  NAND_GATE_1082 UND2_12 ( .A(B[12]), .B(n5), .Y(Y2[12]) );
  NAND_GATE_1081 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  NAND_GATE_1080 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  NAND_GATE_1079 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  NAND_GATE_1078 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  NAND_GATE_1077 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  NAND_GATE_1076 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  NAND_GATE_1075 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  NAND_GATE_1074 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  NAND_GATE_1073 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  NAND_GATE_1072 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  NAND_GATE_1071 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  NAND_GATE_1070 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  NAND_GATE_1069 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  NAND_GATE_1068 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  NAND_GATE_1067 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  NAND_GATE_1066 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  NAND_GATE_1065 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  NAND_GATE_1064 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  NAND_GATE_1063 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  NAND_GATE_1062 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  NAND_GATE_1061 UND2_19 ( .A(B[19]), .B(n4), .Y(Y2[19]) );
  NAND_GATE_1060 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  NAND_GATE_1059 UND1_20 ( .A(A[20]), .B(n1), .Y(Y1[20]) );
  NAND_GATE_1058 UND2_20 ( .A(B[20]), .B(n4), .Y(Y2[20]) );
  NAND_GATE_1057 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  NAND_GATE_1056 UND1_21 ( .A(A[21]), .B(n1), .Y(Y1[21]) );
  NAND_GATE_1055 UND2_21 ( .A(B[21]), .B(n4), .Y(Y2[21]) );
  NAND_GATE_1054 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  NAND_GATE_1053 UND1_22 ( .A(A[22]), .B(n1), .Y(Y1[22]) );
  NAND_GATE_1052 UND2_22 ( .A(B[22]), .B(n4), .Y(Y2[22]) );
  NAND_GATE_1051 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  NAND_GATE_1050 UND1_23 ( .A(A[23]), .B(n1), .Y(Y1[23]) );
  NAND_GATE_1049 UND2_23 ( .A(B[23]), .B(n4), .Y(Y2[23]) );
  NAND_GATE_1048 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  NAND_GATE_1047 UND1_24 ( .A(A[24]), .B(n1), .Y(Y1[24]) );
  NAND_GATE_1046 UND2_24 ( .A(B[24]), .B(n4), .Y(Y2[24]) );
  NAND_GATE_1045 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  NAND_GATE_1044 UND1_25 ( .A(A[25]), .B(n1), .Y(Y1[25]) );
  NAND_GATE_1043 UND2_25 ( .A(B[25]), .B(n4), .Y(Y2[25]) );
  NAND_GATE_1042 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  NAND_GATE_1041 UND1_26 ( .A(A[26]), .B(n1), .Y(Y1[26]) );
  NAND_GATE_1040 UND2_26 ( .A(B[26]), .B(n4), .Y(Y2[26]) );
  NAND_GATE_1039 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  NAND_GATE_1038 UND1_27 ( .A(A[27]), .B(n1), .Y(Y1[27]) );
  NAND_GATE_1037 UND2_27 ( .A(B[27]), .B(n4), .Y(Y2[27]) );
  NAND_GATE_1036 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  NAND_GATE_1035 UND1_28 ( .A(A[28]), .B(n1), .Y(Y1[28]) );
  NAND_GATE_1034 UND2_28 ( .A(B[28]), .B(n4), .Y(Y2[28]) );
  NAND_GATE_1033 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  NAND_GATE_1032 UND1_29 ( .A(A[29]), .B(n1), .Y(Y1[29]) );
  NAND_GATE_1031 UND2_29 ( .A(B[29]), .B(n4), .Y(Y2[29]) );
  NAND_GATE_1030 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  NAND_GATE_1029 UND1_30 ( .A(A[30]), .B(n1), .Y(Y1[30]) );
  NAND_GATE_1028 UND2_30 ( .A(B[30]), .B(n4), .Y(Y2[30]) );
  NAND_GATE_1027 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  NAND_GATE_1026 UND1_31 ( .A(A[31]), .B(n1), .Y(Y1[31]) );
  NAND_GATE_1025 UND2_31 ( .A(B[31]), .B(n4), .Y(Y2[31]) );
  NAND_GATE_1024 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  BUF_X1 U1 ( .A(SB), .Z(n5) );
  BUF_X1 U2 ( .A(SB), .Z(n4) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  BUF_X1 U5 ( .A(SEL), .Z(n2) );
  BUF_X1 U6 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_GEN_N32_2 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  INV_1_39 UIV ( .A(n1), .Y(SB) );
  NAND_GATE_918 UND1_0 ( .A(A[0]), .B(n3), .Y(Y1[0]) );
  NAND_GATE_917 UND2_0 ( .A(B[0]), .B(n6), .Y(Y2[0]) );
  NAND_GATE_916 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_915 UND1_1 ( .A(A[1]), .B(n3), .Y(Y1[1]) );
  NAND_GATE_914 UND2_1 ( .A(B[1]), .B(n6), .Y(Y2[1]) );
  NAND_GATE_913 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_912 UND1_2 ( .A(A[2]), .B(n3), .Y(Y1[2]) );
  NAND_GATE_911 UND2_2 ( .A(B[2]), .B(n6), .Y(Y2[2]) );
  NAND_GATE_910 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_909 UND1_3 ( .A(A[3]), .B(n3), .Y(Y1[3]) );
  NAND_GATE_908 UND2_3 ( .A(B[3]), .B(n6), .Y(Y2[3]) );
  NAND_GATE_907 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_906 UND1_4 ( .A(A[4]), .B(n3), .Y(Y1[4]) );
  NAND_GATE_905 UND2_4 ( .A(B[4]), .B(n6), .Y(Y2[4]) );
  NAND_GATE_904 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_903 UND1_5 ( .A(A[5]), .B(n3), .Y(Y1[5]) );
  NAND_GATE_902 UND2_5 ( .A(B[5]), .B(n6), .Y(Y2[5]) );
  NAND_GATE_901 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_900 UND1_6 ( .A(A[6]), .B(n3), .Y(Y1[6]) );
  NAND_GATE_899 UND2_6 ( .A(B[6]), .B(n5), .Y(Y2[6]) );
  NAND_GATE_898 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_897 UND1_7 ( .A(A[7]), .B(n2), .Y(Y1[7]) );
  NAND_GATE_896 UND2_7 ( .A(B[7]), .B(n5), .Y(Y2[7]) );
  NAND_GATE_895 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  NAND_GATE_894 UND1_8 ( .A(A[8]), .B(n2), .Y(Y1[8]) );
  NAND_GATE_893 UND2_8 ( .A(B[8]), .B(n5), .Y(Y2[8]) );
  NAND_GATE_892 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  NAND_GATE_891 UND1_9 ( .A(A[9]), .B(n2), .Y(Y1[9]) );
  NAND_GATE_890 UND2_9 ( .A(B[9]), .B(n5), .Y(Y2[9]) );
  NAND_GATE_889 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  NAND_GATE_888 UND1_10 ( .A(A[10]), .B(n2), .Y(Y1[10]) );
  NAND_GATE_887 UND2_10 ( .A(B[10]), .B(n5), .Y(Y2[10]) );
  NAND_GATE_886 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  NAND_GATE_885 UND1_11 ( .A(A[11]), .B(n2), .Y(Y1[11]) );
  NAND_GATE_884 UND2_11 ( .A(B[11]), .B(n5), .Y(Y2[11]) );
  NAND_GATE_883 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  NAND_GATE_882 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  NAND_GATE_881 UND2_12 ( .A(B[12]), .B(n5), .Y(Y2[12]) );
  NAND_GATE_880 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  NAND_GATE_879 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  NAND_GATE_878 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  NAND_GATE_877 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  NAND_GATE_876 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  NAND_GATE_875 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  NAND_GATE_874 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  NAND_GATE_873 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  NAND_GATE_872 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  NAND_GATE_871 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  NAND_GATE_870 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  NAND_GATE_869 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  NAND_GATE_868 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  NAND_GATE_867 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  NAND_GATE_866 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  NAND_GATE_865 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  NAND_GATE_864 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  NAND_GATE_863 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  NAND_GATE_862 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  NAND_GATE_861 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  NAND_GATE_860 UND2_19 ( .A(B[19]), .B(n4), .Y(Y2[19]) );
  NAND_GATE_859 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  NAND_GATE_858 UND1_20 ( .A(A[20]), .B(n1), .Y(Y1[20]) );
  NAND_GATE_857 UND2_20 ( .A(B[20]), .B(n4), .Y(Y2[20]) );
  NAND_GATE_856 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  NAND_GATE_855 UND1_21 ( .A(A[21]), .B(n1), .Y(Y1[21]) );
  NAND_GATE_854 UND2_21 ( .A(B[21]), .B(n4), .Y(Y2[21]) );
  NAND_GATE_853 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  NAND_GATE_852 UND1_22 ( .A(A[22]), .B(n1), .Y(Y1[22]) );
  NAND_GATE_851 UND2_22 ( .A(B[22]), .B(n4), .Y(Y2[22]) );
  NAND_GATE_850 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  NAND_GATE_849 UND1_23 ( .A(A[23]), .B(n1), .Y(Y1[23]) );
  NAND_GATE_848 UND2_23 ( .A(B[23]), .B(n4), .Y(Y2[23]) );
  NAND_GATE_847 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  NAND_GATE_846 UND1_24 ( .A(A[24]), .B(n1), .Y(Y1[24]) );
  NAND_GATE_845 UND2_24 ( .A(B[24]), .B(n4), .Y(Y2[24]) );
  NAND_GATE_844 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  NAND_GATE_843 UND1_25 ( .A(A[25]), .B(n1), .Y(Y1[25]) );
  NAND_GATE_842 UND2_25 ( .A(B[25]), .B(n4), .Y(Y2[25]) );
  NAND_GATE_841 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  NAND_GATE_840 UND1_26 ( .A(A[26]), .B(n1), .Y(Y1[26]) );
  NAND_GATE_839 UND2_26 ( .A(B[26]), .B(n4), .Y(Y2[26]) );
  NAND_GATE_838 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  NAND_GATE_837 UND1_27 ( .A(A[27]), .B(n1), .Y(Y1[27]) );
  NAND_GATE_836 UND2_27 ( .A(B[27]), .B(n4), .Y(Y2[27]) );
  NAND_GATE_835 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  NAND_GATE_834 UND1_28 ( .A(A[28]), .B(n1), .Y(Y1[28]) );
  NAND_GATE_833 UND2_28 ( .A(B[28]), .B(n4), .Y(Y2[28]) );
  NAND_GATE_832 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  NAND_GATE_831 UND1_29 ( .A(A[29]), .B(n1), .Y(Y1[29]) );
  NAND_GATE_830 UND2_29 ( .A(B[29]), .B(n4), .Y(Y2[29]) );
  NAND_GATE_829 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  NAND_GATE_828 UND1_30 ( .A(A[30]), .B(n1), .Y(Y1[30]) );
  NAND_GATE_827 UND2_30 ( .A(B[30]), .B(n4), .Y(Y2[30]) );
  NAND_GATE_826 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  NAND_GATE_825 UND1_31 ( .A(A[31]), .B(n1), .Y(Y1[31]) );
  NAND_GATE_824 UND2_31 ( .A(B[31]), .B(n4), .Y(Y2[31]) );
  NAND_GATE_823 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  BUF_X1 U1 ( .A(SB), .Z(n5) );
  BUF_X1 U2 ( .A(SB), .Z(n4) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n3) );
  BUF_X1 U5 ( .A(SEL), .Z(n1) );
  BUF_X1 U6 ( .A(SEL), .Z(n2) );
endmodule


module MUX21_GEN_N32_1 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  INV_1_38 UIV ( .A(n1), .Y(SB) );
  NAND_GATE_822 UND1_0 ( .A(A[0]), .B(n3), .Y(Y1[0]) );
  NAND_GATE_821 UND2_0 ( .A(B[0]), .B(n6), .Y(Y2[0]) );
  NAND_GATE_820 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_819 UND1_1 ( .A(A[1]), .B(n3), .Y(Y1[1]) );
  NAND_GATE_818 UND2_1 ( .A(B[1]), .B(n6), .Y(Y2[1]) );
  NAND_GATE_817 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_816 UND1_2 ( .A(A[2]), .B(n3), .Y(Y1[2]) );
  NAND_GATE_815 UND2_2 ( .A(B[2]), .B(n6), .Y(Y2[2]) );
  NAND_GATE_814 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_813 UND1_3 ( .A(A[3]), .B(n3), .Y(Y1[3]) );
  NAND_GATE_812 UND2_3 ( .A(B[3]), .B(n6), .Y(Y2[3]) );
  NAND_GATE_811 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_810 UND1_4 ( .A(A[4]), .B(n3), .Y(Y1[4]) );
  NAND_GATE_809 UND2_4 ( .A(B[4]), .B(n6), .Y(Y2[4]) );
  NAND_GATE_808 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_807 UND1_5 ( .A(A[5]), .B(n3), .Y(Y1[5]) );
  NAND_GATE_806 UND2_5 ( .A(B[5]), .B(n6), .Y(Y2[5]) );
  NAND_GATE_805 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_804 UND1_6 ( .A(A[6]), .B(n3), .Y(Y1[6]) );
  NAND_GATE_803 UND2_6 ( .A(B[6]), .B(n5), .Y(Y2[6]) );
  NAND_GATE_802 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_801 UND1_7 ( .A(A[7]), .B(n2), .Y(Y1[7]) );
  NAND_GATE_800 UND2_7 ( .A(B[7]), .B(n5), .Y(Y2[7]) );
  NAND_GATE_799 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  NAND_GATE_798 UND1_8 ( .A(A[8]), .B(n2), .Y(Y1[8]) );
  NAND_GATE_797 UND2_8 ( .A(B[8]), .B(n5), .Y(Y2[8]) );
  NAND_GATE_796 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  NAND_GATE_795 UND1_9 ( .A(A[9]), .B(n2), .Y(Y1[9]) );
  NAND_GATE_794 UND2_9 ( .A(B[9]), .B(n5), .Y(Y2[9]) );
  NAND_GATE_793 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  NAND_GATE_792 UND1_10 ( .A(A[10]), .B(n2), .Y(Y1[10]) );
  NAND_GATE_791 UND2_10 ( .A(B[10]), .B(n5), .Y(Y2[10]) );
  NAND_GATE_790 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  NAND_GATE_789 UND1_11 ( .A(A[11]), .B(n2), .Y(Y1[11]) );
  NAND_GATE_788 UND2_11 ( .A(B[11]), .B(n5), .Y(Y2[11]) );
  NAND_GATE_787 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  NAND_GATE_786 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  NAND_GATE_785 UND2_12 ( .A(B[12]), .B(n5), .Y(Y2[12]) );
  NAND_GATE_784 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  NAND_GATE_783 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  NAND_GATE_782 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  NAND_GATE_781 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  NAND_GATE_780 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  NAND_GATE_779 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  NAND_GATE_778 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  NAND_GATE_777 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  NAND_GATE_776 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  NAND_GATE_775 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  NAND_GATE_774 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  NAND_GATE_773 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  NAND_GATE_772 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  NAND_GATE_771 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  NAND_GATE_770 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  NAND_GATE_769 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  NAND_GATE_768 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  NAND_GATE_767 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  NAND_GATE_766 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  NAND_GATE_765 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  NAND_GATE_764 UND2_19 ( .A(B[19]), .B(n4), .Y(Y2[19]) );
  NAND_GATE_763 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  NAND_GATE_762 UND1_20 ( .A(A[20]), .B(n1), .Y(Y1[20]) );
  NAND_GATE_761 UND2_20 ( .A(B[20]), .B(n4), .Y(Y2[20]) );
  NAND_GATE_760 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  NAND_GATE_759 UND1_21 ( .A(A[21]), .B(n1), .Y(Y1[21]) );
  NAND_GATE_758 UND2_21 ( .A(B[21]), .B(n4), .Y(Y2[21]) );
  NAND_GATE_757 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  NAND_GATE_756 UND1_22 ( .A(A[22]), .B(n1), .Y(Y1[22]) );
  NAND_GATE_755 UND2_22 ( .A(B[22]), .B(n4), .Y(Y2[22]) );
  NAND_GATE_754 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  NAND_GATE_753 UND1_23 ( .A(A[23]), .B(n1), .Y(Y1[23]) );
  NAND_GATE_752 UND2_23 ( .A(B[23]), .B(n4), .Y(Y2[23]) );
  NAND_GATE_751 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  NAND_GATE_750 UND1_24 ( .A(A[24]), .B(n1), .Y(Y1[24]) );
  NAND_GATE_749 UND2_24 ( .A(B[24]), .B(n4), .Y(Y2[24]) );
  NAND_GATE_748 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  NAND_GATE_747 UND1_25 ( .A(A[25]), .B(n1), .Y(Y1[25]) );
  NAND_GATE_746 UND2_25 ( .A(B[25]), .B(n4), .Y(Y2[25]) );
  NAND_GATE_745 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  NAND_GATE_744 UND1_26 ( .A(A[26]), .B(n1), .Y(Y1[26]) );
  NAND_GATE_743 UND2_26 ( .A(B[26]), .B(n4), .Y(Y2[26]) );
  NAND_GATE_742 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  NAND_GATE_741 UND1_27 ( .A(A[27]), .B(n1), .Y(Y1[27]) );
  NAND_GATE_740 UND2_27 ( .A(B[27]), .B(n4), .Y(Y2[27]) );
  NAND_GATE_739 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  NAND_GATE_738 UND1_28 ( .A(A[28]), .B(n1), .Y(Y1[28]) );
  NAND_GATE_737 UND2_28 ( .A(B[28]), .B(n4), .Y(Y2[28]) );
  NAND_GATE_736 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  NAND_GATE_735 UND1_29 ( .A(A[29]), .B(n1), .Y(Y1[29]) );
  NAND_GATE_734 UND2_29 ( .A(B[29]), .B(n4), .Y(Y2[29]) );
  NAND_GATE_733 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  NAND_GATE_732 UND1_30 ( .A(A[30]), .B(n1), .Y(Y1[30]) );
  NAND_GATE_731 UND2_30 ( .A(B[30]), .B(n4), .Y(Y2[30]) );
  NAND_GATE_730 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  NAND_GATE_729 UND1_31 ( .A(A[31]), .B(n1), .Y(Y1[31]) );
  NAND_GATE_728 UND2_31 ( .A(B[31]), .B(n4), .Y(Y2[31]) );
  NAND_GATE_727 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  BUF_X1 U1 ( .A(SB), .Z(n5) );
  BUF_X1 U2 ( .A(SB), .Z(n4) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n3) );
  BUF_X1 U5 ( .A(SEL), .Z(n1) );
  BUF_X1 U6 ( .A(SEL), .Z(n2) );
endmodule


module REG_N5_2 ( D, Q, EN, RST, CLK );
  input [4:0] D;
  output [4:0] Q;
  input EN, RST, CLK;


  FD_1_383 FF_0 ( .D(D[0]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[0]) );
  FD_1_382 FF_1 ( .D(D[1]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[1]) );
  FD_1_381 FF_2 ( .D(D[2]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[2]) );
  FD_1_380 FF_3 ( .D(D[3]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[3]) );
  FD_1_379 FF_4 ( .D(D[4]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[4]) );
endmodule


module REG_N5_1 ( D, Q, EN, RST, CLK );
  input [4:0] D;
  output [4:0] Q;
  input EN, RST, CLK;


  FD_1_282 FF_0 ( .D(D[0]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[0]) );
  FD_1_281 FF_1 ( .D(D[1]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[1]) );
  FD_1_280 FF_2 ( .D(D[2]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[2]) );
  FD_1_279 FF_3 ( .D(D[3]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[3]) );
  FD_1_278 FF_4 ( .D(D[4]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[4]) );
endmodule


module XOR_GATE_1 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module AND_GATE_340 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_339 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_338 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_337 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_336 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_335 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_334 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_333 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_332 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_331 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_330 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_329 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_328 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_327 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_326 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_325 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_324 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_323 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_322 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_321 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_320 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_319 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_318 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_317 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_316 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_315 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_314 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_313 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_312 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_311 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_310 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_309 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_308 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_307 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_306 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_305 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_304 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_303 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_302 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_301 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_300 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_299 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_298 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_297 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_296 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_295 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_294 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_293 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_292 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_291 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_290 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_289 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_288 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_287 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_286 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_285 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_284 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_283 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_282 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_281 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_280 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_279 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_278 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_277 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_276 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_275 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_274 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_273 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_272 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_271 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_270 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_269 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_268 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_267 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_266 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_265 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_264 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_263 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_262 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_261 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_260 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_259 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_258 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_257 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_256 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_255 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_254 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_253 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_252 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_251 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_250 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_249 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_248 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_247 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_246 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_245 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_244 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_243 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_242 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_241 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_240 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_239 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_238 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_237 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_236 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_235 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_234 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_233 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_232 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_231 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_230 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_229 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_228 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_227 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_226 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_225 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_224 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_223 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_222 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_221 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_220 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_219 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_218 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_217 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_216 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_215 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_214 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_213 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_212 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_211 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_210 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_209 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_208 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_207 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_206 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_205 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_204 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_203 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_202 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_201 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_200 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_199 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_198 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_197 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_196 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_195 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_194 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_193 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_192 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_191 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_190 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_189 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_188 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_187 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_186 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_185 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_184 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_183 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_182 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_181 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_180 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_179 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_178 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_177 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_176 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_175 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_174 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_173 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_172 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_171 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_170 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_169 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_168 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_167 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_166 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_165 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_164 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_163 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_162 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_161 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_160 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_159 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_158 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_157 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_156 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_155 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_154 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_153 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_152 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_151 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_150 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_149 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_148 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_147 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_146 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_145 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_144 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_143 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_142 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_141 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_140 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_139 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_138 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_137 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_136 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_135 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_134 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_133 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_132 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_131 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_130 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_129 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_128 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_127 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_126 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_125 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_124 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_123 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_122 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_121 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_120 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_119 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_118 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_117 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_116 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_115 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_114 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_113 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_112 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_111 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_110 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_109 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_108 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_107 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_106 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_105 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_104 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_103 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_102 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_101 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_100 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_99 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_98 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_97 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_96 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_95 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_94 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_93 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_92 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_91 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_90 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_89 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_88 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_87 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_86 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_85 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_84 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_83 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_82 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_81 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_80 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_79 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_78 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_77 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_76 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_75 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_74 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_73 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_72 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_71 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_70 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_69 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_68 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_67 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_66 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_65 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_64 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_63 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_62 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_61 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_60 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_59 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_58 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_57 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_56 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_55 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_54 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_53 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_52 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_51 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_50 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_49 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_48 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_47 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_46 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_45 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_44 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_43 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_42 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_41 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_40 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_39 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_38 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_37 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_36 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_35 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_34 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_33 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_32 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_31 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_30 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_29 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_28 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_27 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_26 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_25 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_24 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_23 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_22 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_21 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_20 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_19 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_18 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_17 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_16 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_15 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_14 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_13 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_12 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_11 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_10 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_9 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_8 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_7 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_6 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_5 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_4 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_3 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_2 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module AND_GATE_1 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module INV_169 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_168 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_167 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_166 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_165 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_164 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_163 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_162 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_161 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_160 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_159 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_158 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_157 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_156 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_155 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_154 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_153 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_152 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_151 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_150 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_149 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_148 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_147 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_146 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_145 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_144 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_143 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_142 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_141 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_140 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_139 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_138 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_137 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_136 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_135 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_134 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_133 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_132 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_131 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_130 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_129 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_128 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_127 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_126 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_125 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_124 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_123 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_122 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_121 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_120 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_119 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_118 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_117 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_116 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_115 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_114 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_113 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_112 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_111 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_110 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_109 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_108 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_107 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_106 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_105 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_104 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_103 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_102 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_101 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_100 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_99 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_98 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_97 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_96 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_95 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_94 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_93 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_92 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_91 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_90 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_89 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_88 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_87 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_86 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_85 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_84 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_83 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_82 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_81 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_80 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_79 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_78 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_77 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_76 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_75 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_74 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_73 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_72 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_71 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_70 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_69 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_68 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_67 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_66 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_65 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_64 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_63 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_62 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_61 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_60 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_59 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_58 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_57 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_56 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_55 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_54 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_53 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_52 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_51 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_50 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_49 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_48 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_47 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_46 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_45 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_44 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_43 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_42 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_41 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_40 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_39 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_38 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_37 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_36 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_35 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_34 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_33 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_32 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_31 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_30 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_29 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_28 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_27 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_26 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_25 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_24 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_23 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_22 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_21 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_20 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_19 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_18 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_17 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_16 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_15 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_14 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_13 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_12 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_11 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_10 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_9 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_8 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_7 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_6 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_5 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_4 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_3 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_2 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module INV_1 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module REG_N32_14 ( D, Q, EN, RST, CLK );
  input [31:0] D;
  output [31:0] Q;
  input EN, RST, CLK;
  wire   n1, n2, n3, n4, n5, n6;

  FD_1_548 FF_0 ( .D(D[0]), .CLK(CLK), .EN(n4), .RST(n1), .Q(Q[0]) );
  FD_1_547 FF_1 ( .D(D[1]), .CLK(CLK), .EN(n4), .RST(n1), .Q(Q[1]) );
  FD_1_546 FF_2 ( .D(D[2]), .CLK(CLK), .EN(n4), .RST(n1), .Q(Q[2]) );
  FD_1_545 FF_3 ( .D(D[3]), .CLK(CLK), .EN(n4), .RST(n1), .Q(Q[3]) );
  FD_1_544 FF_4 ( .D(D[4]), .CLK(CLK), .EN(n4), .RST(n1), .Q(Q[4]) );
  FD_1_543 FF_5 ( .D(D[5]), .CLK(CLK), .EN(n4), .RST(n1), .Q(Q[5]) );
  FD_1_542 FF_6 ( .D(D[6]), .CLK(CLK), .EN(n4), .RST(n1), .Q(Q[6]) );
  FD_1_541 FF_7 ( .D(D[7]), .CLK(CLK), .EN(n4), .RST(n1), .Q(Q[7]) );
  FD_1_540 FF_8 ( .D(D[8]), .CLK(CLK), .EN(n4), .RST(n1), .Q(Q[8]) );
  FD_1_539 FF_9 ( .D(D[9]), .CLK(CLK), .EN(n4), .RST(n1), .Q(Q[9]) );
  FD_1_538 FF_10 ( .D(D[10]), .CLK(CLK), .EN(n4), .RST(n1), .Q(Q[10]) );
  FD_1_537 FF_11 ( .D(D[11]), .CLK(CLK), .EN(n4), .RST(n1), .Q(Q[11]) );
  FD_1_536 FF_12 ( .D(D[12]), .CLK(CLK), .EN(n4), .RST(n1), .Q(Q[12]) );
  FD_1_535 FF_13 ( .D(D[13]), .CLK(CLK), .EN(n5), .RST(n2), .Q(Q[13]) );
  FD_1_534 FF_14 ( .D(D[14]), .CLK(CLK), .EN(n5), .RST(n2), .Q(Q[14]) );
  FD_1_533 FF_15 ( .D(D[15]), .CLK(CLK), .EN(n5), .RST(n2), .Q(Q[15]) );
  FD_1_532 FF_16 ( .D(D[16]), .CLK(CLK), .EN(n5), .RST(n2), .Q(Q[16]) );
  FD_1_531 FF_17 ( .D(D[17]), .CLK(CLK), .EN(n5), .RST(n2), .Q(Q[17]) );
  FD_1_530 FF_18 ( .D(D[18]), .CLK(CLK), .EN(n5), .RST(n2), .Q(Q[18]) );
  FD_1_529 FF_19 ( .D(D[19]), .CLK(CLK), .EN(n5), .RST(n2), .Q(Q[19]) );
  FD_1_528 FF_20 ( .D(D[20]), .CLK(CLK), .EN(n5), .RST(n2), .Q(Q[20]) );
  FD_1_527 FF_21 ( .D(D[21]), .CLK(CLK), .EN(n5), .RST(n2), .Q(Q[21]) );
  FD_1_526 FF_22 ( .D(D[22]), .CLK(CLK), .EN(n5), .RST(n2), .Q(Q[22]) );
  FD_1_525 FF_23 ( .D(D[23]), .CLK(CLK), .EN(n5), .RST(n2), .Q(Q[23]) );
  FD_1_524 FF_24 ( .D(D[24]), .CLK(CLK), .EN(n5), .RST(n2), .Q(Q[24]) );
  FD_1_523 FF_25 ( .D(D[25]), .CLK(CLK), .EN(n5), .RST(n2), .Q(Q[25]) );
  FD_1_522 FF_26 ( .D(D[26]), .CLK(CLK), .EN(n6), .RST(n3), .Q(Q[26]) );
  FD_1_521 FF_27 ( .D(D[27]), .CLK(CLK), .EN(n6), .RST(n3), .Q(Q[27]) );
  FD_1_520 FF_28 ( .D(D[28]), .CLK(CLK), .EN(n6), .RST(n3), .Q(Q[28]) );
  FD_1_519 FF_29 ( .D(D[29]), .CLK(CLK), .EN(n6), .RST(n3), .Q(Q[29]) );
  FD_1_518 FF_30 ( .D(D[30]), .CLK(CLK), .EN(n6), .RST(n3), .Q(Q[30]) );
  FD_1_517 FF_31 ( .D(D[31]), .CLK(CLK), .EN(n6), .RST(n3), .Q(Q[31]) );
  BUF_X1 U1 ( .A(EN), .Z(n4) );
  BUF_X1 U2 ( .A(EN), .Z(n5) );
  BUF_X1 U3 ( .A(EN), .Z(n6) );
  BUF_X1 U4 ( .A(RST), .Z(n1) );
  BUF_X1 U5 ( .A(RST), .Z(n2) );
  BUF_X1 U6 ( .A(RST), .Z(n3) );
endmodule


module REG_N32_13 ( D, Q, EN, RST, CLK );
  input [31:0] D;
  output [31:0] Q;
  input EN, RST, CLK;
  wire   n1, n2, n3, n4, n5, n6;

  FD_1_516 FF_0 ( .D(D[0]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[0]) );
  FD_1_515 FF_1 ( .D(D[1]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[1]) );
  FD_1_514 FF_2 ( .D(D[2]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[2]) );
  FD_1_513 FF_3 ( .D(D[3]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[3]) );
  FD_1_512 FF_4 ( .D(D[4]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[4]) );
  FD_1_511 FF_5 ( .D(D[5]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[5]) );
  FD_1_510 FF_6 ( .D(D[6]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[6]) );
  FD_1_509 FF_7 ( .D(D[7]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[7]) );
  FD_1_508 FF_8 ( .D(D[8]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[8]) );
  FD_1_507 FF_9 ( .D(D[9]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[9]) );
  FD_1_506 FF_10 ( .D(D[10]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[10]) );
  FD_1_505 FF_11 ( .D(D[11]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[11]) );
  FD_1_504 FF_12 ( .D(D[12]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[12]) );
  FD_1_503 FF_13 ( .D(D[13]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[13]) );
  FD_1_502 FF_14 ( .D(D[14]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[14]) );
  FD_1_501 FF_15 ( .D(D[15]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[15]) );
  FD_1_500 FF_16 ( .D(D[16]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[16]) );
  FD_1_499 FF_17 ( .D(D[17]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[17]) );
  FD_1_498 FF_18 ( .D(D[18]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[18]) );
  FD_1_497 FF_19 ( .D(D[19]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[19]) );
  FD_1_496 FF_20 ( .D(D[20]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[20]) );
  FD_1_495 FF_21 ( .D(D[21]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[21]) );
  FD_1_494 FF_22 ( .D(D[22]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[22]) );
  FD_1_493 FF_23 ( .D(D[23]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[23]) );
  FD_1_492 FF_24 ( .D(D[24]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[24]) );
  FD_1_491 FF_25 ( .D(D[25]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[25]) );
  FD_1_490 FF_26 ( .D(D[26]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[26]) );
  FD_1_489 FF_27 ( .D(D[27]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[27]) );
  FD_1_488 FF_28 ( .D(D[28]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[28]) );
  FD_1_487 FF_29 ( .D(D[29]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[29]) );
  FD_1_486 FF_30 ( .D(D[30]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[30]) );
  FD_1_485 FF_31 ( .D(D[31]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[31]) );
  CLKBUF_X1 U1 ( .A(EN), .Z(n1) );
  CLKBUF_X1 U2 ( .A(EN), .Z(n2) );
  CLKBUF_X1 U3 ( .A(EN), .Z(n3) );
  BUF_X1 U4 ( .A(RST), .Z(n6) );
  BUF_X1 U5 ( .A(RST), .Z(n4) );
  BUF_X1 U6 ( .A(RST), .Z(n5) );
endmodule


module REG_N32_12 ( D, Q, EN, RST, CLK );
  input [31:0] D;
  output [31:0] Q;
  input EN, RST, CLK;
  wire   n1, n2, n3, n4, n5, n6;

  FD_1_484 FF_0 ( .D(D[0]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[0]) );
  FD_1_483 FF_1 ( .D(D[1]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[1]) );
  FD_1_482 FF_2 ( .D(D[2]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[2]) );
  FD_1_481 FF_3 ( .D(D[3]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[3]) );
  FD_1_480 FF_4 ( .D(D[4]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[4]) );
  FD_1_479 FF_5 ( .D(D[5]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[5]) );
  FD_1_478 FF_6 ( .D(D[6]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[6]) );
  FD_1_477 FF_7 ( .D(D[7]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[7]) );
  FD_1_476 FF_8 ( .D(D[8]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[8]) );
  FD_1_475 FF_9 ( .D(D[9]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[9]) );
  FD_1_474 FF_10 ( .D(D[10]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[10]) );
  FD_1_473 FF_11 ( .D(D[11]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[11]) );
  FD_1_472 FF_12 ( .D(D[12]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[12]) );
  FD_1_471 FF_13 ( .D(D[13]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[13]) );
  FD_1_470 FF_14 ( .D(D[14]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[14]) );
  FD_1_469 FF_15 ( .D(D[15]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[15]) );
  FD_1_468 FF_16 ( .D(D[16]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[16]) );
  FD_1_467 FF_17 ( .D(D[17]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[17]) );
  FD_1_466 FF_18 ( .D(D[18]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[18]) );
  FD_1_465 FF_19 ( .D(D[19]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[19]) );
  FD_1_464 FF_20 ( .D(D[20]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[20]) );
  FD_1_463 FF_21 ( .D(D[21]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[21]) );
  FD_1_462 FF_22 ( .D(D[22]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[22]) );
  FD_1_461 FF_23 ( .D(D[23]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[23]) );
  FD_1_460 FF_24 ( .D(D[24]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[24]) );
  FD_1_459 FF_25 ( .D(D[25]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[25]) );
  FD_1_458 FF_26 ( .D(D[26]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[26]) );
  FD_1_457 FF_27 ( .D(D[27]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[27]) );
  FD_1_456 FF_28 ( .D(D[28]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[28]) );
  FD_1_455 FF_29 ( .D(D[29]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[29]) );
  FD_1_454 FF_30 ( .D(D[30]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[30]) );
  FD_1_453 FF_31 ( .D(D[31]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[31]) );
  CLKBUF_X1 U1 ( .A(EN), .Z(n1) );
  CLKBUF_X1 U2 ( .A(EN), .Z(n2) );
  CLKBUF_X1 U3 ( .A(EN), .Z(n3) );
  BUF_X1 U4 ( .A(RST), .Z(n6) );
  BUF_X1 U5 ( .A(RST), .Z(n4) );
  BUF_X1 U6 ( .A(RST), .Z(n5) );
endmodule


module REG_N32_11 ( D, Q, EN, RST, CLK );
  input [31:0] D;
  output [31:0] Q;
  input EN, RST, CLK;
  wire   n1, n2, n3, n4, n5, n6;

  FD_1_452 FF_0 ( .D(D[0]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[0]) );
  FD_1_451 FF_1 ( .D(D[1]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[1]) );
  FD_1_450 FF_2 ( .D(D[2]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[2]) );
  FD_1_449 FF_3 ( .D(D[3]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[3]) );
  FD_1_448 FF_4 ( .D(D[4]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[4]) );
  FD_1_447 FF_5 ( .D(D[5]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[5]) );
  FD_1_446 FF_6 ( .D(D[6]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[6]) );
  FD_1_445 FF_7 ( .D(D[7]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[7]) );
  FD_1_444 FF_8 ( .D(D[8]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[8]) );
  FD_1_443 FF_9 ( .D(D[9]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[9]) );
  FD_1_442 FF_10 ( .D(D[10]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[10]) );
  FD_1_441 FF_11 ( .D(D[11]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[11]) );
  FD_1_440 FF_12 ( .D(D[12]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[12]) );
  FD_1_439 FF_13 ( .D(D[13]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[13]) );
  FD_1_438 FF_14 ( .D(D[14]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[14]) );
  FD_1_437 FF_15 ( .D(D[15]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[15]) );
  FD_1_436 FF_16 ( .D(D[16]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[16]) );
  FD_1_435 FF_17 ( .D(D[17]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[17]) );
  FD_1_434 FF_18 ( .D(D[18]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[18]) );
  FD_1_433 FF_19 ( .D(D[19]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[19]) );
  FD_1_432 FF_20 ( .D(D[20]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[20]) );
  FD_1_431 FF_21 ( .D(D[21]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[21]) );
  FD_1_430 FF_22 ( .D(D[22]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[22]) );
  FD_1_429 FF_23 ( .D(D[23]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[23]) );
  FD_1_428 FF_24 ( .D(D[24]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[24]) );
  FD_1_427 FF_25 ( .D(D[25]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[25]) );
  FD_1_426 FF_26 ( .D(D[26]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[26]) );
  FD_1_425 FF_27 ( .D(D[27]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[27]) );
  FD_1_424 FF_28 ( .D(D[28]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[28]) );
  FD_1_423 FF_29 ( .D(D[29]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[29]) );
  FD_1_422 FF_30 ( .D(D[30]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[30]) );
  FD_1_421 FF_31 ( .D(D[31]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[31]) );
  CLKBUF_X1 U1 ( .A(EN), .Z(n1) );
  CLKBUF_X1 U2 ( .A(EN), .Z(n2) );
  CLKBUF_X1 U3 ( .A(EN), .Z(n3) );
  BUF_X1 U4 ( .A(RST), .Z(n6) );
  BUF_X1 U5 ( .A(RST), .Z(n4) );
  BUF_X1 U6 ( .A(RST), .Z(n5) );
endmodule


module REG_N32_10 ( D, Q, EN, RST, CLK );
  input [31:0] D;
  output [31:0] Q;
  input EN, RST, CLK;
  wire   n1, n2, n3, n4, n5, n6;

  FD_1_415 FF_0 ( .D(D[0]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[0]) );
  FD_1_414 FF_1 ( .D(D[1]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[1]) );
  FD_1_413 FF_2 ( .D(D[2]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[2]) );
  FD_1_412 FF_3 ( .D(D[3]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[3]) );
  FD_1_411 FF_4 ( .D(D[4]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[4]) );
  FD_1_410 FF_5 ( .D(D[5]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[5]) );
  FD_1_409 FF_6 ( .D(D[6]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[6]) );
  FD_1_408 FF_7 ( .D(D[7]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[7]) );
  FD_1_407 FF_8 ( .D(D[8]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[8]) );
  FD_1_406 FF_9 ( .D(D[9]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[9]) );
  FD_1_405 FF_10 ( .D(D[10]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[10]) );
  FD_1_404 FF_11 ( .D(D[11]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[11]) );
  FD_1_403 FF_12 ( .D(D[12]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[12]) );
  FD_1_402 FF_13 ( .D(D[13]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[13]) );
  FD_1_401 FF_14 ( .D(D[14]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[14]) );
  FD_1_400 FF_15 ( .D(D[15]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[15]) );
  FD_1_399 FF_16 ( .D(D[16]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[16]) );
  FD_1_398 FF_17 ( .D(D[17]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[17]) );
  FD_1_397 FF_18 ( .D(D[18]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[18]) );
  FD_1_396 FF_19 ( .D(D[19]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[19]) );
  FD_1_395 FF_20 ( .D(D[20]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[20]) );
  FD_1_394 FF_21 ( .D(D[21]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[21]) );
  FD_1_393 FF_22 ( .D(D[22]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[22]) );
  FD_1_392 FF_23 ( .D(D[23]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[23]) );
  FD_1_391 FF_24 ( .D(D[24]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[24]) );
  FD_1_390 FF_25 ( .D(D[25]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[25]) );
  FD_1_389 FF_26 ( .D(D[26]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[26]) );
  FD_1_388 FF_27 ( .D(D[27]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[27]) );
  FD_1_387 FF_28 ( .D(D[28]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[28]) );
  FD_1_386 FF_29 ( .D(D[29]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[29]) );
  FD_1_385 FF_30 ( .D(D[30]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[30]) );
  FD_1_384 FF_31 ( .D(D[31]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[31]) );
  CLKBUF_X1 U1 ( .A(EN), .Z(n1) );
  CLKBUF_X1 U2 ( .A(EN), .Z(n2) );
  CLKBUF_X1 U3 ( .A(EN), .Z(n3) );
  BUF_X1 U4 ( .A(RST), .Z(n6) );
  BUF_X1 U5 ( .A(RST), .Z(n4) );
  BUF_X1 U6 ( .A(RST), .Z(n5) );
endmodule


module REG_N32_9 ( D, Q, EN, RST, CLK );
  input [31:0] D;
  output [31:0] Q;
  input EN, RST, CLK;
  wire   n1, n2, n3, n4, n5, n6;

  FD_1_378 FF_0 ( .D(D[0]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[0]) );
  FD_1_377 FF_1 ( .D(D[1]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[1]) );
  FD_1_376 FF_2 ( .D(D[2]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[2]) );
  FD_1_375 FF_3 ( .D(D[3]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[3]) );
  FD_1_374 FF_4 ( .D(D[4]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[4]) );
  FD_1_373 FF_5 ( .D(D[5]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[5]) );
  FD_1_372 FF_6 ( .D(D[6]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[6]) );
  FD_1_371 FF_7 ( .D(D[7]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[7]) );
  FD_1_370 FF_8 ( .D(D[8]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[8]) );
  FD_1_369 FF_9 ( .D(D[9]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[9]) );
  FD_1_368 FF_10 ( .D(D[10]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[10]) );
  FD_1_367 FF_11 ( .D(D[11]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[11]) );
  FD_1_366 FF_12 ( .D(D[12]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[12]) );
  FD_1_365 FF_13 ( .D(D[13]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[13]) );
  FD_1_364 FF_14 ( .D(D[14]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[14]) );
  FD_1_363 FF_15 ( .D(D[15]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[15]) );
  FD_1_362 FF_16 ( .D(D[16]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[16]) );
  FD_1_361 FF_17 ( .D(D[17]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[17]) );
  FD_1_360 FF_18 ( .D(D[18]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[18]) );
  FD_1_359 FF_19 ( .D(D[19]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[19]) );
  FD_1_358 FF_20 ( .D(D[20]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[20]) );
  FD_1_357 FF_21 ( .D(D[21]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[21]) );
  FD_1_356 FF_22 ( .D(D[22]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[22]) );
  FD_1_355 FF_23 ( .D(D[23]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[23]) );
  FD_1_354 FF_24 ( .D(D[24]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[24]) );
  FD_1_353 FF_25 ( .D(D[25]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[25]) );
  FD_1_352 FF_26 ( .D(D[26]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[26]) );
  FD_1_351 FF_27 ( .D(D[27]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[27]) );
  FD_1_350 FF_28 ( .D(D[28]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[28]) );
  FD_1_349 FF_29 ( .D(D[29]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[29]) );
  FD_1_348 FF_30 ( .D(D[30]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[30]) );
  FD_1_347 FF_31 ( .D(D[31]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[31]) );
  BUF_X1 U1 ( .A(EN), .Z(n3) );
  BUF_X1 U2 ( .A(EN), .Z(n1) );
  BUF_X1 U3 ( .A(EN), .Z(n2) );
  BUF_X1 U4 ( .A(RST), .Z(n6) );
  BUF_X1 U5 ( .A(RST), .Z(n5) );
  BUF_X1 U6 ( .A(RST), .Z(n4) );
endmodule


module REG_N32_8 ( D, Q, EN, RST, CLK );
  input [31:0] D;
  output [31:0] Q;
  input EN, RST, CLK;
  wire   n1, n2, n3, n4, n5, n6;

  FD_1_346 FF_0 ( .D(D[0]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[0]) );
  FD_1_345 FF_1 ( .D(D[1]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[1]) );
  FD_1_344 FF_2 ( .D(D[2]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[2]) );
  FD_1_343 FF_3 ( .D(D[3]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[3]) );
  FD_1_342 FF_4 ( .D(D[4]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[4]) );
  FD_1_341 FF_5 ( .D(D[5]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[5]) );
  FD_1_340 FF_6 ( .D(D[6]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[6]) );
  FD_1_339 FF_7 ( .D(D[7]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[7]) );
  FD_1_338 FF_8 ( .D(D[8]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[8]) );
  FD_1_337 FF_9 ( .D(D[9]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[9]) );
  FD_1_336 FF_10 ( .D(D[10]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[10]) );
  FD_1_335 FF_11 ( .D(D[11]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[11]) );
  FD_1_334 FF_12 ( .D(D[12]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[12]) );
  FD_1_333 FF_13 ( .D(D[13]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[13]) );
  FD_1_332 FF_14 ( .D(D[14]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[14]) );
  FD_1_331 FF_15 ( .D(D[15]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[15]) );
  FD_1_330 FF_16 ( .D(D[16]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[16]) );
  FD_1_329 FF_17 ( .D(D[17]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[17]) );
  FD_1_328 FF_18 ( .D(D[18]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[18]) );
  FD_1_327 FF_19 ( .D(D[19]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[19]) );
  FD_1_326 FF_20 ( .D(D[20]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[20]) );
  FD_1_325 FF_21 ( .D(D[21]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[21]) );
  FD_1_324 FF_22 ( .D(D[22]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[22]) );
  FD_1_323 FF_23 ( .D(D[23]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[23]) );
  FD_1_322 FF_24 ( .D(D[24]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[24]) );
  FD_1_321 FF_25 ( .D(D[25]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[25]) );
  FD_1_320 FF_26 ( .D(D[26]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[26]) );
  FD_1_319 FF_27 ( .D(D[27]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[27]) );
  FD_1_318 FF_28 ( .D(D[28]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[28]) );
  FD_1_317 FF_29 ( .D(D[29]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[29]) );
  FD_1_316 FF_30 ( .D(D[30]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[30]) );
  FD_1_315 FF_31 ( .D(D[31]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[31]) );
  BUF_X1 U1 ( .A(EN), .Z(n3) );
  BUF_X1 U2 ( .A(EN), .Z(n1) );
  BUF_X1 U3 ( .A(EN), .Z(n2) );
  BUF_X1 U4 ( .A(RST), .Z(n6) );
  BUF_X1 U5 ( .A(RST), .Z(n4) );
  BUF_X1 U6 ( .A(RST), .Z(n5) );
endmodule


module REG_N32_7 ( D, Q, EN, RST, CLK );
  input [31:0] D;
  output [31:0] Q;
  input EN, RST, CLK;
  wire   n1, n2, n3, n4, n5, n6;

  FD_1_314 FF_0 ( .D(D[0]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[0]) );
  FD_1_313 FF_1 ( .D(D[1]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[1]) );
  FD_1_312 FF_2 ( .D(D[2]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[2]) );
  FD_1_311 FF_3 ( .D(D[3]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[3]) );
  FD_1_310 FF_4 ( .D(D[4]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[4]) );
  FD_1_309 FF_5 ( .D(D[5]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[5]) );
  FD_1_308 FF_6 ( .D(D[6]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[6]) );
  FD_1_307 FF_7 ( .D(D[7]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[7]) );
  FD_1_306 FF_8 ( .D(D[8]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[8]) );
  FD_1_305 FF_9 ( .D(D[9]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[9]) );
  FD_1_304 FF_10 ( .D(D[10]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[10]) );
  FD_1_303 FF_11 ( .D(D[11]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[11]) );
  FD_1_302 FF_12 ( .D(D[12]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[12]) );
  FD_1_301 FF_13 ( .D(D[13]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[13]) );
  FD_1_300 FF_14 ( .D(D[14]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[14]) );
  FD_1_299 FF_15 ( .D(D[15]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[15]) );
  FD_1_298 FF_16 ( .D(D[16]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[16]) );
  FD_1_297 FF_17 ( .D(D[17]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[17]) );
  FD_1_296 FF_18 ( .D(D[18]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[18]) );
  FD_1_295 FF_19 ( .D(D[19]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[19]) );
  FD_1_294 FF_20 ( .D(D[20]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[20]) );
  FD_1_293 FF_21 ( .D(D[21]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[21]) );
  FD_1_292 FF_22 ( .D(D[22]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[22]) );
  FD_1_291 FF_23 ( .D(D[23]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[23]) );
  FD_1_290 FF_24 ( .D(D[24]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[24]) );
  FD_1_289 FF_25 ( .D(D[25]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[25]) );
  FD_1_288 FF_26 ( .D(D[26]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[26]) );
  FD_1_287 FF_27 ( .D(D[27]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[27]) );
  FD_1_286 FF_28 ( .D(D[28]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[28]) );
  FD_1_285 FF_29 ( .D(D[29]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[29]) );
  FD_1_284 FF_30 ( .D(D[30]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[30]) );
  FD_1_283 FF_31 ( .D(D[31]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[31]) );
  BUF_X1 U1 ( .A(EN), .Z(n3) );
  BUF_X1 U2 ( .A(EN), .Z(n1) );
  BUF_X1 U3 ( .A(EN), .Z(n2) );
  BUF_X1 U4 ( .A(RST), .Z(n6) );
  BUF_X1 U5 ( .A(RST), .Z(n4) );
  BUF_X1 U6 ( .A(RST), .Z(n5) );
endmodule


module REG_N32_6 ( D, Q, EN, RST, CLK );
  input [31:0] D;
  output [31:0] Q;
  input EN, RST, CLK;
  wire   n1, n2, n3, n4, n5, n6;

  FD_1_277 FF_0 ( .D(D[0]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[0]) );
  FD_1_276 FF_1 ( .D(D[1]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[1]) );
  FD_1_275 FF_2 ( .D(D[2]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[2]) );
  FD_1_274 FF_3 ( .D(D[3]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[3]) );
  FD_1_273 FF_4 ( .D(D[4]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[4]) );
  FD_1_272 FF_5 ( .D(D[5]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[5]) );
  FD_1_271 FF_6 ( .D(D[6]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[6]) );
  FD_1_270 FF_7 ( .D(D[7]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[7]) );
  FD_1_269 FF_8 ( .D(D[8]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[8]) );
  FD_1_268 FF_9 ( .D(D[9]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[9]) );
  FD_1_267 FF_10 ( .D(D[10]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[10]) );
  FD_1_266 FF_11 ( .D(D[11]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[11]) );
  FD_1_265 FF_12 ( .D(D[12]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[12]) );
  FD_1_264 FF_13 ( .D(D[13]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[13]) );
  FD_1_263 FF_14 ( .D(D[14]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[14]) );
  FD_1_262 FF_15 ( .D(D[15]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[15]) );
  FD_1_261 FF_16 ( .D(D[16]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[16]) );
  FD_1_260 FF_17 ( .D(D[17]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[17]) );
  FD_1_259 FF_18 ( .D(D[18]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[18]) );
  FD_1_258 FF_19 ( .D(D[19]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[19]) );
  FD_1_257 FF_20 ( .D(D[20]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[20]) );
  FD_1_256 FF_21 ( .D(D[21]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[21]) );
  FD_1_255 FF_22 ( .D(D[22]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[22]) );
  FD_1_254 FF_23 ( .D(D[23]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[23]) );
  FD_1_253 FF_24 ( .D(D[24]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[24]) );
  FD_1_252 FF_25 ( .D(D[25]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[25]) );
  FD_1_251 FF_26 ( .D(D[26]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[26]) );
  FD_1_250 FF_27 ( .D(D[27]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[27]) );
  FD_1_249 FF_28 ( .D(D[28]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[28]) );
  FD_1_248 FF_29 ( .D(D[29]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[29]) );
  FD_1_247 FF_30 ( .D(D[30]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[30]) );
  FD_1_246 FF_31 ( .D(D[31]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[31]) );
  BUF_X1 U1 ( .A(EN), .Z(n3) );
  BUF_X1 U2 ( .A(EN), .Z(n1) );
  BUF_X1 U3 ( .A(EN), .Z(n2) );
  BUF_X1 U4 ( .A(RST), .Z(n6) );
  BUF_X1 U5 ( .A(RST), .Z(n4) );
  BUF_X1 U6 ( .A(RST), .Z(n5) );
endmodule


module REG_N32_5 ( D, Q, EN, RST, CLK );
  input [31:0] D;
  output [31:0] Q;
  input EN, RST, CLK;
  wire   n1, n2, n3, n4, n5, n6;

  FD_1_245 FF_0 ( .D(D[0]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[0]) );
  FD_1_244 FF_1 ( .D(D[1]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[1]) );
  FD_1_243 FF_2 ( .D(D[2]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[2]) );
  FD_1_242 FF_3 ( .D(D[3]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[3]) );
  FD_1_241 FF_4 ( .D(D[4]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[4]) );
  FD_1_240 FF_5 ( .D(D[5]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[5]) );
  FD_1_239 FF_6 ( .D(D[6]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[6]) );
  FD_1_238 FF_7 ( .D(D[7]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[7]) );
  FD_1_237 FF_8 ( .D(D[8]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[8]) );
  FD_1_236 FF_9 ( .D(D[9]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[9]) );
  FD_1_235 FF_10 ( .D(D[10]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[10]) );
  FD_1_234 FF_11 ( .D(D[11]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[11]) );
  FD_1_233 FF_12 ( .D(D[12]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[12]) );
  FD_1_232 FF_13 ( .D(D[13]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[13]) );
  FD_1_231 FF_14 ( .D(D[14]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[14]) );
  FD_1_230 FF_15 ( .D(D[15]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[15]) );
  FD_1_229 FF_16 ( .D(D[16]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[16]) );
  FD_1_228 FF_17 ( .D(D[17]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[17]) );
  FD_1_227 FF_18 ( .D(D[18]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[18]) );
  FD_1_226 FF_19 ( .D(D[19]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[19]) );
  FD_1_225 FF_20 ( .D(D[20]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[20]) );
  FD_1_224 FF_21 ( .D(D[21]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[21]) );
  FD_1_223 FF_22 ( .D(D[22]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[22]) );
  FD_1_222 FF_23 ( .D(D[23]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[23]) );
  FD_1_221 FF_24 ( .D(D[24]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[24]) );
  FD_1_220 FF_25 ( .D(D[25]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[25]) );
  FD_1_219 FF_26 ( .D(D[26]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[26]) );
  FD_1_218 FF_27 ( .D(D[27]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[27]) );
  FD_1_217 FF_28 ( .D(D[28]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[28]) );
  FD_1_216 FF_29 ( .D(D[29]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[29]) );
  FD_1_215 FF_30 ( .D(D[30]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[30]) );
  FD_1_214 FF_31 ( .D(D[31]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[31]) );
  BUF_X1 U1 ( .A(EN), .Z(n3) );
  BUF_X1 U2 ( .A(EN), .Z(n1) );
  BUF_X1 U3 ( .A(EN), .Z(n2) );
  BUF_X1 U4 ( .A(RST), .Z(n6) );
  BUF_X1 U5 ( .A(RST), .Z(n4) );
  BUF_X1 U6 ( .A(RST), .Z(n5) );
endmodule


module REG_N32_4 ( D, Q, EN, RST, CLK );
  input [31:0] D;
  output [31:0] Q;
  input EN, RST, CLK;
  wire   n1, n2, n3, n4, n5, n6;

  FD_1_213 FF_0 ( .D(D[0]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[0]) );
  FD_1_212 FF_1 ( .D(D[1]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[1]) );
  FD_1_211 FF_2 ( .D(D[2]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[2]) );
  FD_1_210 FF_3 ( .D(D[3]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[3]) );
  FD_1_209 FF_4 ( .D(D[4]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[4]) );
  FD_1_208 FF_5 ( .D(D[5]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[5]) );
  FD_1_207 FF_6 ( .D(D[6]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[6]) );
  FD_1_206 FF_7 ( .D(D[7]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[7]) );
  FD_1_205 FF_8 ( .D(D[8]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[8]) );
  FD_1_204 FF_9 ( .D(D[9]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[9]) );
  FD_1_203 FF_10 ( .D(D[10]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[10]) );
  FD_1_202 FF_11 ( .D(D[11]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[11]) );
  FD_1_201 FF_12 ( .D(D[12]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[12]) );
  FD_1_200 FF_13 ( .D(D[13]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[13]) );
  FD_1_199 FF_14 ( .D(D[14]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[14]) );
  FD_1_198 FF_15 ( .D(D[15]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[15]) );
  FD_1_197 FF_16 ( .D(D[16]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[16]) );
  FD_1_196 FF_17 ( .D(D[17]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[17]) );
  FD_1_195 FF_18 ( .D(D[18]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[18]) );
  FD_1_194 FF_19 ( .D(D[19]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[19]) );
  FD_1_193 FF_20 ( .D(D[20]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[20]) );
  FD_1_192 FF_21 ( .D(D[21]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[21]) );
  FD_1_191 FF_22 ( .D(D[22]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[22]) );
  FD_1_190 FF_23 ( .D(D[23]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[23]) );
  FD_1_189 FF_24 ( .D(D[24]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[24]) );
  FD_1_188 FF_25 ( .D(D[25]), .CLK(CLK), .EN(n2), .RST(n5), .Q(Q[25]) );
  FD_1_187 FF_26 ( .D(D[26]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[26]) );
  FD_1_186 FF_27 ( .D(D[27]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[27]) );
  FD_1_185 FF_28 ( .D(D[28]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[28]) );
  FD_1_184 FF_29 ( .D(D[29]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[29]) );
  FD_1_183 FF_30 ( .D(D[30]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[30]) );
  FD_1_182 FF_31 ( .D(D[31]), .CLK(CLK), .EN(n3), .RST(n6), .Q(Q[31]) );
  BUF_X1 U1 ( .A(EN), .Z(n3) );
  BUF_X1 U2 ( .A(EN), .Z(n1) );
  BUF_X1 U3 ( .A(EN), .Z(n2) );
  BUF_X1 U4 ( .A(RST), .Z(n6) );
  BUF_X1 U5 ( .A(RST), .Z(n4) );
  BUF_X1 U6 ( .A(RST), .Z(n5) );
endmodule


module REG_N32_3 ( D, Q, EN, RST, CLK );
  input [31:0] D;
  output [31:0] Q;
  input EN, RST, CLK;
  wire   n1, n2, n3;

  FD_1_181 FF_0 ( .D(D[0]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[0]) );
  FD_1_180 FF_1 ( .D(D[1]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[1]) );
  FD_1_179 FF_2 ( .D(D[2]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[2]) );
  FD_1_178 FF_3 ( .D(D[3]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[3]) );
  FD_1_177 FF_4 ( .D(D[4]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[4]) );
  FD_1_176 FF_5 ( .D(D[5]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[5]) );
  FD_1_175 FF_6 ( .D(D[6]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[6]) );
  FD_1_174 FF_7 ( .D(D[7]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[7]) );
  FD_1_173 FF_8 ( .D(D[8]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[8]) );
  FD_1_172 FF_9 ( .D(D[9]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[9]) );
  FD_1_171 FF_10 ( .D(D[10]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[10]) );
  FD_1_170 FF_11 ( .D(D[11]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[11]) );
  FD_1_169 FF_12 ( .D(D[12]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[12]) );
  FD_1_168 FF_13 ( .D(D[13]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[13]) );
  FD_1_167 FF_14 ( .D(D[14]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[14]) );
  FD_1_166 FF_15 ( .D(D[15]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[15]) );
  FD_1_165 FF_16 ( .D(D[16]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[16]) );
  FD_1_164 FF_17 ( .D(D[17]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[17]) );
  FD_1_163 FF_18 ( .D(D[18]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[18]) );
  FD_1_162 FF_19 ( .D(D[19]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[19]) );
  FD_1_161 FF_20 ( .D(D[20]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[20]) );
  FD_1_160 FF_21 ( .D(D[21]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[21]) );
  FD_1_159 FF_22 ( .D(D[22]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[22]) );
  FD_1_158 FF_23 ( .D(D[23]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[23]) );
  FD_1_157 FF_24 ( .D(D[24]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[24]) );
  FD_1_156 FF_25 ( .D(D[25]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[25]) );
  FD_1_155 FF_26 ( .D(D[26]), .CLK(CLK), .EN(EN), .RST(n3), .Q(Q[26]) );
  FD_1_154 FF_27 ( .D(D[27]), .CLK(CLK), .EN(EN), .RST(n3), .Q(Q[27]) );
  FD_1_153 FF_28 ( .D(D[28]), .CLK(CLK), .EN(EN), .RST(n3), .Q(Q[28]) );
  FD_1_152 FF_29 ( .D(D[29]), .CLK(CLK), .EN(EN), .RST(n3), .Q(Q[29]) );
  FD_1_151 FF_30 ( .D(D[30]), .CLK(CLK), .EN(EN), .RST(n3), .Q(Q[30]) );
  FD_1_150 FF_31 ( .D(D[31]), .CLK(CLK), .EN(EN), .RST(n3), .Q(Q[31]) );
  BUF_X1 U1 ( .A(RST), .Z(n1) );
  BUF_X1 U2 ( .A(RST), .Z(n2) );
  BUF_X1 U3 ( .A(RST), .Z(n3) );
endmodule


module REG_N32_2 ( D, Q, EN, RST, CLK );
  input [31:0] D;
  output [31:0] Q;
  input EN, RST, CLK;
  wire   n1, n2, n3, n4, n5, n6;

  FD_1_147 FF_0 ( .D(D[0]), .CLK(CLK), .EN(n4), .RST(n2), .Q(Q[0]) );
  FD_1_146 FF_1 ( .D(D[1]), .CLK(CLK), .EN(n4), .RST(n2), .Q(Q[1]) );
  FD_1_145 FF_2 ( .D(D[2]), .CLK(CLK), .EN(n4), .RST(n2), .Q(Q[2]) );
  FD_1_144 FF_3 ( .D(D[3]), .CLK(CLK), .EN(n4), .RST(n2), .Q(Q[3]) );
  FD_1_143 FF_4 ( .D(D[4]), .CLK(CLK), .EN(n4), .RST(n2), .Q(Q[4]) );
  FD_1_142 FF_5 ( .D(D[5]), .CLK(CLK), .EN(n4), .RST(n2), .Q(Q[5]) );
  FD_1_141 FF_6 ( .D(D[6]), .CLK(CLK), .EN(n4), .RST(n2), .Q(Q[6]) );
  FD_1_140 FF_7 ( .D(D[7]), .CLK(CLK), .EN(n4), .RST(n2), .Q(Q[7]) );
  FD_1_139 FF_8 ( .D(D[8]), .CLK(CLK), .EN(n4), .RST(n2), .Q(Q[8]) );
  FD_1_138 FF_9 ( .D(D[9]), .CLK(CLK), .EN(n4), .RST(n3), .Q(Q[9]) );
  FD_1_137 FF_10 ( .D(D[10]), .CLK(CLK), .EN(n4), .RST(n3), .Q(Q[10]) );
  FD_1_136 FF_11 ( .D(D[11]), .CLK(CLK), .EN(n4), .RST(n3), .Q(Q[11]) );
  FD_1_135 FF_12 ( .D(D[12]), .CLK(CLK), .EN(n4), .RST(n1), .Q(Q[12]) );
  FD_1_134 FF_13 ( .D(D[13]), .CLK(CLK), .EN(n5), .RST(n1), .Q(Q[13]) );
  FD_1_133 FF_14 ( .D(D[14]), .CLK(CLK), .EN(n5), .RST(n1), .Q(Q[14]) );
  FD_1_132 FF_15 ( .D(D[15]), .CLK(CLK), .EN(n5), .RST(n1), .Q(Q[15]) );
  FD_1_131 FF_16 ( .D(D[16]), .CLK(CLK), .EN(n5), .RST(n1), .Q(Q[16]) );
  FD_1_130 FF_17 ( .D(D[17]), .CLK(CLK), .EN(n5), .RST(n1), .Q(Q[17]) );
  FD_1_129 FF_18 ( .D(D[18]), .CLK(CLK), .EN(n5), .RST(n1), .Q(Q[18]) );
  FD_1_128 FF_19 ( .D(D[19]), .CLK(CLK), .EN(n5), .RST(n1), .Q(Q[19]) );
  FD_1_127 FF_20 ( .D(D[20]), .CLK(CLK), .EN(n5), .RST(n1), .Q(Q[20]) );
  FD_1_126 FF_21 ( .D(D[21]), .CLK(CLK), .EN(n5), .RST(n1), .Q(Q[21]) );
  FD_1_125 FF_22 ( .D(D[22]), .CLK(CLK), .EN(n5), .RST(n1), .Q(Q[22]) );
  FD_1_124 FF_23 ( .D(D[23]), .CLK(CLK), .EN(n5), .RST(n2), .Q(Q[23]) );
  FD_1_123 FF_24 ( .D(D[24]), .CLK(CLK), .EN(n5), .RST(n2), .Q(Q[24]) );
  FD_1_122 FF_25 ( .D(D[25]), .CLK(CLK), .EN(n5), .RST(n2), .Q(Q[25]) );
  FD_1_121 FF_26 ( .D(D[26]), .CLK(CLK), .EN(n6), .RST(n2), .Q(Q[26]) );
  FD_1_120 FF_27 ( .D(D[27]), .CLK(CLK), .EN(n6), .RST(n1), .Q(Q[27]) );
  FD_1_119 FF_28 ( .D(D[28]), .CLK(CLK), .EN(n6), .RST(n1), .Q(Q[28]) );
  FD_1_118 FF_29 ( .D(D[29]), .CLK(CLK), .EN(n6), .RST(n3), .Q(Q[29]) );
  FD_1_117 FF_30 ( .D(D[30]), .CLK(CLK), .EN(n6), .RST(n3), .Q(Q[30]) );
  FD_1_116 FF_31 ( .D(D[31]), .CLK(CLK), .EN(n6), .RST(n3), .Q(Q[31]) );
  BUF_X1 U1 ( .A(EN), .Z(n6) );
  BUF_X1 U2 ( .A(EN), .Z(n4) );
  BUF_X1 U3 ( .A(EN), .Z(n5) );
  BUF_X1 U4 ( .A(RST), .Z(n2) );
  BUF_X1 U5 ( .A(RST), .Z(n1) );
  BUF_X1 U6 ( .A(RST), .Z(n3) );
endmodule


module REG_N32_1 ( D, Q, EN, RST, CLK );
  input [31:0] D;
  output [31:0] Q;
  input EN, RST, CLK;
  wire   n1, n2, n3;

  FD_1_97 FF_0 ( .D(D[0]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[0]) );
  FD_1_96 FF_1 ( .D(D[1]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[1]) );
  FD_1_95 FF_2 ( .D(D[2]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[2]) );
  FD_1_94 FF_3 ( .D(D[3]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[3]) );
  FD_1_93 FF_4 ( .D(D[4]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[4]) );
  FD_1_92 FF_5 ( .D(D[5]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[5]) );
  FD_1_91 FF_6 ( .D(D[6]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[6]) );
  FD_1_90 FF_7 ( .D(D[7]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[7]) );
  FD_1_89 FF_8 ( .D(D[8]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[8]) );
  FD_1_88 FF_9 ( .D(D[9]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[9]) );
  FD_1_87 FF_10 ( .D(D[10]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[10]) );
  FD_1_86 FF_11 ( .D(D[11]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[11]) );
  FD_1_85 FF_12 ( .D(D[12]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[12]) );
  FD_1_84 FF_13 ( .D(D[13]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[13]) );
  FD_1_83 FF_14 ( .D(D[14]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[14]) );
  FD_1_82 FF_15 ( .D(D[15]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[15]) );
  FD_1_81 FF_16 ( .D(D[16]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[16]) );
  FD_1_80 FF_17 ( .D(D[17]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[17]) );
  FD_1_79 FF_18 ( .D(D[18]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[18]) );
  FD_1_78 FF_19 ( .D(D[19]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[19]) );
  FD_1_77 FF_20 ( .D(D[20]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[20]) );
  FD_1_76 FF_21 ( .D(D[21]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[21]) );
  FD_1_75 FF_22 ( .D(D[22]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[22]) );
  FD_1_74 FF_23 ( .D(D[23]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[23]) );
  FD_1_73 FF_24 ( .D(D[24]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[24]) );
  FD_1_72 FF_25 ( .D(D[25]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[25]) );
  FD_1_71 FF_26 ( .D(D[26]), .CLK(CLK), .EN(EN), .RST(n3), .Q(Q[26]) );
  FD_1_70 FF_27 ( .D(D[27]), .CLK(CLK), .EN(EN), .RST(n3), .Q(Q[27]) );
  FD_1_69 FF_28 ( .D(D[28]), .CLK(CLK), .EN(EN), .RST(n3), .Q(Q[28]) );
  FD_1_68 FF_29 ( .D(D[29]), .CLK(CLK), .EN(EN), .RST(n3), .Q(Q[29]) );
  FD_1_67 FF_30 ( .D(D[30]), .CLK(CLK), .EN(EN), .RST(n3), .Q(Q[30]) );
  FD_1_66 FF_31 ( .D(D[31]), .CLK(CLK), .EN(EN), .RST(n3), .Q(Q[31]) );
  BUF_X1 U1 ( .A(RST), .Z(n1) );
  BUF_X1 U2 ( .A(RST), .Z(n2) );
  BUF_X1 U3 ( .A(RST), .Z(n3) );
endmodule


module FD_181 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_180 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_179 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_178 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_177 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_176 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_175 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_174 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_173 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_172 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_171 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_170 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_169 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_168 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_167 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_166 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_165 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_164 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_163 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_162 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_161 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_160 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_159 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n3, n4;

  DFF_X1 Q_reg ( .D(n3), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n4), .ZN(n3) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n1), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n1) );
endmodule


module FD_158 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_157 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_156 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_155 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_154 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_153 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_152 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_151 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_150 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_149 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_148 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_147 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_146 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_145 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_144 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_143 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_142 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_141 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_140 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_139 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_138 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_137 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_136 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_135 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_134 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_133 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_132 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_131 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_130 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_129 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_128 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_127 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_126 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n2, n3;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  AND2_X1 U3 ( .A1(n2), .A2(n3), .ZN(n1) );
  INV_X1 U4 ( .A(RST), .ZN(n2) );
  MUX2_X1 U5 ( .A(Q), .B(D), .S(EN), .Z(n3) );
endmodule


module FD_125 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n2, n3, n4;

  DFF_X1 Q_reg ( .D(n4), .CK(CLK), .Q(Q) );
  MUX2_X2 U3 ( .A(Q), .B(D), .S(EN), .Z(n2) );
  INV_X1 U4 ( .A(RST), .ZN(n1) );
  NAND2_X1 U5 ( .A1(n2), .A2(n1), .ZN(n3) );
  INV_X1 U6 ( .A(n3), .ZN(n4) );
endmodule


module FD_124 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n2, n3, n4, n5, n6, n7, n8;

  DFF_X1 Q_reg ( .D(n6), .CK(CLK), .Q(Q) );
  INV_X1 U3 ( .A(RST), .ZN(n5) );
  NAND2_X1 U4 ( .A1(D), .A2(n4), .ZN(n2) );
  NAND2_X1 U5 ( .A1(n2), .A2(n3), .ZN(n6) );
  OR2_X1 U6 ( .A1(RST), .A2(n7), .ZN(n3) );
  AND2_X1 U7 ( .A1(EN), .A2(n5), .ZN(n4) );
  NAND2_X1 U8 ( .A1(Q), .A2(n8), .ZN(n7) );
  INV_X1 U9 ( .A(EN), .ZN(n8) );
endmodule


module FD_123 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_122 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_121 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_120 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_119 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_118 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_117 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_116 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_115 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_114 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_113 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_112 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_111 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_110 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_109 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_108 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_107 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_106 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_105 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_104 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_103 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_102 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n9, n1, n6, n7, n8;

  DFF_X1 Q_reg ( .D(n6), .CK(CLK), .Q(n9), .QN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(Q) );
  NOR2_X1 U4 ( .A1(RST), .A2(n8), .ZN(n6) );
  AOI22_X1 U5 ( .A1(EN), .A2(D), .B1(n9), .B2(n7), .ZN(n8) );
  INV_X1 U6 ( .A(EN), .ZN(n7) );
endmodule


module FD_101 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_100 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_99 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_98 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_97 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_96 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_95 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_94 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_93 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_92 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_91 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_90 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_89 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_88 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_87 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_86 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_85 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_84 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_83 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_82 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_81 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_80 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_79 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_78 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_77 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_76 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_75 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_74 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_73 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_72 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_71 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_70 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_69 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_68 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_67 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_66 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_65 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_64 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_63 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_62 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_61 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_60 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_59 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_58 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_57 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_56 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_55 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_54 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_53 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_52 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_51 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_50 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n2, n3;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  AND2_X1 U3 ( .A1(n2), .A2(n3), .ZN(n1) );
  INV_X1 U4 ( .A(RST), .ZN(n2) );
  MUX2_X1 U5 ( .A(Q), .B(D), .S(EN), .Z(n3) );
endmodule


module FD_49 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n2, n3, n4, n5, n6, n7;

  DFF_X1 Q_reg ( .D(n6), .CK(CLK), .Q(Q) );
  AND2_X1 U3 ( .A1(EN), .A2(n7), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Q), .A2(n4), .ZN(n5) );
  NAND2_X1 U5 ( .A1(D), .A2(n3), .ZN(n1) );
  NAND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(n6) );
  OR2_X1 U7 ( .A1(RST), .A2(n5), .ZN(n2) );
  INV_X1 U8 ( .A(EN), .ZN(n4) );
  INV_X1 U9 ( .A(RST), .ZN(n7) );
endmodule


module FD_48 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_47 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_46 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_45 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_44 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_43 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_42 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_41 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_40 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_39 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_38 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_37 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_36 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_35 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_34 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_33 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_32 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_31 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_30 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_29 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_28 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_27 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_26 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_25 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_24 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_23 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_22 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_21 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_20 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_19 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_18 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_17 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_16 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_15 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_14 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_13 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_12 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_11 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_10 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_9 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_8 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_7 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_6 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_5 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_4 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_3 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_2 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module FD_1 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n1, n4, n5;

  DFF_X1 Q_reg ( .D(n1), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n5), .ZN(n1) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U5 ( .A(EN), .ZN(n4) );
endmodule


module GENERAL_PROPAGATE_0 ( Pi, Po );
  input [1:0] Pi;
  output Po;


  AND_GATE_1_440 AND_INST ( .A(Pi[1]), .B(Pi[0]), .Y(Po) );
endmodule


module MUX41_GEN_N16_0 ( A, B, C, D, SEL, Y );
  input [15:0] A;
  input [15:0] B;
  input [15:0] C;
  input [15:0] D;
  input [1:0] SEL;
  output [15:0] Y;
  wire   n3, n4, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n1;

  NAND2_X1 U38 ( .A1(n3), .A2(n4), .ZN(Y[9]) );
  NAND2_X1 U39 ( .A1(n9), .A2(n10), .ZN(Y[8]) );
  NAND2_X1 U40 ( .A1(n11), .A2(n12), .ZN(Y[7]) );
  NAND2_X1 U41 ( .A1(n13), .A2(n14), .ZN(Y[6]) );
  NAND2_X1 U42 ( .A1(n15), .A2(n16), .ZN(Y[5]) );
  NAND2_X1 U43 ( .A1(n17), .A2(n18), .ZN(Y[4]) );
  NAND2_X1 U44 ( .A1(n19), .A2(n20), .ZN(Y[3]) );
  NAND2_X1 U45 ( .A1(n21), .A2(n22), .ZN(Y[2]) );
  NAND2_X1 U46 ( .A1(n23), .A2(n24), .ZN(Y[1]) );
  NAND2_X1 U47 ( .A1(n25), .A2(n26), .ZN(Y[15]) );
  NAND2_X1 U48 ( .A1(n27), .A2(n28), .ZN(Y[14]) );
  NAND2_X1 U49 ( .A1(n29), .A2(n30), .ZN(Y[13]) );
  NAND2_X1 U50 ( .A1(n31), .A2(n32), .ZN(Y[12]) );
  NAND2_X1 U51 ( .A1(n33), .A2(n34), .ZN(Y[11]) );
  NAND2_X1 U52 ( .A1(n35), .A2(n36), .ZN(Y[10]) );
  NAND2_X1 U53 ( .A1(n37), .A2(n38), .ZN(Y[0]) );
  AND2_X2 U1 ( .A1(SEL[0]), .A2(SEL[1]), .ZN(n8) );
  NOR2_X2 U2 ( .A1(n39), .A2(SEL[1]), .ZN(n1) );
  NOR3_X2 U3 ( .A1(n1), .A2(n8), .A3(n5), .ZN(n7) );
  AND2_X1 U4 ( .A1(SEL[1]), .A2(n39), .ZN(n5) );
  INV_X1 U5 ( .A(SEL[0]), .ZN(n39) );
  AOI22_X1 U6 ( .A1(D[13]), .A2(n7), .B1(A[13]), .B2(n8), .ZN(n29) );
  AOI22_X1 U7 ( .A1(D[11]), .A2(n7), .B1(A[11]), .B2(n8), .ZN(n33) );
  AOI22_X1 U8 ( .A1(D[12]), .A2(n7), .B1(A[12]), .B2(n8), .ZN(n31) );
  AOI22_X1 U9 ( .A1(D[10]), .A2(n7), .B1(A[10]), .B2(n8), .ZN(n35) );
  AOI22_X1 U10 ( .A1(D[7]), .A2(n7), .B1(A[7]), .B2(n8), .ZN(n11) );
  AOI22_X1 U11 ( .A1(D[15]), .A2(n7), .B1(A[15]), .B2(n8), .ZN(n25) );
  AOI22_X1 U12 ( .A1(D[6]), .A2(n7), .B1(A[6]), .B2(n8), .ZN(n13) );
  AOI22_X1 U13 ( .A1(D[9]), .A2(n7), .B1(A[9]), .B2(n8), .ZN(n3) );
  AOI22_X1 U14 ( .A1(D[8]), .A2(n7), .B1(A[8]), .B2(n8), .ZN(n9) );
  AOI22_X1 U15 ( .A1(D[5]), .A2(n7), .B1(A[5]), .B2(n8), .ZN(n15) );
  AOI22_X1 U16 ( .A1(D[4]), .A2(n7), .B1(A[4]), .B2(n8), .ZN(n17) );
  AOI22_X1 U17 ( .A1(D[3]), .A2(n7), .B1(A[3]), .B2(n8), .ZN(n19) );
  AOI22_X1 U18 ( .A1(D[2]), .A2(n7), .B1(A[2]), .B2(n8), .ZN(n21) );
  AOI22_X1 U19 ( .A1(D[0]), .A2(n7), .B1(A[0]), .B2(n8), .ZN(n37) );
  AOI22_X1 U20 ( .A1(D[1]), .A2(n7), .B1(A[1]), .B2(n8), .ZN(n23) );
  AOI22_X1 U21 ( .A1(D[14]), .A2(n7), .B1(A[14]), .B2(n8), .ZN(n27) );
  AOI22_X1 U22 ( .A1(B[0]), .A2(n5), .B1(C[0]), .B2(n1), .ZN(n38) );
  AOI22_X1 U23 ( .A1(B[1]), .A2(n5), .B1(C[1]), .B2(n1), .ZN(n24) );
  AOI22_X1 U24 ( .A1(B[2]), .A2(n5), .B1(C[2]), .B2(n1), .ZN(n22) );
  AOI22_X1 U25 ( .A1(B[3]), .A2(n5), .B1(C[3]), .B2(n1), .ZN(n20) );
  AOI22_X1 U26 ( .A1(B[4]), .A2(n5), .B1(C[4]), .B2(n1), .ZN(n18) );
  AOI22_X1 U27 ( .A1(B[5]), .A2(n5), .B1(C[5]), .B2(n1), .ZN(n16) );
  AOI22_X1 U28 ( .A1(B[6]), .A2(n5), .B1(C[6]), .B2(n1), .ZN(n14) );
  AOI22_X1 U29 ( .A1(B[7]), .A2(n5), .B1(C[7]), .B2(n1), .ZN(n12) );
  AOI22_X1 U30 ( .A1(B[8]), .A2(n5), .B1(C[8]), .B2(n1), .ZN(n10) );
  AOI22_X1 U31 ( .A1(B[9]), .A2(n5), .B1(C[9]), .B2(n1), .ZN(n4) );
  AOI22_X1 U32 ( .A1(B[10]), .A2(n5), .B1(C[10]), .B2(n1), .ZN(n36) );
  AOI22_X1 U33 ( .A1(B[11]), .A2(n5), .B1(C[11]), .B2(n1), .ZN(n34) );
  AOI22_X1 U34 ( .A1(B[12]), .A2(n5), .B1(C[12]), .B2(n1), .ZN(n32) );
  AOI22_X1 U35 ( .A1(B[13]), .A2(n5), .B1(C[13]), .B2(n1), .ZN(n30) );
  AOI22_X1 U36 ( .A1(B[14]), .A2(n5), .B1(C[14]), .B2(n1), .ZN(n28) );
  AOI22_X1 U37 ( .A1(B[15]), .A2(n5), .B1(C[15]), .B2(n1), .ZN(n26) );
endmodule


module REG_N16_1_0 ( D, Q, EN, RST, CLK );
  input [15:0] D;
  output [15:0] Q;
  input EN, RST, CLK;
  wire   n1, n2, n3, n4;

  FD_1_64 FF_0 ( .D(D[0]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[0]) );
  FD_1_63 FF_1 ( .D(D[1]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[1]) );
  FD_1_62 FF_2 ( .D(D[2]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[2]) );
  FD_1_61 FF_3 ( .D(D[3]), .CLK(CLK), .EN(n1), .RST(n3), .Q(Q[3]) );
  FD_1_60 FF_4 ( .D(D[4]), .CLK(CLK), .EN(n1), .RST(n3), .Q(Q[4]) );
  FD_1_59 FF_5 ( .D(D[5]), .CLK(CLK), .EN(n1), .RST(n3), .Q(Q[5]) );
  FD_1_58 FF_6 ( .D(D[6]), .CLK(CLK), .EN(n1), .RST(n3), .Q(Q[6]) );
  FD_1_57 FF_7 ( .D(D[7]), .CLK(CLK), .EN(n1), .RST(n3), .Q(Q[7]) );
  FD_1_56 FF_8 ( .D(D[8]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[8]) );
  FD_1_55 FF_9 ( .D(D[9]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[9]) );
  FD_1_54 FF_10 ( .D(D[10]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[10]) );
  FD_1_53 FF_11 ( .D(D[11]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[11]) );
  FD_1_52 FF_12 ( .D(D[12]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[12]) );
  FD_1_51 FF_13 ( .D(D[13]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[13]) );
  FD_1_50 FF_14 ( .D(D[14]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[14]) );
  FD_1_49 FF_15 ( .D(D[15]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[15]) );
  BUF_X1 U1 ( .A(RST), .Z(n3) );
  BUF_X1 U2 ( .A(RST), .Z(n4) );
  CLKBUF_X1 U3 ( .A(EN), .Z(n1) );
  CLKBUF_X1 U4 ( .A(EN), .Z(n2) );
endmodule


module MUX21_GEN_N16_0 ( A, B, SEL, Y );
  input [15:0] A;
  input [15:0] B;
  output [15:0] Y;
  input SEL;
  wire   SB;
  wire   [15:0] Y1;
  wire   [15:0] Y2;

  INV_1_11 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_240 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_239 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_238 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_237 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_236 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_235 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_234 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_233 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_232 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_231 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_230 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_229 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_228 UND1_4 ( .A(A[4]), .B(SEL), .Y(Y1[4]) );
  NAND_GATE_227 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  NAND_GATE_226 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_225 UND1_5 ( .A(A[5]), .B(SEL), .Y(Y1[5]) );
  NAND_GATE_224 UND2_5 ( .A(B[5]), .B(SB), .Y(Y2[5]) );
  NAND_GATE_223 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_222 UND1_6 ( .A(A[6]), .B(SEL), .Y(Y1[6]) );
  NAND_GATE_221 UND2_6 ( .A(B[6]), .B(SB), .Y(Y2[6]) );
  NAND_GATE_220 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_219 UND1_7 ( .A(A[7]), .B(SEL), .Y(Y1[7]) );
  NAND_GATE_218 UND2_7 ( .A(B[7]), .B(SB), .Y(Y2[7]) );
  NAND_GATE_217 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  NAND_GATE_216 UND1_8 ( .A(A[8]), .B(SEL), .Y(Y1[8]) );
  NAND_GATE_215 UND2_8 ( .A(B[8]), .B(SB), .Y(Y2[8]) );
  NAND_GATE_214 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  NAND_GATE_213 UND1_9 ( .A(A[9]), .B(SEL), .Y(Y1[9]) );
  NAND_GATE_212 UND2_9 ( .A(B[9]), .B(SB), .Y(Y2[9]) );
  NAND_GATE_211 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  NAND_GATE_210 UND1_10 ( .A(A[10]), .B(SEL), .Y(Y1[10]) );
  NAND_GATE_209 UND2_10 ( .A(B[10]), .B(SB), .Y(Y2[10]) );
  NAND_GATE_208 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  NAND_GATE_207 UND1_11 ( .A(A[11]), .B(SEL), .Y(Y1[11]) );
  NAND_GATE_206 UND2_11 ( .A(B[11]), .B(SB), .Y(Y2[11]) );
  NAND_GATE_205 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  NAND_GATE_204 UND1_12 ( .A(A[12]), .B(SEL), .Y(Y1[12]) );
  NAND_GATE_203 UND2_12 ( .A(B[12]), .B(SB), .Y(Y2[12]) );
  NAND_GATE_202 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  NAND_GATE_201 UND1_13 ( .A(A[13]), .B(SEL), .Y(Y1[13]) );
  NAND_GATE_200 UND2_13 ( .A(B[13]), .B(SB), .Y(Y2[13]) );
  NAND_GATE_199 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  NAND_GATE_198 UND1_14 ( .A(A[14]), .B(SEL), .Y(Y1[14]) );
  NAND_GATE_197 UND2_14 ( .A(B[14]), .B(SB), .Y(Y2[14]) );
  NAND_GATE_196 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  NAND_GATE_195 UND1_15 ( .A(A[15]), .B(SEL), .Y(Y1[15]) );
  NAND_GATE_194 UND2_15 ( .A(B[15]), .B(SB), .Y(Y2[15]) );
  NAND_GATE_193 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
endmodule


module BOOTH_ENCODER_0 ( TO_ENC, ENC );
  input [2:0] TO_ENC;
  output [2:0] ENC;
  wire   n1, n2, n3, n4;

  INV_X1 U1 ( .A(TO_ENC[1]), .ZN(n3) );
  NAND2_X2 U2 ( .A1(TO_ENC[1]), .A2(TO_ENC[0]), .ZN(n2) );
  OAI21_X1 U3 ( .B1(TO_ENC[0]), .B2(TO_ENC[1]), .A(n1), .ZN(ENC[0]) );
  XNOR2_X2 U4 ( .A(n2), .B(n1), .ZN(ENC[1]) );
  INV_X2 U5 ( .A(TO_ENC[2]), .ZN(n1) );
  INV_X1 U6 ( .A(TO_ENC[0]), .ZN(n4) );
  NAND3_X1 U7 ( .A1(TO_ENC[2]), .A2(n4), .A3(n3), .ZN(ENC[2]) );
endmodule


module RCA_GEN_NO_C_N19_0 ( A, B, S, Co );
  input [18:0] A;
  input [18:0] B;
  output [18:0] S;
  output Co;

  wire   [17:0] CTMP;

  HA_7 HA_INST ( .A(A[0]), .B(B[0]), .S(S[0]), .Co(CTMP[0]) );
  FA_190 FAI_0 ( .A(A[1]), .B(B[1]), .Ci(CTMP[0]), .S(S[1]), .Co(CTMP[1]) );
  FA_189 FAI_1 ( .A(A[2]), .B(B[2]), .Ci(CTMP[1]), .S(S[2]), .Co(CTMP[2]) );
  FA_188 FAI_2 ( .A(A[3]), .B(B[3]), .Ci(CTMP[2]), .S(S[3]), .Co(CTMP[3]) );
  FA_187 FAI_3 ( .A(A[4]), .B(B[4]), .Ci(CTMP[3]), .S(S[4]), .Co(CTMP[4]) );
  FA_186 FAI_4 ( .A(A[5]), .B(B[5]), .Ci(CTMP[4]), .S(S[5]), .Co(CTMP[5]) );
  FA_185 FAI_5 ( .A(A[6]), .B(B[6]), .Ci(CTMP[5]), .S(S[6]), .Co(CTMP[6]) );
  FA_184 FAI_6 ( .A(A[7]), .B(B[7]), .Ci(CTMP[6]), .S(S[7]), .Co(CTMP[7]) );
  FA_183 FAI_7 ( .A(A[8]), .B(B[8]), .Ci(CTMP[7]), .S(S[8]), .Co(CTMP[8]) );
  FA_182 FAI_8 ( .A(A[9]), .B(B[9]), .Ci(CTMP[8]), .S(S[9]), .Co(CTMP[9]) );
  FA_181 FAI_9 ( .A(A[10]), .B(B[10]), .Ci(CTMP[9]), .S(S[10]), .Co(CTMP[10])
         );
  FA_180 FAI_10 ( .A(A[11]), .B(B[11]), .Ci(CTMP[10]), .S(S[11]), .Co(CTMP[11]) );
  FA_179 FAI_11 ( .A(A[12]), .B(B[12]), .Ci(CTMP[11]), .S(S[12]), .Co(CTMP[12]) );
  FA_178 FAI_12 ( .A(A[13]), .B(B[13]), .Ci(CTMP[12]), .S(S[13]), .Co(CTMP[13]) );
  FA_177 FAI_13 ( .A(A[14]), .B(B[14]), .Ci(CTMP[13]), .S(S[14]), .Co(CTMP[14]) );
  FA_176 FAI_14 ( .A(A[15]), .B(B[15]), .Ci(CTMP[14]), .S(S[15]), .Co(CTMP[15]) );
  FA_175 FAI_15 ( .A(A[16]), .B(B[16]), .Ci(CTMP[15]), .S(S[16]), .Co(CTMP[16]) );
  FA_174 FAI_16 ( .A(A[17]), .B(B[17]), .Ci(CTMP[16]), .S(S[17]), .Co(CTMP[17]) );
  FA_173 FAI_17 ( .A(A[18]), .B(B[18]), .Ci(CTMP[17]), .S(S[18]), .Co(Co) );
endmodule


module MUX51_GEN_N19_0 ( A, B, C, D, E, SEL, Y );
  input [18:0] A;
  input [18:0] B;
  input [18:0] C;
  input [18:0] D;
  input [18:0] E;
  input [2:0] SEL;
  output [18:0] Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98;

  BUF_X2 U1 ( .A(n93), .Z(n3) );
  NAND2_X4 U2 ( .A1(C[15]), .A2(n94), .ZN(n81) );
  NAND4_X2 U3 ( .A1(n83), .A2(n82), .A3(n81), .A4(n80), .ZN(Y[15]) );
  NAND2_X2 U4 ( .A1(C[11]), .A2(n94), .ZN(n62) );
  NAND2_X4 U5 ( .A1(C[13]), .A2(n94), .ZN(n72) );
  NAND4_X2 U6 ( .A1(n64), .A2(n63), .A3(n62), .A4(n61), .ZN(Y[11]) );
  NAND2_X2 U7 ( .A1(C[14]), .A2(n94), .ZN(n76) );
  NAND4_X2 U8 ( .A1(n78), .A2(n77), .A3(n76), .A4(n75), .ZN(Y[14]) );
  NAND2_X1 U9 ( .A1(C[10]), .A2(n94), .ZN(n57) );
  NAND4_X1 U10 ( .A1(n59), .A2(n58), .A3(n57), .A4(n56), .ZN(Y[10]) );
  NAND4_X2 U11 ( .A1(n74), .A2(n73), .A3(n72), .A4(n71), .ZN(Y[13]) );
  NAND3_X1 U12 ( .A1(n18), .A2(n17), .A3(n16), .ZN(Y[1]) );
  AOI22_X1 U13 ( .A1(E[2]), .A2(n3), .B1(B[2]), .B2(n92), .ZN(n19) );
  NAND2_X1 U14 ( .A1(C[6]), .A2(n94), .ZN(n37) );
  NAND2_X1 U15 ( .A1(C[9]), .A2(n94), .ZN(n52) );
  NOR2_X1 U16 ( .A1(n11), .A2(n10), .ZN(n93) );
  NAND3_X1 U17 ( .A1(SEL[2]), .A2(n8), .A3(n7), .ZN(n91) );
  BUF_X2 U18 ( .A(n91), .Z(n2) );
  INV_X2 U19 ( .A(SEL[1]), .ZN(n7) );
  AOI22_X2 U20 ( .A1(E[1]), .A2(n93), .B1(B[1]), .B2(n92), .ZN(n16) );
  INV_X2 U21 ( .A(n12), .ZN(n92) );
  INV_X1 U22 ( .A(n9), .ZN(n1) );
  AOI22_X2 U23 ( .A1(A[4]), .A2(n95), .B1(C[4]), .B2(n94), .ZN(n30) );
  AOI211_X1 U24 ( .C1(E[5]), .C2(n3), .A(n32), .B(n4), .ZN(n33) );
  INV_X1 U25 ( .A(n9), .ZN(n95) );
  INV_X1 U26 ( .A(n22), .ZN(n94) );
  INV_X1 U27 ( .A(n22), .ZN(n6) );
  INV_X1 U28 ( .A(n2), .ZN(n40) );
  INV_X1 U29 ( .A(n2), .ZN(n45) );
  INV_X1 U30 ( .A(n2), .ZN(n50) );
  INV_X1 U31 ( .A(n2), .ZN(n55) );
  INV_X1 U32 ( .A(n2), .ZN(n60) );
  INV_X1 U33 ( .A(n2), .ZN(n65) );
  INV_X1 U34 ( .A(n2), .ZN(n70) );
  INV_X1 U35 ( .A(n2), .ZN(n84) );
  INV_X1 U36 ( .A(n2), .ZN(n79) );
  INV_X1 U37 ( .A(SEL[0]), .ZN(n8) );
  NOR2_X1 U38 ( .A1(n2), .A2(n31), .ZN(n32) );
  AND2_X1 U39 ( .A1(B[5]), .A2(n92), .ZN(n4) );
  AND2_X1 U40 ( .A1(SEL[2]), .A2(SEL[1]), .ZN(n5) );
  AOI22_X1 U41 ( .A1(C[0]), .A2(n6), .B1(A[0]), .B2(n1), .ZN(n15) );
  AOI22_X1 U42 ( .A1(E[0]), .A2(n93), .B1(B[0]), .B2(n92), .ZN(n13) );
  AOI22_X1 U43 ( .A1(C[1]), .A2(n6), .B1(A[1]), .B2(n1), .ZN(n18) );
  AOI22_X1 U44 ( .A1(D[15]), .A2(n79), .B1(B[15]), .B2(n92), .ZN(n83) );
  AOI22_X1 U45 ( .A1(E[4]), .A2(n3), .B1(B[4]), .B2(n92), .ZN(n28) );
  AOI22_X1 U46 ( .A1(C[2]), .A2(n6), .B1(A[2]), .B2(n95), .ZN(n21) );
  NAND4_X1 U47 ( .A1(n44), .A2(n43), .A3(n42), .A4(n41), .ZN(Y[7]) );
  AOI22_X1 U48 ( .A1(D[7]), .A2(n40), .B1(B[7]), .B2(n92), .ZN(n44) );
  NAND4_X1 U49 ( .A1(n49), .A2(n48), .A3(n47), .A4(n46), .ZN(Y[8]) );
  AOI22_X1 U50 ( .A1(D[8]), .A2(n45), .B1(B[8]), .B2(n92), .ZN(n49) );
  NAND4_X1 U51 ( .A1(n54), .A2(n53), .A3(n52), .A4(n51), .ZN(Y[9]) );
  AOI22_X1 U52 ( .A1(D[9]), .A2(n50), .B1(B[9]), .B2(n92), .ZN(n54) );
  AOI22_X1 U53 ( .A1(D[10]), .A2(n55), .B1(B[10]), .B2(n92), .ZN(n59) );
  AOI22_X1 U54 ( .A1(D[11]), .A2(n60), .B1(B[11]), .B2(n92), .ZN(n64) );
  NAND4_X1 U55 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(Y[12]) );
  AOI22_X1 U56 ( .A1(D[12]), .A2(n65), .B1(B[12]), .B2(n92), .ZN(n69) );
  AOI22_X1 U57 ( .A1(D[13]), .A2(n70), .B1(B[13]), .B2(n92), .ZN(n74) );
  AOI22_X1 U58 ( .A1(D[14]), .A2(n79), .B1(B[14]), .B2(n92), .ZN(n78) );
  NAND4_X1 U59 ( .A1(n39), .A2(n38), .A3(n37), .A4(n36), .ZN(Y[6]) );
  AOI22_X1 U60 ( .A1(D[6]), .A2(n40), .B1(B[6]), .B2(n92), .ZN(n39) );
  AOI22_X1 U61 ( .A1(D[18]), .A2(n84), .B1(B[18]), .B2(n92), .ZN(n98) );
  AOI22_X1 U62 ( .A1(A[18]), .A2(n95), .B1(C[18]), .B2(n94), .ZN(n96) );
  AOI22_X1 U63 ( .A1(D[17]), .A2(n84), .B1(B[17]), .B2(n92), .ZN(n90) );
  AOI22_X1 U64 ( .A1(A[17]), .A2(n95), .B1(C[17]), .B2(n94), .ZN(n88) );
  AOI22_X1 U65 ( .A1(D[16]), .A2(n84), .B1(B[16]), .B2(n92), .ZN(n87) );
  AOI22_X1 U66 ( .A1(A[16]), .A2(n95), .B1(C[16]), .B2(n94), .ZN(n85) );
  NAND3_X1 U67 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n7), .ZN(n22) );
  NAND2_X1 U68 ( .A1(SEL[0]), .A2(n5), .ZN(n9) );
  INV_X1 U69 ( .A(n2), .ZN(n27) );
  NAND2_X1 U70 ( .A1(D[0]), .A2(n27), .ZN(n14) );
  NAND2_X1 U71 ( .A1(n9), .A2(n22), .ZN(n11) );
  NAND2_X1 U72 ( .A1(n8), .A2(n5), .ZN(n12) );
  NAND2_X1 U73 ( .A1(n12), .A2(n91), .ZN(n10) );
  NAND3_X1 U74 ( .A1(n15), .A2(n14), .A3(n13), .ZN(Y[0]) );
  NAND2_X1 U75 ( .A1(D[1]), .A2(n27), .ZN(n17) );
  NAND2_X1 U76 ( .A1(D[2]), .A2(n27), .ZN(n20) );
  NAND3_X1 U77 ( .A1(n21), .A2(n20), .A3(n19), .ZN(Y[2]) );
  NAND2_X1 U78 ( .A1(E[3]), .A2(n3), .ZN(n26) );
  NAND2_X1 U79 ( .A1(B[3]), .A2(n92), .ZN(n25) );
  NAND2_X1 U80 ( .A1(D[3]), .A2(n27), .ZN(n24) );
  AOI22_X1 U81 ( .A1(C[3]), .A2(n94), .B1(A[3]), .B2(n95), .ZN(n23) );
  NAND4_X1 U82 ( .A1(n26), .A2(n25), .A3(n24), .A4(n23), .ZN(Y[3]) );
  NAND2_X1 U83 ( .A1(D[4]), .A2(n27), .ZN(n29) );
  NAND3_X1 U84 ( .A1(n30), .A2(n29), .A3(n28), .ZN(Y[4]) );
  NAND2_X1 U85 ( .A1(A[5]), .A2(n95), .ZN(n35) );
  NAND2_X1 U86 ( .A1(C[5]), .A2(n94), .ZN(n34) );
  INV_X1 U87 ( .A(D[5]), .ZN(n31) );
  NAND3_X1 U88 ( .A1(n35), .A2(n34), .A3(n33), .ZN(Y[5]) );
  NAND2_X1 U89 ( .A1(E[6]), .A2(n3), .ZN(n38) );
  NAND2_X1 U90 ( .A1(A[6]), .A2(n95), .ZN(n36) );
  NAND2_X1 U91 ( .A1(E[7]), .A2(n3), .ZN(n43) );
  NAND2_X1 U92 ( .A1(C[7]), .A2(n94), .ZN(n42) );
  NAND2_X1 U93 ( .A1(A[7]), .A2(n95), .ZN(n41) );
  NAND2_X1 U94 ( .A1(E[8]), .A2(n3), .ZN(n48) );
  NAND2_X1 U95 ( .A1(C[8]), .A2(n94), .ZN(n47) );
  NAND2_X1 U96 ( .A1(A[8]), .A2(n95), .ZN(n46) );
  NAND2_X1 U97 ( .A1(E[9]), .A2(n3), .ZN(n53) );
  NAND2_X1 U98 ( .A1(A[9]), .A2(n95), .ZN(n51) );
  NAND2_X1 U99 ( .A1(E[10]), .A2(n3), .ZN(n58) );
  NAND2_X1 U100 ( .A1(A[10]), .A2(n95), .ZN(n56) );
  NAND2_X1 U101 ( .A1(E[11]), .A2(n3), .ZN(n63) );
  NAND2_X1 U102 ( .A1(A[11]), .A2(n95), .ZN(n61) );
  NAND2_X1 U103 ( .A1(E[12]), .A2(n3), .ZN(n68) );
  NAND2_X1 U104 ( .A1(C[12]), .A2(n94), .ZN(n67) );
  NAND2_X1 U105 ( .A1(A[12]), .A2(n95), .ZN(n66) );
  NAND2_X1 U106 ( .A1(E[13]), .A2(n3), .ZN(n73) );
  NAND2_X1 U107 ( .A1(A[13]), .A2(n95), .ZN(n71) );
  NAND2_X1 U108 ( .A1(E[14]), .A2(n3), .ZN(n77) );
  NAND2_X1 U109 ( .A1(A[14]), .A2(n95), .ZN(n75) );
  NAND2_X1 U110 ( .A1(E[15]), .A2(n3), .ZN(n82) );
  NAND2_X1 U111 ( .A1(A[15]), .A2(n95), .ZN(n80) );
  NAND2_X1 U112 ( .A1(E[16]), .A2(n3), .ZN(n86) );
  NAND3_X1 U113 ( .A1(n87), .A2(n86), .A3(n85), .ZN(Y[16]) );
  NAND2_X1 U114 ( .A1(E[17]), .A2(n3), .ZN(n89) );
  NAND3_X1 U115 ( .A1(n90), .A2(n89), .A3(n88), .ZN(Y[17]) );
  NAND2_X1 U116 ( .A1(E[18]), .A2(n3), .ZN(n97) );
  NAND3_X1 U117 ( .A1(n98), .A2(n97), .A3(n96), .ZN(Y[18]) );
endmodule


module PG_BLOCK_0 ( Gi_0, Gi_1, Pi_0, Pi_1, Po, Go );
  input Gi_0, Gi_1, Pi_0, Pi_1;
  output Po, Go;


  GENERAL_GENERATE_27 GEN_BLOCK ( .Gi_0(Gi_0), .Gi_1(Gi_1), .Pi(Pi_1), .Go(Go)
         );
  GENERAL_PROPAGATE_0 PRO_BLOCK ( .Pi({Pi_1, Pi_0}), .Po(Po) );
endmodule


module GENERAL_GENERATE_0 ( Gi_0, Gi_1, Pi, Go );
  input Gi_0, Gi_1, Pi;
  output Go;
  wire   OUT_AND;

  AND_GATE_1_482 AND_INST ( .A(Pi), .B(Gi_0), .Y(OUT_AND) );
  OR_GATE_242 OR_INST ( .A(Gi_1), .B(OUT_AND), .Y(Go) );
endmodule


module PG_NETWORK_N32 ( A, B, Ci, G, P );
  input [31:0] A;
  input [31:0] B;
  output [31:0] G;
  output [31:0] P;
  input Ci;
  wire   G_tmp, P_tmp;
  assign P[0] = 1'b0;

  AND_GATE_1_514 FIRST_GEN_BLOCK ( .A(A[0]), .B(B[0]), .Y(G_tmp) );
  XOR_GATE_1_450 FIRST_PRO_BLOCK ( .A(A[0]), .B(B[0]), .Y(P_tmp) );
  GENERAL_GENERATE_28 FIRST_GENERATE ( .Gi_0(Ci), .Gi_1(G_tmp), .Pi(P_tmp), 
        .Go(G[0]) );
  AND_GATE_1_513 GEN_BLOCK_1 ( .A(A[1]), .B(B[1]), .Y(G[1]) );
  XOR_GATE_1_449 PRO_BLOCK_1 ( .A(A[1]), .B(B[1]), .Y(P[1]) );
  AND_GATE_1_512 GEN_BLOCK_2 ( .A(A[2]), .B(B[2]), .Y(G[2]) );
  XOR_GATE_1_448 PRO_BLOCK_2 ( .A(A[2]), .B(B[2]), .Y(P[2]) );
  AND_GATE_1_511 GEN_BLOCK_3 ( .A(A[3]), .B(B[3]), .Y(G[3]) );
  XOR_GATE_1_447 PRO_BLOCK_3 ( .A(A[3]), .B(B[3]), .Y(P[3]) );
  AND_GATE_1_510 GEN_BLOCK_4 ( .A(A[4]), .B(B[4]), .Y(G[4]) );
  XOR_GATE_1_446 PRO_BLOCK_4 ( .A(A[4]), .B(B[4]), .Y(P[4]) );
  AND_GATE_1_509 GEN_BLOCK_5 ( .A(A[5]), .B(B[5]), .Y(G[5]) );
  XOR_GATE_1_445 PRO_BLOCK_5 ( .A(A[5]), .B(B[5]), .Y(P[5]) );
  AND_GATE_1_508 GEN_BLOCK_6 ( .A(A[6]), .B(B[6]), .Y(G[6]) );
  XOR_GATE_1_444 PRO_BLOCK_6 ( .A(A[6]), .B(B[6]), .Y(P[6]) );
  AND_GATE_1_507 GEN_BLOCK_7 ( .A(A[7]), .B(B[7]), .Y(G[7]) );
  XOR_GATE_1_443 PRO_BLOCK_7 ( .A(A[7]), .B(B[7]), .Y(P[7]) );
  AND_GATE_1_506 GEN_BLOCK_8 ( .A(A[8]), .B(B[8]), .Y(G[8]) );
  XOR_GATE_1_442 PRO_BLOCK_8 ( .A(A[8]), .B(B[8]), .Y(P[8]) );
  AND_GATE_1_505 GEN_BLOCK_9 ( .A(A[9]), .B(B[9]), .Y(G[9]) );
  XOR_GATE_1_441 PRO_BLOCK_9 ( .A(A[9]), .B(B[9]), .Y(P[9]) );
  AND_GATE_1_504 GEN_BLOCK_10 ( .A(A[10]), .B(B[10]), .Y(G[10]) );
  XOR_GATE_1_440 PRO_BLOCK_10 ( .A(A[10]), .B(B[10]), .Y(P[10]) );
  AND_GATE_1_503 GEN_BLOCK_11 ( .A(A[11]), .B(B[11]), .Y(G[11]) );
  XOR_GATE_1_439 PRO_BLOCK_11 ( .A(A[11]), .B(B[11]), .Y(P[11]) );
  AND_GATE_1_502 GEN_BLOCK_12 ( .A(A[12]), .B(B[12]), .Y(G[12]) );
  XOR_GATE_1_438 PRO_BLOCK_12 ( .A(A[12]), .B(B[12]), .Y(P[12]) );
  AND_GATE_1_501 GEN_BLOCK_13 ( .A(A[13]), .B(B[13]), .Y(G[13]) );
  XOR_GATE_1_437 PRO_BLOCK_13 ( .A(A[13]), .B(B[13]), .Y(P[13]) );
  AND_GATE_1_500 GEN_BLOCK_14 ( .A(A[14]), .B(B[14]), .Y(G[14]) );
  XOR_GATE_1_436 PRO_BLOCK_14 ( .A(A[14]), .B(B[14]), .Y(P[14]) );
  AND_GATE_1_499 GEN_BLOCK_15 ( .A(A[15]), .B(B[15]), .Y(G[15]) );
  XOR_GATE_1_435 PRO_BLOCK_15 ( .A(A[15]), .B(B[15]), .Y(P[15]) );
  AND_GATE_1_498 GEN_BLOCK_16 ( .A(A[16]), .B(B[16]), .Y(G[16]) );
  XOR_GATE_1_434 PRO_BLOCK_16 ( .A(A[16]), .B(B[16]), .Y(P[16]) );
  AND_GATE_1_497 GEN_BLOCK_17 ( .A(A[17]), .B(B[17]), .Y(G[17]) );
  XOR_GATE_1_433 PRO_BLOCK_17 ( .A(A[17]), .B(B[17]), .Y(P[17]) );
  AND_GATE_1_496 GEN_BLOCK_18 ( .A(A[18]), .B(B[18]), .Y(G[18]) );
  XOR_GATE_1_432 PRO_BLOCK_18 ( .A(A[18]), .B(B[18]), .Y(P[18]) );
  AND_GATE_1_495 GEN_BLOCK_19 ( .A(A[19]), .B(B[19]), .Y(G[19]) );
  XOR_GATE_1_431 PRO_BLOCK_19 ( .A(A[19]), .B(B[19]), .Y(P[19]) );
  AND_GATE_1_494 GEN_BLOCK_20 ( .A(A[20]), .B(B[20]), .Y(G[20]) );
  XOR_GATE_1_430 PRO_BLOCK_20 ( .A(A[20]), .B(B[20]), .Y(P[20]) );
  AND_GATE_1_493 GEN_BLOCK_21 ( .A(A[21]), .B(B[21]), .Y(G[21]) );
  XOR_GATE_1_429 PRO_BLOCK_21 ( .A(A[21]), .B(B[21]), .Y(P[21]) );
  AND_GATE_1_492 GEN_BLOCK_22 ( .A(A[22]), .B(B[22]), .Y(G[22]) );
  XOR_GATE_1_428 PRO_BLOCK_22 ( .A(A[22]), .B(B[22]), .Y(P[22]) );
  AND_GATE_1_491 GEN_BLOCK_23 ( .A(A[23]), .B(B[23]), .Y(G[23]) );
  XOR_GATE_1_427 PRO_BLOCK_23 ( .A(A[23]), .B(B[23]), .Y(P[23]) );
  AND_GATE_1_490 GEN_BLOCK_24 ( .A(A[24]), .B(B[24]), .Y(G[24]) );
  XOR_GATE_1_426 PRO_BLOCK_24 ( .A(A[24]), .B(B[24]), .Y(P[24]) );
  AND_GATE_1_489 GEN_BLOCK_25 ( .A(A[25]), .B(B[25]), .Y(G[25]) );
  XOR_GATE_1_425 PRO_BLOCK_25 ( .A(A[25]), .B(B[25]), .Y(P[25]) );
  AND_GATE_1_488 GEN_BLOCK_26 ( .A(A[26]), .B(B[26]), .Y(G[26]) );
  XOR_GATE_1_424 PRO_BLOCK_26 ( .A(A[26]), .B(B[26]), .Y(P[26]) );
  AND_GATE_1_487 GEN_BLOCK_27 ( .A(A[27]), .B(B[27]), .Y(G[27]) );
  XOR_GATE_1_423 PRO_BLOCK_27 ( .A(A[27]), .B(B[27]), .Y(P[27]) );
  AND_GATE_1_486 GEN_BLOCK_28 ( .A(A[28]), .B(B[28]), .Y(G[28]) );
  XOR_GATE_1_422 PRO_BLOCK_28 ( .A(A[28]), .B(B[28]), .Y(P[28]) );
  AND_GATE_1_485 GEN_BLOCK_29 ( .A(A[29]), .B(B[29]), .Y(G[29]) );
  XOR_GATE_1_421 PRO_BLOCK_29 ( .A(A[29]), .B(B[29]), .Y(P[29]) );
  AND_GATE_1_484 GEN_BLOCK_30 ( .A(A[30]), .B(B[30]), .Y(G[30]) );
  XOR_GATE_1_420 PRO_BLOCK_30 ( .A(A[30]), .B(B[30]), .Y(P[30]) );
  AND_GATE_1_483 GEN_BLOCK_31 ( .A(A[31]), .B(B[31]), .Y(G[31]) );
  XOR_GATE_1_419 PRO_BLOCK_31 ( .A(A[31]), .B(B[31]), .Y(P[31]) );
endmodule


module FSM_DIVISOR ( CLK, RST, EN, SEL_R_MUX_IN, SEL_Q_MUX_IN, SEL_D_MUX, 
        SEL_ADD_IN_D_MUX, SEL_ADD_IN_R_MUX, SEL_SIGN_MUX, EN_D, EN_Z, EN_Q, 
        EN_R, EN_SIGN, MSB_REM );
  output [1:0] SEL_ADD_IN_D_MUX;
  output [1:0] SEL_ADD_IN_R_MUX;
  output [1:0] SEL_SIGN_MUX;
  input CLK, RST, EN, MSB_REM;
  output SEL_R_MUX_IN, SEL_Q_MUX_IN, SEL_D_MUX, EN_D, EN_Z, EN_Q, EN_R,
         EN_SIGN;
  wire   \CURRENT_STATE[3] , N27, N28, N29, N30, N31, N32, N33, N34, N35, N36,
         N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N60, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n54,
         n55, n56, n57, n58, n61, n62, n63, n64, n65, n66, n67, n68, n69, n71,
         n72, n73, n74, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n144, n145, n146, n147, n1, n2, n3, n4, n5,
         n53, n59, n60, n70, n75, n76, SEL_D_MUX, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89;
  wire   [31:0] CNT;
  assign EN_Z = SEL_D_MUX;
  assign EN_SIGN = SEL_D_MUX;

  DFFR_X1 \CURRENT_STATE_reg[0]  ( .D(n144), .CK(CLK), .RN(n78), .Q(n1), .QN(
        n145) );
  DFFR_X1 \CURRENT_STATE_reg[3]  ( .D(n142), .CK(CLK), .RN(n78), .Q(
        \CURRENT_STATE[3] ), .QN(n2) );
  DFFR_X1 \CURRENT_STATE_reg[1]  ( .D(n141), .CK(CLK), .RN(n78), .QN(n146) );
  DFF_X1 \CNT_reg[19]  ( .D(n140), .CK(CLK), .Q(CNT[19]) );
  DFF_X1 \CNT_reg[0]  ( .D(n139), .CK(CLK), .Q(CNT[0]) );
  DFF_X1 \CNT_reg[1]  ( .D(n138), .CK(CLK), .Q(CNT[1]) );
  DFF_X1 \CNT_reg[2]  ( .D(n137), .CK(CLK), .Q(CNT[2]) );
  DFF_X1 \CNT_reg[3]  ( .D(n136), .CK(CLK), .Q(CNT[3]) );
  DFF_X1 \CNT_reg[4]  ( .D(n135), .CK(CLK), .Q(CNT[4]) );
  DFF_X1 \CNT_reg[5]  ( .D(n134), .CK(CLK), .Q(CNT[5]) );
  DFF_X1 \CNT_reg[6]  ( .D(n133), .CK(CLK), .Q(CNT[6]) );
  DFF_X1 \CNT_reg[7]  ( .D(n132), .CK(CLK), .Q(CNT[7]) );
  DFF_X1 \CNT_reg[8]  ( .D(n131), .CK(CLK), .Q(CNT[8]) );
  DFF_X1 \CNT_reg[9]  ( .D(n130), .CK(CLK), .Q(CNT[9]) );
  DFF_X1 \CNT_reg[10]  ( .D(n129), .CK(CLK), .Q(CNT[10]) );
  DFF_X1 \CNT_reg[11]  ( .D(n128), .CK(CLK), .Q(CNT[11]) );
  DFF_X1 \CNT_reg[12]  ( .D(n127), .CK(CLK), .Q(CNT[12]) );
  DFF_X1 \CNT_reg[13]  ( .D(n126), .CK(CLK), .Q(CNT[13]) );
  DFF_X1 \CNT_reg[14]  ( .D(n125), .CK(CLK), .Q(CNT[14]) );
  DFF_X1 \CNT_reg[15]  ( .D(n124), .CK(CLK), .Q(CNT[15]) );
  DFF_X1 \CNT_reg[16]  ( .D(n123), .CK(CLK), .Q(CNT[16]) );
  DFF_X1 \CNT_reg[17]  ( .D(n122), .CK(CLK), .Q(CNT[17]) );
  DFF_X1 \CNT_reg[18]  ( .D(n121), .CK(CLK), .Q(CNT[18]) );
  DFF_X1 \CNT_reg[20]  ( .D(n120), .CK(CLK), .Q(CNT[20]) );
  DFF_X1 \CNT_reg[21]  ( .D(n119), .CK(CLK), .Q(CNT[21]) );
  DFF_X1 \CNT_reg[22]  ( .D(n118), .CK(CLK), .Q(CNT[22]) );
  DFF_X1 \CNT_reg[23]  ( .D(n117), .CK(CLK), .Q(CNT[23]) );
  DFF_X1 \CNT_reg[24]  ( .D(n116), .CK(CLK), .Q(CNT[24]) );
  DFF_X1 \CNT_reg[25]  ( .D(n115), .CK(CLK), .Q(CNT[25]) );
  DFF_X1 \CNT_reg[26]  ( .D(n114), .CK(CLK), .Q(CNT[26]) );
  DFF_X1 \CNT_reg[27]  ( .D(n113), .CK(CLK), .Q(CNT[27]) );
  DFF_X1 \CNT_reg[28]  ( .D(n112), .CK(CLK), .Q(CNT[28]) );
  DFF_X1 \CNT_reg[29]  ( .D(n111), .CK(CLK), .Q(CNT[29]) );
  DFF_X1 \CNT_reg[30]  ( .D(n110), .CK(CLK), .Q(CNT[30]) );
  DFF_X1 \CNT_reg[31]  ( .D(n109), .CK(CLK), .Q(CNT[31]), .QN(n4) );
  DFFR_X1 \CURRENT_STATE_reg[2]  ( .D(n108), .CK(CLK), .RN(n78), .Q(n3), .QN(
        n147) );
  NAND2_X1 U83 ( .A1(n50), .A2(n3), .ZN(n58) );
  NAND2_X1 U87 ( .A1(n62), .A2(n51), .ZN(SEL_SIGN_MUX[1]) );
  NAND3_X1 U90 ( .A1(n54), .A2(n64), .A3(n65), .ZN(SEL_ADD_IN_R_MUX[1]) );
  NAND2_X1 U92 ( .A1(n47), .A2(n68), .ZN(SEL_ADD_IN_R_MUX[0]) );
  NAND2_X1 U94 ( .A1(n69), .A2(n64), .ZN(SEL_Q_MUX_IN) );
  NAND2_X1 U95 ( .A1(n69), .A2(n5), .ZN(SEL_ADD_IN_D_MUX[1]) );
  NAND2_X1 U97 ( .A1(n52), .A2(n63), .ZN(SEL_ADD_IN_D_MUX[0]) );
  NAND3_X1 U99 ( .A1(n54), .A2(n64), .A3(n62), .ZN(EN_R) );
  NAND2_X1 U101 ( .A1(n72), .A2(n47), .ZN(n71) );
  NAND2_X1 U102 ( .A1(n49), .A2(n73), .ZN(n47) );
  NAND3_X1 U104 ( .A1(n52), .A2(n64), .A3(n72), .ZN(EN_Q) );
  NAND3_X1 U107 ( .A1(n73), .A2(n1), .A3(n147), .ZN(n9) );
  NAND2_X1 U112 ( .A1(n66), .A2(n73), .ZN(n52) );
  NAND2_X1 U114 ( .A1(n74), .A2(n5), .ZN(EN_D) );
  NAND2_X1 U117 ( .A1(n146), .A2(n2), .ZN(n51) );
  NAND3_X1 U121 ( .A1(n147), .A2(n73), .A3(n145), .ZN(n74) );
  FSM_DIVISOR_DW01_inc_0 add_63 ( .A(CNT), .SUM({N58, N57, N56, N55, N54, N53, 
        N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, 
        N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27}) );
  INV_X1 U3 ( .A(MSB_REM), .ZN(n50) );
  INV_X1 U4 ( .A(n71), .ZN(n62) );
  INV_X1 U5 ( .A(n63), .ZN(SEL_SIGN_MUX[0]) );
  INV_X1 U6 ( .A(n67), .ZN(n72) );
  BUF_X1 U7 ( .A(n12), .Z(n76) );
  BUF_X1 U8 ( .A(n12), .Z(n70) );
  BUF_X1 U9 ( .A(n12), .Z(n75) );
  AOI211_X1 U10 ( .C1(n61), .C2(n66), .A(EN_D), .B(n71), .ZN(n63) );
  AOI21_X1 U11 ( .B1(n66), .B2(n2), .A(n67), .ZN(n65) );
  OAI21_X1 U12 ( .B1(n7), .B2(n51), .A(n9), .ZN(n67) );
  INV_X1 U13 ( .A(n51), .ZN(n61) );
  OR3_X1 U14 ( .A1(n1), .A2(n3), .A3(n51), .ZN(n5) );
  INV_X1 U15 ( .A(n49), .ZN(n7) );
  AND2_X1 U16 ( .A1(n54), .A2(n52), .ZN(n69) );
  NOR2_X1 U17 ( .A1(n60), .A2(n9), .ZN(n12) );
  INV_X1 U18 ( .A(n64), .ZN(SEL_R_MUX_IN) );
  NOR2_X1 U19 ( .A1(n10), .A2(n61), .ZN(n6) );
  BUF_X1 U20 ( .A(n13), .Z(n60) );
  BUF_X1 U21 ( .A(n13), .Z(n53) );
  BUF_X1 U22 ( .A(n13), .Z(n59) );
  NOR2_X1 U23 ( .A1(n57), .A2(n9), .ZN(n45) );
  INV_X1 U24 ( .A(N60), .ZN(n57) );
  AOI21_X1 U25 ( .B1(n147), .B2(n61), .A(EN_D), .ZN(n64) );
  INV_X1 U26 ( .A(n11), .ZN(n109) );
  AOI22_X1 U27 ( .A1(N58), .A2(n70), .B1(CNT[31]), .B2(n53), .ZN(n11) );
  NOR2_X1 U28 ( .A1(n145), .A2(n147), .ZN(n66) );
  NAND4_X1 U29 ( .A1(\CURRENT_STATE[3] ), .A2(n145), .A3(n146), .A4(n147), 
        .ZN(n54) );
  NOR2_X1 U30 ( .A1(n1), .A2(n147), .ZN(n49) );
  INV_X1 U31 ( .A(n21), .ZN(n117) );
  AOI22_X1 U32 ( .A1(N50), .A2(n70), .B1(CNT[23]), .B2(n53), .ZN(n21) );
  NOR2_X1 U33 ( .A1(\CURRENT_STATE[3] ), .A2(n146), .ZN(n73) );
  OAI211_X1 U34 ( .C1(n146), .C2(EN), .A(n46), .B(n47), .ZN(n141) );
  OAI21_X1 U35 ( .B1(n48), .B2(n45), .A(EN), .ZN(n46) );
  AOI21_X1 U36 ( .B1(n49), .B2(n50), .A(n51), .ZN(n48) );
  OAI21_X1 U37 ( .B1(n145), .B2(n6), .A(n55), .ZN(n144) );
  OAI21_X1 U38 ( .B1(n56), .B2(n45), .A(EN), .ZN(n55) );
  AOI211_X1 U39 ( .C1(n146), .C2(n58), .A(n1), .B(\CURRENT_STATE[3] ), .ZN(n56) );
  INV_X1 U40 ( .A(n14), .ZN(n110) );
  AOI22_X1 U41 ( .A1(N57), .A2(n70), .B1(CNT[30]), .B2(n53), .ZN(n14) );
  INV_X1 U42 ( .A(n15), .ZN(n111) );
  AOI22_X1 U43 ( .A1(N56), .A2(n70), .B1(CNT[29]), .B2(n53), .ZN(n15) );
  INV_X1 U44 ( .A(n16), .ZN(n112) );
  AOI22_X1 U45 ( .A1(N55), .A2(n70), .B1(CNT[28]), .B2(n53), .ZN(n16) );
  INV_X1 U46 ( .A(n19), .ZN(n115) );
  AOI22_X1 U47 ( .A1(N52), .A2(n70), .B1(CNT[25]), .B2(n53), .ZN(n19) );
  INV_X1 U48 ( .A(n17), .ZN(n113) );
  AOI22_X1 U49 ( .A1(N54), .A2(n70), .B1(CNT[27]), .B2(n53), .ZN(n17) );
  INV_X1 U50 ( .A(n20), .ZN(n116) );
  AOI22_X1 U51 ( .A1(N51), .A2(n70), .B1(CNT[24]), .B2(n53), .ZN(n20) );
  INV_X1 U52 ( .A(n18), .ZN(n114) );
  AOI22_X1 U53 ( .A1(N53), .A2(n70), .B1(CNT[26]), .B2(n53), .ZN(n18) );
  OAI211_X1 U54 ( .C1(n45), .C2(SEL_D_MUX), .A(n78), .B(EN), .ZN(n13) );
  OAI221_X1 U55 ( .B1(n147), .B2(n6), .C1(\CURRENT_STATE[3] ), .C2(n7), .A(n8), 
        .ZN(n108) );
  OR3_X1 U56 ( .A1(n9), .A2(N60), .A3(n10), .ZN(n8) );
  OAI221_X1 U57 ( .B1(n10), .B2(n52), .C1(EN), .C2(n2), .A(n54), .ZN(n142) );
  INV_X1 U58 ( .A(n22), .ZN(n118) );
  AOI22_X1 U59 ( .A1(N49), .A2(n70), .B1(CNT[22]), .B2(n53), .ZN(n22) );
  INV_X1 U60 ( .A(n24), .ZN(n120) );
  AOI22_X1 U61 ( .A1(N47), .A2(n70), .B1(CNT[20]), .B2(n53), .ZN(n24) );
  INV_X1 U62 ( .A(n27), .ZN(n123) );
  AOI22_X1 U63 ( .A1(N43), .A2(n75), .B1(CNT[16]), .B2(n59), .ZN(n27) );
  INV_X1 U64 ( .A(n30), .ZN(n126) );
  AOI22_X1 U65 ( .A1(N40), .A2(n75), .B1(CNT[13]), .B2(n59), .ZN(n30) );
  INV_X1 U66 ( .A(n43), .ZN(n139) );
  AOI22_X1 U67 ( .A1(N27), .A2(n76), .B1(CNT[0]), .B2(n60), .ZN(n43) );
  INV_X1 U68 ( .A(n28), .ZN(n124) );
  AOI22_X1 U69 ( .A1(N42), .A2(n75), .B1(CNT[15]), .B2(n59), .ZN(n28) );
  INV_X1 U70 ( .A(n34), .ZN(n130) );
  AOI22_X1 U71 ( .A1(N36), .A2(n75), .B1(CNT[9]), .B2(n59), .ZN(n34) );
  INV_X1 U72 ( .A(n40), .ZN(n136) );
  AOI22_X1 U73 ( .A1(N30), .A2(n76), .B1(CNT[3]), .B2(n60), .ZN(n40) );
  INV_X1 U74 ( .A(n23), .ZN(n119) );
  AOI22_X1 U75 ( .A1(N48), .A2(n70), .B1(CNT[21]), .B2(n53), .ZN(n23) );
  INV_X1 U76 ( .A(n29), .ZN(n125) );
  AOI22_X1 U77 ( .A1(N41), .A2(n75), .B1(CNT[14]), .B2(n59), .ZN(n29) );
  INV_X1 U78 ( .A(n35), .ZN(n131) );
  AOI22_X1 U79 ( .A1(N35), .A2(n75), .B1(CNT[8]), .B2(n59), .ZN(n35) );
  INV_X1 U80 ( .A(n25), .ZN(n121) );
  AOI22_X1 U81 ( .A1(N45), .A2(n70), .B1(CNT[18]), .B2(n53), .ZN(n25) );
  INV_X1 U82 ( .A(n38), .ZN(n134) );
  AOI22_X1 U84 ( .A1(N32), .A2(n75), .B1(CNT[5]), .B2(n59), .ZN(n38) );
  INV_X1 U85 ( .A(n33), .ZN(n129) );
  AOI22_X1 U86 ( .A1(N37), .A2(n75), .B1(CNT[10]), .B2(n59), .ZN(n33) );
  INV_X1 U88 ( .A(n36), .ZN(n132) );
  AOI22_X1 U89 ( .A1(N34), .A2(n75), .B1(CNT[7]), .B2(n59), .ZN(n36) );
  INV_X1 U91 ( .A(n32), .ZN(n128) );
  AOI22_X1 U93 ( .A1(N38), .A2(n75), .B1(CNT[11]), .B2(n59), .ZN(n32) );
  INV_X1 U96 ( .A(n26), .ZN(n122) );
  AOI22_X1 U98 ( .A1(N44), .A2(n75), .B1(CNT[17]), .B2(n59), .ZN(n26) );
  INV_X1 U100 ( .A(n39), .ZN(n135) );
  AOI22_X1 U103 ( .A1(N31), .A2(n76), .B1(CNT[4]), .B2(n60), .ZN(n39) );
  INV_X1 U105 ( .A(n31), .ZN(n127) );
  AOI22_X1 U106 ( .A1(N39), .A2(n75), .B1(CNT[12]), .B2(n59), .ZN(n31) );
  INV_X1 U108 ( .A(n37), .ZN(n133) );
  AOI22_X1 U109 ( .A1(N33), .A2(n75), .B1(CNT[6]), .B2(n59), .ZN(n37) );
  INV_X1 U110 ( .A(n44), .ZN(n140) );
  AOI22_X1 U111 ( .A1(N46), .A2(n76), .B1(CNT[19]), .B2(n60), .ZN(n44) );
  INV_X1 U113 ( .A(n41), .ZN(n137) );
  AOI22_X1 U115 ( .A1(N29), .A2(n76), .B1(CNT[2]), .B2(n60), .ZN(n41) );
  INV_X1 U116 ( .A(n42), .ZN(n138) );
  AOI22_X1 U118 ( .A1(N28), .A2(n76), .B1(CNT[1]), .B2(n60), .ZN(n42) );
  INV_X1 U119 ( .A(EN), .ZN(n10) );
  INV_X1 U120 ( .A(SEL_Q_MUX_IN), .ZN(n68) );
  INV_X1 U122 ( .A(n5), .ZN(SEL_D_MUX) );
  INV_X1 U123 ( .A(RST), .ZN(n78) );
  NOR3_X1 U124 ( .A1(CNT[23]), .A2(CNT[25]), .A3(CNT[24]), .ZN(n82) );
  NOR4_X1 U125 ( .A1(CNT[29]), .A2(CNT[28]), .A3(CNT[27]), .A4(CNT[26]), .ZN(
        n81) );
  NOR3_X1 U126 ( .A1(CNT[30]), .A2(CNT[5]), .A3(CNT[4]), .ZN(n80) );
  NOR4_X1 U127 ( .A1(CNT[9]), .A2(CNT[8]), .A3(CNT[7]), .A4(CNT[6]), .ZN(n79)
         );
  NAND4_X1 U128 ( .A1(n82), .A2(n81), .A3(n80), .A4(n79), .ZN(n89) );
  AND2_X1 U129 ( .A1(CNT[2]), .A2(CNT[1]), .ZN(n83) );
  AOI211_X1 U130 ( .C1(n83), .C2(CNT[3]), .A(CNT[11]), .B(CNT[10]), .ZN(n87)
         );
  NOR4_X1 U131 ( .A1(CNT[15]), .A2(CNT[14]), .A3(CNT[13]), .A4(CNT[12]), .ZN(
        n86) );
  NOR3_X1 U132 ( .A1(CNT[16]), .A2(CNT[18]), .A3(CNT[17]), .ZN(n85) );
  NOR4_X1 U133 ( .A1(CNT[22]), .A2(CNT[21]), .A3(CNT[20]), .A4(CNT[19]), .ZN(
        n84) );
  NAND4_X1 U134 ( .A1(n87), .A2(n86), .A3(n85), .A4(n84), .ZN(n88) );
  OAI21_X1 U135 ( .B1(n89), .B2(n88), .A(n4), .ZN(N60) );
endmodule


module NR_DIVISOR_DATAPATH ( CLK, RST, Z, D, Q, R, MSB_REM, ADD_IN_D, ADD_IN_R, 
        SIGN, ADD_OUT, SEL_R_MUX_IN, SEL_Q_MUX_IN, SEL_D_MUX, SEL_ADD_IN_D_MUX, 
        SEL_ADD_IN_R_MUX, SEL_SIGN_MUX, EN_D, EN_Z, EN_Q, EN_R, EN_SIGN );
  input [15:0] Z;
  input [15:0] D;
  output [15:0] Q;
  output [15:0] R;
  output [15:0] ADD_IN_D;
  output [15:0] ADD_IN_R;
  input [15:0] ADD_OUT;
  input [1:0] SEL_ADD_IN_D_MUX;
  input [1:0] SEL_ADD_IN_R_MUX;
  input [1:0] SEL_SIGN_MUX;
  input CLK, RST, SEL_R_MUX_IN, SEL_Q_MUX_IN, SEL_D_MUX, EN_D, EN_Z, EN_Q,
         EN_R, EN_SIGN;
  output MSB_REM, SIGN;
  wire   \Q_MUX_IN[0] , XOR_SIGN, SIGN_REG_OUT, SIGN_SIG, n1;
  wire   [15:0] R_MUX_OUT;
  wire   [15:0] Q_MUX_OUT;
  wire   [15:0] D_MUX_OUT;
  wire   [15:0] D_REG_OUT;
  wire   [15:0] Z_REG_OUT;
  assign MSB_REM = ADD_OUT[15];

  MUX21_GEN_N16_0 R_MUX_IN ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(ADD_OUT), 
        .SEL(SEL_R_MUX_IN), .Y(R_MUX_OUT) );
  REG_N16_1_0 REG_R ( .D(R_MUX_OUT), .Q(R), .EN(EN_R), .RST(n1), .CLK(CLK) );
  MUX21_GEN_N16_2 Q_MUX21_IN ( .A(ADD_OUT), .B({Q[14:0], \Q_MUX_IN[0] }), 
        .SEL(SEL_Q_MUX_IN), .Y(Q_MUX_OUT) );
  REG_N16_1_3 REG_Q ( .D(Q_MUX_OUT), .Q(Q), .EN(EN_Q), .RST(n1), .CLK(CLK) );
  MUX21_GEN_N16_1 D_MUX ( .A(D), .B(ADD_OUT), .SEL(SEL_D_MUX), .Y(D_MUX_OUT)
         );
  REG_N16_1_2 REG_D ( .D(D_MUX_OUT), .Q(D_REG_OUT), .EN(EN_D), .RST(1'b0), 
        .CLK(CLK) );
  REG_N16_1_1 REG_Z ( .D(Z), .Q(Z_REG_OUT), .EN(EN_Z), .RST(n1), .CLK(CLK) );
  MUX41_GEN_N16_0 ADD_IN_D_MUX ( .A(Q), .B(R), .C(D_REG_OUT), .D(Z_REG_OUT), 
        .SEL(SEL_ADD_IN_D_MUX), .Y(ADD_IN_D) );
  MUX41_GEN_N16_1 ADD_IN_R_MUX ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({R[14:0], 
        Q[15]}), .C(R), .D({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL(
        SEL_ADD_IN_R_MUX), .Y(ADD_IN_R) );
  XOR_GATE_1_451 SIGN_XOR ( .A(Z[15]), .B(D[15]), .Y(XOR_SIGN) );
  FD_1_65 SIGN_FD ( .D(XOR_SIGN), .CLK(CLK), .EN(EN_SIGN), .RST(n1), .Q(
        SIGN_REG_OUT) );
  MUX41_1 ADD_IN_SIGN_MUX ( .A(SIGN_SIG), .B(Z[15]), .C(D[15]), .D(
        SIGN_REG_OUT), .SEL(SEL_SIGN_MUX), .Y(SIGN) );
  INV_X1 U2 ( .A(ADD_OUT[15]), .ZN(\Q_MUX_IN[0] ) );
  INV_X1 U3 ( .A(R[15]), .ZN(SIGN_SIG) );
  BUF_X1 U4 ( .A(RST), .Z(n1) );
endmodule


module BOOTHMUL_COMP_3 ( PREVIOUS, A, NEG_A, B, P );
  input [16:0] PREVIOUS;
  input [15:0] A;
  input [15:0] NEG_A;
  input [15:0] B;
  output [20:0] P;
  wire   \SEL[1][2] , \SEL[1][1] , \SEL[1][0] , \SEL[0][2] , \SEL[0][1] ,
         \SEL[0][0] , \IN_B_RCA[1][18] , \IN_B_RCA[1][17] , \IN_B_RCA[1][16] ,
         \IN_B_RCA[1][15] , \IN_B_RCA[1][14] , \IN_B_RCA[1][13] ,
         \IN_B_RCA[1][12] , \IN_B_RCA[1][11] , \IN_B_RCA[1][10] ,
         \IN_B_RCA[1][9] , \IN_B_RCA[1][8] , \IN_B_RCA[1][7] ,
         \IN_B_RCA[1][6] , \IN_B_RCA[1][5] , \IN_B_RCA[1][4] ,
         \IN_B_RCA[1][3] , \IN_B_RCA[1][2] , \IN_B_RCA[1][1] ,
         \IN_B_RCA[1][0] , \IN_B_RCA[0][18] , \IN_B_RCA[0][17] ,
         \IN_B_RCA[0][16] , \IN_B_RCA[0][15] , \IN_B_RCA[0][14] ,
         \IN_B_RCA[0][13] , \IN_B_RCA[0][12] , \IN_B_RCA[0][11] ,
         \IN_B_RCA[0][10] , \IN_B_RCA[0][9] , \IN_B_RCA[0][8] ,
         \IN_B_RCA[0][7] , \IN_B_RCA[0][6] , \IN_B_RCA[0][5] ,
         \IN_B_RCA[0][4] , \IN_B_RCA[0][3] , \IN_B_RCA[0][2] ,
         \IN_B_RCA[0][1] , \IN_B_RCA[0][0] , \IN_A_RCA[1][18] ,
         \IN_A_RCA[1][15] , \IN_A_RCA[1][14] , \IN_A_RCA[1][13] ,
         \IN_A_RCA[1][12] , \IN_A_RCA[1][11] , \IN_A_RCA[1][10] ,
         \IN_A_RCA[1][9] , \IN_A_RCA[1][8] , \IN_A_RCA[1][7] ,
         \IN_A_RCA[1][6] , \IN_A_RCA[1][5] , \IN_A_RCA[1][4] ,
         \IN_A_RCA[1][3] , \IN_A_RCA[1][2] , \IN_A_RCA[1][1] ,
         \IN_A_RCA[1][0] ;

  MUX51_GEN_N19_2 MUX_INST_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({A[15], A, 1'b0, 1'b0}), .C({NEG_A[15], NEG_A, 1'b0, 1'b0}), .D({A, 1'b0, 
        1'b0, 1'b0}), .E({NEG_A, 1'b0, 1'b0, 1'b0}), .SEL({\SEL[0][2] , 
        \SEL[0][1] , \SEL[0][0] }), .Y({\IN_B_RCA[0][18] , \IN_B_RCA[0][17] , 
        \IN_B_RCA[0][16] , \IN_B_RCA[0][15] , \IN_B_RCA[0][14] , 
        \IN_B_RCA[0][13] , \IN_B_RCA[0][12] , \IN_B_RCA[0][11] , 
        \IN_B_RCA[0][10] , \IN_B_RCA[0][9] , \IN_B_RCA[0][8] , 
        \IN_B_RCA[0][7] , \IN_B_RCA[0][6] , \IN_B_RCA[0][5] , \IN_B_RCA[0][4] , 
        \IN_B_RCA[0][3] , \IN_B_RCA[0][2] , \IN_B_RCA[0][1] , \IN_B_RCA[0][0] }) );
  MUX51_GEN_N19_1 MUX_INST_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({A[15], A, 1'b0, 1'b0}), .C({NEG_A[15], NEG_A, 1'b0, 1'b0}), .D({A, 1'b0, 
        1'b0, 1'b0}), .E({NEG_A, 1'b0, 1'b0, 1'b0}), .SEL({\SEL[1][2] , 
        \SEL[1][1] , \SEL[1][0] }), .Y({\IN_B_RCA[1][18] , \IN_B_RCA[1][17] , 
        \IN_B_RCA[1][16] , \IN_B_RCA[1][15] , \IN_B_RCA[1][14] , 
        \IN_B_RCA[1][13] , \IN_B_RCA[1][12] , \IN_B_RCA[1][11] , 
        \IN_B_RCA[1][10] , \IN_B_RCA[1][9] , \IN_B_RCA[1][8] , 
        \IN_B_RCA[1][7] , \IN_B_RCA[1][6] , \IN_B_RCA[1][5] , \IN_B_RCA[1][4] , 
        \IN_B_RCA[1][3] , \IN_B_RCA[1][2] , \IN_B_RCA[1][1] , \IN_B_RCA[1][0] }) );
  RCA_GEN_NO_C_N19_2 RCA_INST_1_0 ( .A({PREVIOUS[16], PREVIOUS[16], PREVIOUS}), 
        .B({\IN_B_RCA[0][18] , \IN_B_RCA[0][17] , \IN_B_RCA[0][16] , 
        \IN_B_RCA[0][15] , \IN_B_RCA[0][14] , \IN_B_RCA[0][13] , 
        \IN_B_RCA[0][12] , \IN_B_RCA[0][11] , \IN_B_RCA[0][10] , 
        \IN_B_RCA[0][9] , \IN_B_RCA[0][8] , \IN_B_RCA[0][7] , \IN_B_RCA[0][6] , 
        \IN_B_RCA[0][5] , \IN_B_RCA[0][4] , \IN_B_RCA[0][3] , \IN_B_RCA[0][2] , 
        \IN_B_RCA[0][1] , \IN_B_RCA[0][0] }), .S({\IN_A_RCA[1][18] , 
        \IN_A_RCA[1][15] , \IN_A_RCA[1][14] , \IN_A_RCA[1][13] , 
        \IN_A_RCA[1][12] , \IN_A_RCA[1][11] , \IN_A_RCA[1][10] , 
        \IN_A_RCA[1][9] , \IN_A_RCA[1][8] , \IN_A_RCA[1][7] , \IN_A_RCA[1][6] , 
        \IN_A_RCA[1][5] , \IN_A_RCA[1][4] , \IN_A_RCA[1][3] , \IN_A_RCA[1][2] , 
        \IN_A_RCA[1][1] , \IN_A_RCA[1][0] , P[1:0]}) );
  RCA_GEN_NO_C_N19_1 RCA_INST_1_1 ( .A({\IN_A_RCA[1][18] , \IN_A_RCA[1][18] , 
        \IN_A_RCA[1][18] , \IN_A_RCA[1][15] , \IN_A_RCA[1][14] , 
        \IN_A_RCA[1][13] , \IN_A_RCA[1][12] , \IN_A_RCA[1][11] , 
        \IN_A_RCA[1][10] , \IN_A_RCA[1][9] , \IN_A_RCA[1][8] , 
        \IN_A_RCA[1][7] , \IN_A_RCA[1][6] , \IN_A_RCA[1][5] , \IN_A_RCA[1][4] , 
        \IN_A_RCA[1][3] , \IN_A_RCA[1][2] , \IN_A_RCA[1][1] , \IN_A_RCA[1][0] }), .B({\IN_B_RCA[1][18] , \IN_B_RCA[1][17] , \IN_B_RCA[1][16] , 
        \IN_B_RCA[1][15] , \IN_B_RCA[1][14] , \IN_B_RCA[1][13] , 
        \IN_B_RCA[1][12] , \IN_B_RCA[1][11] , \IN_B_RCA[1][10] , 
        \IN_B_RCA[1][9] , \IN_B_RCA[1][8] , \IN_B_RCA[1][7] , \IN_B_RCA[1][6] , 
        \IN_B_RCA[1][5] , \IN_B_RCA[1][4] , \IN_B_RCA[1][3] , \IN_B_RCA[1][2] , 
        \IN_B_RCA[1][1] , \IN_B_RCA[1][0] }), .S(P[20:2]) );
  BOOTH_ENCODER_2 ENCODERS_6 ( .TO_ENC(B[13:11]), .ENC({\SEL[0][2] , 
        \SEL[0][1] , \SEL[0][0] }) );
  BOOTH_ENCODER_1 ENCODERS_7 ( .TO_ENC(B[15:13]), .ENC({\SEL[1][2] , 
        \SEL[1][1] , \SEL[1][0] }) );
endmodule


module REG_N10 ( D, Q, EN, RST, CLK );
  input [9:0] D;
  output [9:0] Q;
  input EN, RST, CLK;
  wire   n1;

  FD_75 FF_0 ( .D(D[0]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[0]) );
  FD_74 FF_1 ( .D(D[1]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[1]) );
  FD_73 FF_2 ( .D(D[2]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[2]) );
  FD_72 FF_3 ( .D(D[3]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[3]) );
  FD_71 FF_4 ( .D(D[4]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[4]) );
  FD_70 FF_5 ( .D(D[5]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[5]) );
  FD_69 FF_6 ( .D(D[6]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[6]) );
  FD_68 FF_7 ( .D(D[7]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[7]) );
  FD_67 FF_8 ( .D(D[8]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[8]) );
  FD_66 FF_9 ( .D(D[9]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[9]) );
  BUF_X1 U1 ( .A(RST), .Z(n1) );
endmodule


module BOOTHMUL_COMP_2 ( PREVIOUS, A, NEG_A, B, P );
  input [16:0] PREVIOUS;
  input [15:0] A;
  input [15:0] NEG_A;
  input [15:0] B;
  output [22:0] P;
  wire   \SEL[2][2] , \SEL[2][1] , \SEL[2][0] , \SEL[1][2] , \SEL[1][1] ,
         \SEL[1][0] , \SEL[0][2] , \SEL[0][1] , \SEL[0][0] , \IN_B_RCA[2][18] ,
         \IN_B_RCA[2][17] , \IN_B_RCA[2][16] , \IN_B_RCA[2][15] ,
         \IN_B_RCA[2][14] , \IN_B_RCA[2][13] , \IN_B_RCA[2][12] ,
         \IN_B_RCA[2][11] , \IN_B_RCA[2][10] , \IN_B_RCA[2][9] ,
         \IN_B_RCA[2][8] , \IN_B_RCA[2][7] , \IN_B_RCA[2][6] ,
         \IN_B_RCA[2][5] , \IN_B_RCA[2][4] , \IN_B_RCA[2][3] ,
         \IN_B_RCA[2][2] , \IN_B_RCA[2][1] , \IN_B_RCA[2][0] ,
         \IN_B_RCA[1][18] , \IN_B_RCA[1][17] , \IN_B_RCA[1][16] ,
         \IN_B_RCA[1][15] , \IN_B_RCA[1][14] , \IN_B_RCA[1][13] ,
         \IN_B_RCA[1][12] , \IN_B_RCA[1][11] , \IN_B_RCA[1][10] ,
         \IN_B_RCA[1][9] , \IN_B_RCA[1][8] , \IN_B_RCA[1][7] ,
         \IN_B_RCA[1][6] , \IN_B_RCA[1][5] , \IN_B_RCA[1][4] ,
         \IN_B_RCA[1][3] , \IN_B_RCA[1][2] , \IN_B_RCA[1][1] ,
         \IN_B_RCA[1][0] , \IN_B_RCA[0][18] , \IN_B_RCA[0][17] ,
         \IN_B_RCA[0][16] , \IN_B_RCA[0][15] , \IN_B_RCA[0][14] ,
         \IN_B_RCA[0][13] , \IN_B_RCA[0][12] , \IN_B_RCA[0][11] ,
         \IN_B_RCA[0][10] , \IN_B_RCA[0][9] , \IN_B_RCA[0][8] ,
         \IN_B_RCA[0][7] , \IN_B_RCA[0][6] , \IN_B_RCA[0][5] ,
         \IN_B_RCA[0][4] , \IN_B_RCA[0][3] , \IN_B_RCA[0][2] ,
         \IN_B_RCA[0][1] , \IN_B_RCA[0][0] , \IN_A_RCA[2][18] ,
         \IN_A_RCA[2][15] , \IN_A_RCA[2][14] , \IN_A_RCA[2][13] ,
         \IN_A_RCA[2][12] , \IN_A_RCA[2][11] , \IN_A_RCA[2][10] ,
         \IN_A_RCA[2][9] , \IN_A_RCA[2][8] , \IN_A_RCA[2][7] ,
         \IN_A_RCA[2][6] , \IN_A_RCA[2][5] , \IN_A_RCA[2][4] ,
         \IN_A_RCA[2][3] , \IN_A_RCA[2][2] , \IN_A_RCA[2][1] ,
         \IN_A_RCA[2][0] , \IN_A_RCA[1][18] , \IN_A_RCA[1][15] ,
         \IN_A_RCA[1][14] , \IN_A_RCA[1][13] , \IN_A_RCA[1][12] ,
         \IN_A_RCA[1][11] , \IN_A_RCA[1][10] , \IN_A_RCA[1][9] ,
         \IN_A_RCA[1][8] , \IN_A_RCA[1][7] , \IN_A_RCA[1][6] ,
         \IN_A_RCA[1][5] , \IN_A_RCA[1][4] , \IN_A_RCA[1][3] ,
         \IN_A_RCA[1][2] , \IN_A_RCA[1][1] , \IN_A_RCA[1][0] , n1, n2, n3, n4,
         n5;

  MUX51_GEN_N19_5 MUX_INST_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({A[15], A, 1'b0, 1'b0}), .C({NEG_A[15], NEG_A, 1'b0, 1'b0}), .D({A, 1'b0, 
        1'b0, 1'b0}), .E({NEG_A, 1'b0, 1'b0, 1'b0}), .SEL({\SEL[0][2] , 
        \SEL[0][1] , \SEL[0][0] }), .Y({\IN_B_RCA[0][18] , \IN_B_RCA[0][17] , 
        \IN_B_RCA[0][16] , \IN_B_RCA[0][15] , \IN_B_RCA[0][14] , 
        \IN_B_RCA[0][13] , \IN_B_RCA[0][12] , \IN_B_RCA[0][11] , 
        \IN_B_RCA[0][10] , \IN_B_RCA[0][9] , \IN_B_RCA[0][8] , 
        \IN_B_RCA[0][7] , \IN_B_RCA[0][6] , \IN_B_RCA[0][5] , \IN_B_RCA[0][4] , 
        \IN_B_RCA[0][3] , \IN_B_RCA[0][2] , \IN_B_RCA[0][1] , \IN_B_RCA[0][0] }) );
  MUX51_GEN_N19_4 MUX_INST_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({A[15], A, 1'b0, 1'b0}), .C({NEG_A[15], NEG_A, 1'b0, 1'b0}), .D({A, 1'b0, 
        1'b0, 1'b0}), .E({NEG_A, 1'b0, 1'b0, 1'b0}), .SEL({\SEL[1][2] , 
        \SEL[1][1] , \SEL[1][0] }), .Y({\IN_B_RCA[1][18] , \IN_B_RCA[1][17] , 
        \IN_B_RCA[1][16] , \IN_B_RCA[1][15] , \IN_B_RCA[1][14] , 
        \IN_B_RCA[1][13] , \IN_B_RCA[1][12] , \IN_B_RCA[1][11] , 
        \IN_B_RCA[1][10] , \IN_B_RCA[1][9] , \IN_B_RCA[1][8] , 
        \IN_B_RCA[1][7] , \IN_B_RCA[1][6] , \IN_B_RCA[1][5] , \IN_B_RCA[1][4] , 
        \IN_B_RCA[1][3] , \IN_B_RCA[1][2] , \IN_B_RCA[1][1] , \IN_B_RCA[1][0] }) );
  MUX51_GEN_N19_3 MUX_INST_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({A[15], A, 1'b0, 1'b0}), .C({NEG_A[15], NEG_A, 1'b0, 1'b0}), .D({A, 1'b0, 
        1'b0, 1'b0}), .E({NEG_A, 1'b0, 1'b0, 1'b0}), .SEL({\SEL[2][2] , 
        \SEL[2][1] , \SEL[2][0] }), .Y({\IN_B_RCA[2][18] , \IN_B_RCA[2][17] , 
        \IN_B_RCA[2][16] , \IN_B_RCA[2][15] , \IN_B_RCA[2][14] , 
        \IN_B_RCA[2][13] , \IN_B_RCA[2][12] , \IN_B_RCA[2][11] , 
        \IN_B_RCA[2][10] , \IN_B_RCA[2][9] , \IN_B_RCA[2][8] , 
        \IN_B_RCA[2][7] , \IN_B_RCA[2][6] , \IN_B_RCA[2][5] , \IN_B_RCA[2][4] , 
        \IN_B_RCA[2][3] , \IN_B_RCA[2][2] , \IN_B_RCA[2][1] , \IN_B_RCA[2][0] }) );
  RCA_GEN_NO_C_N19_5 RCA_INST_1_0 ( .A({PREVIOUS[16], PREVIOUS[16], PREVIOUS}), 
        .B({\IN_B_RCA[0][18] , \IN_B_RCA[0][17] , \IN_B_RCA[0][16] , 
        \IN_B_RCA[0][15] , \IN_B_RCA[0][14] , \IN_B_RCA[0][13] , 
        \IN_B_RCA[0][12] , \IN_B_RCA[0][11] , \IN_B_RCA[0][10] , 
        \IN_B_RCA[0][9] , \IN_B_RCA[0][8] , \IN_B_RCA[0][7] , \IN_B_RCA[0][6] , 
        \IN_B_RCA[0][5] , \IN_B_RCA[0][4] , \IN_B_RCA[0][3] , \IN_B_RCA[0][2] , 
        \IN_B_RCA[0][1] , \IN_B_RCA[0][0] }), .S({\IN_A_RCA[1][18] , 
        \IN_A_RCA[1][15] , \IN_A_RCA[1][14] , \IN_A_RCA[1][13] , 
        \IN_A_RCA[1][12] , \IN_A_RCA[1][11] , \IN_A_RCA[1][10] , 
        \IN_A_RCA[1][9] , \IN_A_RCA[1][8] , \IN_A_RCA[1][7] , \IN_A_RCA[1][6] , 
        \IN_A_RCA[1][5] , \IN_A_RCA[1][4] , \IN_A_RCA[1][3] , \IN_A_RCA[1][2] , 
        \IN_A_RCA[1][1] , \IN_A_RCA[1][0] , P[1:0]}) );
  RCA_GEN_NO_C_N19_4 RCA_INST_1_1 ( .A({\IN_A_RCA[1][18] , \IN_A_RCA[1][18] , 
        \IN_A_RCA[1][18] , \IN_A_RCA[1][15] , \IN_A_RCA[1][14] , 
        \IN_A_RCA[1][13] , \IN_A_RCA[1][12] , \IN_A_RCA[1][11] , 
        \IN_A_RCA[1][10] , \IN_A_RCA[1][9] , \IN_A_RCA[1][8] , 
        \IN_A_RCA[1][7] , \IN_A_RCA[1][6] , \IN_A_RCA[1][5] , \IN_A_RCA[1][4] , 
        \IN_A_RCA[1][3] , \IN_A_RCA[1][2] , \IN_A_RCA[1][1] , \IN_A_RCA[1][0] }), .B({\IN_B_RCA[1][18] , \IN_B_RCA[1][17] , \IN_B_RCA[1][16] , 
        \IN_B_RCA[1][15] , \IN_B_RCA[1][14] , \IN_B_RCA[1][13] , 
        \IN_B_RCA[1][12] , \IN_B_RCA[1][11] , \IN_B_RCA[1][10] , 
        \IN_B_RCA[1][9] , \IN_B_RCA[1][8] , \IN_B_RCA[1][7] , \IN_B_RCA[1][6] , 
        \IN_B_RCA[1][5] , \IN_B_RCA[1][4] , \IN_B_RCA[1][3] , \IN_B_RCA[1][2] , 
        \IN_B_RCA[1][1] , \IN_B_RCA[1][0] }), .S({\IN_A_RCA[2][18] , 
        \IN_A_RCA[2][15] , \IN_A_RCA[2][14] , \IN_A_RCA[2][13] , 
        \IN_A_RCA[2][12] , \IN_A_RCA[2][11] , \IN_A_RCA[2][10] , 
        \IN_A_RCA[2][9] , \IN_A_RCA[2][8] , \IN_A_RCA[2][7] , \IN_A_RCA[2][6] , 
        \IN_A_RCA[2][5] , \IN_A_RCA[2][4] , \IN_A_RCA[2][3] , \IN_A_RCA[2][2] , 
        \IN_A_RCA[2][1] , \IN_A_RCA[2][0] , P[3:2]}) );
  RCA_GEN_NO_C_N19_3 RCA_INST_1_2 ( .A({n3, n2, \IN_A_RCA[2][18] , 
        \IN_A_RCA[2][15] , \IN_A_RCA[2][14] , \IN_A_RCA[2][13] , 
        \IN_A_RCA[2][12] , \IN_A_RCA[2][11] , \IN_A_RCA[2][10] , 
        \IN_A_RCA[2][9] , \IN_A_RCA[2][8] , \IN_A_RCA[2][7] , \IN_A_RCA[2][6] , 
        \IN_A_RCA[2][5] , \IN_A_RCA[2][4] , \IN_A_RCA[2][3] , \IN_A_RCA[2][2] , 
        \IN_A_RCA[2][1] , \IN_A_RCA[2][0] }), .B({\IN_B_RCA[2][18] , 
        \IN_B_RCA[2][17] , \IN_B_RCA[2][16] , \IN_B_RCA[2][15] , 
        \IN_B_RCA[2][14] , \IN_B_RCA[2][13] , \IN_B_RCA[2][12] , 
        \IN_B_RCA[2][11] , \IN_B_RCA[2][10] , \IN_B_RCA[2][9] , 
        \IN_B_RCA[2][8] , \IN_B_RCA[2][7] , \IN_B_RCA[2][6] , \IN_B_RCA[2][5] , 
        \IN_B_RCA[2][4] , \IN_B_RCA[2][3] , \IN_B_RCA[2][2] , \IN_B_RCA[2][1] , 
        \IN_B_RCA[2][0] }), .S(P[22:4]) );
  BOOTH_ENCODER_5 ENCODERS_3 ( .TO_ENC(B[7:5]), .ENC({\SEL[0][2] , \SEL[0][1] , 
        \SEL[0][0] }) );
  BOOTH_ENCODER_4 ENCODERS_4 ( .TO_ENC({B[9:8], n5}), .ENC({\SEL[1][2] , 
        \SEL[1][1] , \SEL[1][0] }) );
  BOOTH_ENCODER_3 ENCODERS_5 ( .TO_ENC(B[11:9]), .ENC({\SEL[2][2] , 
        \SEL[2][1] , \SEL[2][0] }) );
  INV_X1 U2 ( .A(\IN_A_RCA[2][18] ), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(n2) );
  CLKBUF_X1 U4 ( .A(n2), .Z(n3) );
  INV_X1 U5 ( .A(B[7]), .ZN(n4) );
  INV_X1 U6 ( .A(n4), .ZN(n5) );
endmodule


module REG_N16_0 ( D, Q, EN, RST, CLK );
  input [15:0] D;
  output [15:0] Q;
  input EN, RST, CLK;
  wire   n1, n2;

  FD_123 FF_0 ( .D(D[0]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[0]) );
  FD_122 FF_1 ( .D(D[1]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[1]) );
  FD_121 FF_2 ( .D(D[2]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[2]) );
  FD_120 FF_3 ( .D(D[3]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[3]) );
  FD_119 FF_4 ( .D(D[4]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[4]) );
  FD_118 FF_5 ( .D(D[5]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[5]) );
  FD_117 FF_6 ( .D(D[6]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[6]) );
  FD_116 FF_7 ( .D(D[7]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[7]) );
  FD_115 FF_8 ( .D(D[8]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[8]) );
  FD_114 FF_9 ( .D(D[9]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[9]) );
  FD_113 FF_10 ( .D(D[10]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[10]) );
  FD_112 FF_11 ( .D(D[11]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[11]) );
  FD_111 FF_12 ( .D(D[12]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[12]) );
  FD_110 FF_13 ( .D(D[13]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[13]) );
  FD_109 FF_14 ( .D(D[14]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[14]) );
  FD_108 FF_15 ( .D(D[15]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[15]) );
  BUF_X1 U1 ( .A(RST), .Z(n1) );
  BUF_X1 U2 ( .A(RST), .Z(n2) );
endmodule


module REG_N17_0 ( D, Q, EN, RST, CLK );
  input [16:0] D;
  output [16:0] Q;
  input EN, RST, CLK;
  wire   n1, n2;

  FD_140 FF_0 ( .D(D[0]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[0]) );
  FD_139 FF_1 ( .D(D[1]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[1]) );
  FD_138 FF_2 ( .D(D[2]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[2]) );
  FD_137 FF_3 ( .D(D[3]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[3]) );
  FD_136 FF_4 ( .D(D[4]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[4]) );
  FD_135 FF_5 ( .D(D[5]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[5]) );
  FD_134 FF_6 ( .D(D[6]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[6]) );
  FD_133 FF_7 ( .D(D[7]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[7]) );
  FD_132 FF_8 ( .D(D[8]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[8]) );
  FD_131 FF_9 ( .D(D[9]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[9]) );
  FD_130 FF_10 ( .D(D[10]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[10]) );
  FD_129 FF_11 ( .D(D[11]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[11]) );
  FD_128 FF_12 ( .D(D[12]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[12]) );
  FD_127 FF_13 ( .D(D[13]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[13]) );
  FD_126 FF_14 ( .D(D[14]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[14]) );
  FD_125 FF_15 ( .D(D[15]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[15]) );
  FD_124 FF_16 ( .D(D[16]), .CLK(CLK), .EN(EN), .RST(n2), .Q(Q[16]) );
  BUF_X1 U1 ( .A(RST), .Z(n1) );
  BUF_X1 U2 ( .A(RST), .Z(n2) );
endmodule


module REG_N4 ( D, Q, EN, RST, CLK );
  input [3:0] D;
  output [3:0] Q;
  input EN, RST, CLK;


  FD_144 FF_0 ( .D(D[0]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[0]) );
  FD_143 FF_1 ( .D(D[1]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[1]) );
  FD_142 FF_2 ( .D(D[2]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[2]) );
  FD_141 FF_3 ( .D(D[3]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[3]) );
endmodule


module BOOTHMUL_COMP_1 ( A, NEG_A, B, P );
  input [15:0] A;
  input [15:0] NEG_A;
  input [15:0] B;
  output [20:0] P;
  wire   \SEL[2][2] , \SEL[2][1] , \SEL[2][0] , \SEL[1][2] , \SEL[1][1] ,
         \SEL[1][0] , \SEL[0][2] , \SEL[0][1] , \SEL[0][0] , \IN_B_RCA[1][18] ,
         \IN_B_RCA[1][17] , \IN_B_RCA[1][16] , \IN_B_RCA[1][15] ,
         \IN_B_RCA[1][14] , \IN_B_RCA[1][13] , \IN_B_RCA[1][12] ,
         \IN_B_RCA[1][11] , \IN_B_RCA[1][10] , \IN_B_RCA[1][9] ,
         \IN_B_RCA[1][8] , \IN_B_RCA[1][7] , \IN_B_RCA[1][6] ,
         \IN_B_RCA[1][5] , \IN_B_RCA[1][4] , \IN_B_RCA[1][3] ,
         \IN_B_RCA[1][2] , \IN_B_RCA[1][1] , \IN_B_RCA[1][0] ,
         \IN_B_RCA[0][18] , \IN_B_RCA[0][17] , \IN_B_RCA[0][16] ,
         \IN_B_RCA[0][15] , \IN_B_RCA[0][14] , \IN_B_RCA[0][13] ,
         \IN_B_RCA[0][12] , \IN_B_RCA[0][11] , \IN_B_RCA[0][10] ,
         \IN_B_RCA[0][9] , \IN_B_RCA[0][8] , \IN_B_RCA[0][7] ,
         \IN_B_RCA[0][6] , \IN_B_RCA[0][5] , \IN_B_RCA[0][4] ,
         \IN_B_RCA[0][3] , \IN_B_RCA[0][2] , \IN_B_RCA[0][1] ,
         \IN_B_RCA[0][0] , \IN_A_RCA[1][18] , \IN_A_RCA[1][15] ,
         \IN_A_RCA[1][14] , \IN_A_RCA[1][13] , \IN_A_RCA[1][12] ,
         \IN_A_RCA[1][11] , \IN_A_RCA[1][10] , \IN_A_RCA[1][9] ,
         \IN_A_RCA[1][8] , \IN_A_RCA[1][7] , \IN_A_RCA[1][6] ,
         \IN_A_RCA[1][5] , \IN_A_RCA[1][4] , \IN_A_RCA[1][3] ,
         \IN_A_RCA[1][2] , \IN_A_RCA[1][1] , \IN_A_RCA[1][0] ,
         \IN_A_RCA[0][18] , \IN_A_RCA[0][17] , \IN_A_RCA[0][16] ,
         \IN_A_RCA[0][15] , \IN_A_RCA[0][14] , \IN_A_RCA[0][13] ,
         \IN_A_RCA[0][12] , \IN_A_RCA[0][11] , \IN_A_RCA[0][10] ,
         \IN_A_RCA[0][9] , \IN_A_RCA[0][8] , \IN_A_RCA[0][7] ,
         \IN_A_RCA[0][6] , \IN_A_RCA[0][5] , \IN_A_RCA[0][4] ,
         \IN_A_RCA[0][3] , \IN_A_RCA[0][2] , \IN_A_RCA[0][1] ,
         \IN_A_RCA[0][0] , n1, n2, n3, n4, n5;

  MUX51_GEN_N19_0 FIRST_MUX ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n5, n5, n5, n5, A[14:0]}), .C({NEG_A[15], NEG_A[15], NEG_A[15], NEG_A}), 
        .D({n5, n5, n5, A[14:0], 1'b0}), .E({NEG_A[15], NEG_A[15], NEG_A[15], 
        n3, n1, n4, n2, NEG_A[10:0], 1'b0}), .SEL({\SEL[0][2] , \SEL[0][1] , 
        \SEL[0][0] }), .Y({\IN_A_RCA[0][18] , \IN_A_RCA[0][17] , 
        \IN_A_RCA[0][16] , \IN_A_RCA[0][15] , \IN_A_RCA[0][14] , 
        \IN_A_RCA[0][13] , \IN_A_RCA[0][12] , \IN_A_RCA[0][11] , 
        \IN_A_RCA[0][10] , \IN_A_RCA[0][9] , \IN_A_RCA[0][8] , 
        \IN_A_RCA[0][7] , \IN_A_RCA[0][6] , \IN_A_RCA[0][5] , \IN_A_RCA[0][4] , 
        \IN_A_RCA[0][3] , \IN_A_RCA[0][2] , \IN_A_RCA[0][1] , \IN_A_RCA[0][0] }) );
  MUX51_GEN_N19_7 MUX_INST_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n5, n5, A[14:0], 1'b0, 1'b0}), .C({NEG_A[15], NEG_A[15], n3, n1, n4, n2, 
        NEG_A[10:0], 1'b0, 1'b0}), .D({n5, A[14:0], 1'b0, 1'b0, 1'b0}), .E({
        NEG_A[15], n3, n1, n4, n2, NEG_A[10:0], 1'b0, 1'b0, 1'b0}), .SEL({
        \SEL[1][2] , \SEL[1][1] , \SEL[1][0] }), .Y({\IN_B_RCA[0][18] , 
        \IN_B_RCA[0][17] , \IN_B_RCA[0][16] , \IN_B_RCA[0][15] , 
        \IN_B_RCA[0][14] , \IN_B_RCA[0][13] , \IN_B_RCA[0][12] , 
        \IN_B_RCA[0][11] , \IN_B_RCA[0][10] , \IN_B_RCA[0][9] , 
        \IN_B_RCA[0][8] , \IN_B_RCA[0][7] , \IN_B_RCA[0][6] , \IN_B_RCA[0][5] , 
        \IN_B_RCA[0][4] , \IN_B_RCA[0][3] , \IN_B_RCA[0][2] , \IN_B_RCA[0][1] , 
        \IN_B_RCA[0][0] }) );
  MUX51_GEN_N19_6 MUX_INST_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n5, n5, A[14:0], 1'b0, 1'b0}), .C({NEG_A[15], NEG_A[15], n3, n1, n4, n2, 
        NEG_A[10:0], 1'b0, 1'b0}), .D({n5, A[14:0], 1'b0, 1'b0, 1'b0}), .E({
        NEG_A[15], n3, n1, n4, n2, NEG_A[10:0], 1'b0, 1'b0, 1'b0}), .SEL({
        \SEL[2][2] , \SEL[2][1] , \SEL[2][0] }), .Y({\IN_B_RCA[1][18] , 
        \IN_B_RCA[1][17] , \IN_B_RCA[1][16] , \IN_B_RCA[1][15] , 
        \IN_B_RCA[1][14] , \IN_B_RCA[1][13] , \IN_B_RCA[1][12] , 
        \IN_B_RCA[1][11] , \IN_B_RCA[1][10] , \IN_B_RCA[1][9] , 
        \IN_B_RCA[1][8] , \IN_B_RCA[1][7] , \IN_B_RCA[1][6] , \IN_B_RCA[1][5] , 
        \IN_B_RCA[1][4] , \IN_B_RCA[1][3] , \IN_B_RCA[1][2] , \IN_B_RCA[1][1] , 
        \IN_B_RCA[1][0] }) );
  RCA_GEN_NO_C_N19_0 RCA_INST_1_0 ( .A({\IN_A_RCA[0][18] , \IN_A_RCA[0][17] , 
        \IN_A_RCA[0][16] , \IN_A_RCA[0][15] , \IN_A_RCA[0][14] , 
        \IN_A_RCA[0][13] , \IN_A_RCA[0][12] , \IN_A_RCA[0][11] , 
        \IN_A_RCA[0][10] , \IN_A_RCA[0][9] , \IN_A_RCA[0][8] , 
        \IN_A_RCA[0][7] , \IN_A_RCA[0][6] , \IN_A_RCA[0][5] , \IN_A_RCA[0][4] , 
        \IN_A_RCA[0][3] , \IN_A_RCA[0][2] , \IN_A_RCA[0][1] , \IN_A_RCA[0][0] }), .B({\IN_B_RCA[0][18] , \IN_B_RCA[0][17] , \IN_B_RCA[0][16] , 
        \IN_B_RCA[0][15] , \IN_B_RCA[0][14] , \IN_B_RCA[0][13] , 
        \IN_B_RCA[0][12] , \IN_B_RCA[0][11] , \IN_B_RCA[0][10] , 
        \IN_B_RCA[0][9] , \IN_B_RCA[0][8] , \IN_B_RCA[0][7] , \IN_B_RCA[0][6] , 
        \IN_B_RCA[0][5] , \IN_B_RCA[0][4] , \IN_B_RCA[0][3] , \IN_B_RCA[0][2] , 
        \IN_B_RCA[0][1] , \IN_B_RCA[0][0] }), .S({\IN_A_RCA[1][18] , 
        \IN_A_RCA[1][15] , \IN_A_RCA[1][14] , \IN_A_RCA[1][13] , 
        \IN_A_RCA[1][12] , \IN_A_RCA[1][11] , \IN_A_RCA[1][10] , 
        \IN_A_RCA[1][9] , \IN_A_RCA[1][8] , \IN_A_RCA[1][7] , \IN_A_RCA[1][6] , 
        \IN_A_RCA[1][5] , \IN_A_RCA[1][4] , \IN_A_RCA[1][3] , \IN_A_RCA[1][2] , 
        \IN_A_RCA[1][1] , \IN_A_RCA[1][0] , P[1:0]}) );
  RCA_GEN_NO_C_N19_6 RCA_INST_1_1 ( .A({\IN_A_RCA[1][18] , \IN_A_RCA[1][18] , 
        \IN_A_RCA[1][18] , \IN_A_RCA[1][15] , \IN_A_RCA[1][14] , 
        \IN_A_RCA[1][13] , \IN_A_RCA[1][12] , \IN_A_RCA[1][11] , 
        \IN_A_RCA[1][10] , \IN_A_RCA[1][9] , \IN_A_RCA[1][8] , 
        \IN_A_RCA[1][7] , \IN_A_RCA[1][6] , \IN_A_RCA[1][5] , \IN_A_RCA[1][4] , 
        \IN_A_RCA[1][3] , \IN_A_RCA[1][2] , \IN_A_RCA[1][1] , \IN_A_RCA[1][0] }), .B({\IN_B_RCA[1][18] , \IN_B_RCA[1][17] , \IN_B_RCA[1][16] , 
        \IN_B_RCA[1][15] , \IN_B_RCA[1][14] , \IN_B_RCA[1][13] , 
        \IN_B_RCA[1][12] , \IN_B_RCA[1][11] , \IN_B_RCA[1][10] , 
        \IN_B_RCA[1][9] , \IN_B_RCA[1][8] , \IN_B_RCA[1][7] , \IN_B_RCA[1][6] , 
        \IN_B_RCA[1][5] , \IN_B_RCA[1][4] , \IN_B_RCA[1][3] , \IN_B_RCA[1][2] , 
        \IN_B_RCA[1][1] , \IN_B_RCA[1][0] }), .S(P[20:2]) );
  BOOTH_ENCODER_0 ENCODERS_0 ( .TO_ENC({B[1:0], 1'b0}), .ENC({\SEL[0][2] , 
        \SEL[0][1] , \SEL[0][0] }) );
  BOOTH_ENCODER_7 ENCODERS_1 ( .TO_ENC(B[3:1]), .ENC({\SEL[1][2] , \SEL[1][1] , 
        \SEL[1][0] }) );
  BOOTH_ENCODER_6 ENCODERS_2 ( .TO_ENC(B[5:3]), .ENC({\SEL[2][2] , \SEL[2][1] , 
        \SEL[2][0] }) );
  CLKBUF_X1 U2 ( .A(NEG_A[13]), .Z(n1) );
  CLKBUF_X1 U3 ( .A(NEG_A[11]), .Z(n2) );
  CLKBUF_X1 U4 ( .A(NEG_A[14]), .Z(n3) );
  CLKBUF_X1 U5 ( .A(NEG_A[12]), .Z(n4) );
  BUF_X1 U6 ( .A(A[15]), .Z(n5) );
endmodule


module RCA_GEN_NO_C_N16 ( A, B, S, Co );
  input [15:0] A;
  input [15:0] B;
  output [15:0] S;
  output Co;

  wire   [14:0] CTMP;

  HA_8 HA_INST ( .A(A[0]), .B(B[0]), .S(S[0]), .Co(CTMP[0]) );
  FA_205 FAI_0 ( .A(A[1]), .B(B[1]), .Ci(CTMP[0]), .S(S[1]), .Co(CTMP[1]) );
  FA_204 FAI_1 ( .A(A[2]), .B(B[2]), .Ci(CTMP[1]), .S(S[2]), .Co(CTMP[2]) );
  FA_203 FAI_2 ( .A(A[3]), .B(B[3]), .Ci(CTMP[2]), .S(S[3]), .Co(CTMP[3]) );
  FA_202 FAI_3 ( .A(A[4]), .B(B[4]), .Ci(CTMP[3]), .S(S[4]), .Co(CTMP[4]) );
  FA_201 FAI_4 ( .A(A[5]), .B(B[5]), .Ci(CTMP[4]), .S(S[5]), .Co(CTMP[5]) );
  FA_200 FAI_5 ( .A(A[6]), .B(B[6]), .Ci(CTMP[5]), .S(S[6]), .Co(CTMP[6]) );
  FA_199 FAI_6 ( .A(A[7]), .B(B[7]), .Ci(CTMP[6]), .S(S[7]), .Co(CTMP[7]) );
  FA_198 FAI_7 ( .A(A[8]), .B(B[8]), .Ci(CTMP[7]), .S(S[8]), .Co(CTMP[8]) );
  FA_197 FAI_8 ( .A(A[9]), .B(B[9]), .Ci(CTMP[8]), .S(S[9]), .Co(CTMP[9]) );
  FA_196 FAI_9 ( .A(A[10]), .B(B[10]), .Ci(CTMP[9]), .S(S[10]), .Co(CTMP[10])
         );
  FA_195 FAI_10 ( .A(A[11]), .B(B[11]), .Ci(CTMP[10]), .S(S[11]), .Co(CTMP[11]) );
  FA_194 FAI_11 ( .A(A[12]), .B(B[12]), .Ci(CTMP[11]), .S(S[12]), .Co(CTMP[12]) );
  FA_193 FAI_12 ( .A(A[13]), .B(B[13]), .Ci(CTMP[12]), .S(S[13]), .Co(CTMP[13]) );
  FA_192 FAI_13 ( .A(A[14]), .B(B[14]), .Ci(CTMP[13]), .S(S[14]), .Co(CTMP[14]) );
  FA_191 FAI_14 ( .A(A[15]), .B(B[15]), .Ci(CTMP[14]), .S(S[15]), .Co(Co) );
endmodule


module MUX81_GEN_N32 ( A, B, C, D, E, F, G, H, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [31:0] F;
  input [31:0] G;
  input [31:0] H;
  input [2:0] SEL;
  output [31:0] Y;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n1, n2, n3, n4,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164;

  BUF_X1 U1 ( .A(n12), .Z(n153) );
  BUF_X1 U2 ( .A(n12), .Z(n154) );
  BUF_X1 U3 ( .A(n12), .Z(n155) );
  NOR4_X1 U4 ( .A1(n161), .A2(n149), .A3(n156), .A4(n141), .ZN(n12) );
  OR4_X1 U5 ( .A1(n3), .A2(n146), .A3(n152), .A4(n164), .ZN(n141) );
  BUF_X1 U6 ( .A(n16), .Z(n3) );
  BUF_X1 U7 ( .A(n16), .Z(n2) );
  BUF_X1 U8 ( .A(n16), .Z(n1) );
  NOR3_X1 U9 ( .A1(n143), .A2(n142), .A3(n144), .ZN(n16) );
  BUF_X1 U10 ( .A(n11), .Z(n156) );
  AOI22_X1 U11 ( .A1(G[25]), .A2(n157), .B1(H[25]), .B2(n154), .ZN(n71) );
  AOI22_X1 U12 ( .A1(G[26]), .A2(n157), .B1(H[26]), .B2(n154), .ZN(n67) );
  AOI22_X1 U13 ( .A1(G[27]), .A2(n157), .B1(H[27]), .B2(n154), .ZN(n63) );
  AOI22_X1 U14 ( .A1(G[28]), .A2(n157), .B1(H[28]), .B2(n154), .ZN(n59) );
  AOI22_X1 U15 ( .A1(G[29]), .A2(n157), .B1(H[29]), .B2(n154), .ZN(n55) );
  AOI22_X1 U16 ( .A1(G[30]), .A2(n157), .B1(H[30]), .B2(n154), .ZN(n47) );
  BUF_X1 U17 ( .A(n14), .Z(n149) );
  BUF_X1 U18 ( .A(n10), .Z(n161) );
  BUF_X1 U19 ( .A(n15), .Z(n146) );
  BUF_X1 U20 ( .A(n13), .Z(n152) );
  BUF_X1 U21 ( .A(n9), .Z(n164) );
  BUF_X1 U22 ( .A(n9), .Z(n163) );
  BUF_X1 U23 ( .A(n13), .Z(n151) );
  BUF_X1 U24 ( .A(n15), .Z(n145) );
  BUF_X1 U25 ( .A(n11), .Z(n157) );
  BUF_X1 U26 ( .A(n15), .Z(n4) );
  BUF_X1 U27 ( .A(n9), .Z(n162) );
  BUF_X1 U28 ( .A(n13), .Z(n150) );
  BUF_X1 U29 ( .A(n10), .Z(n160) );
  BUF_X1 U30 ( .A(n14), .Z(n148) );
  BUF_X1 U31 ( .A(n10), .Z(n159) );
  BUF_X1 U32 ( .A(n14), .Z(n147) );
  AOI22_X1 U33 ( .A1(D[31]), .A2(n4), .B1(A[31]), .B2(n1), .ZN(n41) );
  BUF_X1 U34 ( .A(n11), .Z(n158) );
  NOR3_X1 U35 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n143), .ZN(n15) );
  NOR3_X1 U36 ( .A1(n143), .A2(SEL[1]), .A3(n144), .ZN(n13) );
  NOR3_X1 U37 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n144), .ZN(n11) );
  NOR3_X1 U38 ( .A1(n142), .A2(SEL[2]), .A3(n144), .ZN(n10) );
  NOR3_X1 U39 ( .A1(n142), .A2(SEL[0]), .A3(n143), .ZN(n9) );
  NOR3_X1 U40 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n142), .ZN(n14) );
  AOI22_X1 U41 ( .A1(G[1]), .A2(n156), .B1(H[1]), .B2(n153), .ZN(n95) );
  AOI22_X1 U42 ( .A1(G[2]), .A2(n157), .B1(H[2]), .B2(n154), .ZN(n51) );
  AOI22_X1 U43 ( .A1(G[3]), .A2(n158), .B1(H[3]), .B2(n154), .ZN(n39) );
  AOI22_X1 U44 ( .A1(G[4]), .A2(n158), .B1(H[4]), .B2(n155), .ZN(n35) );
  AOI22_X1 U45 ( .A1(G[5]), .A2(n158), .B1(H[5]), .B2(n155), .ZN(n31) );
  AOI22_X1 U46 ( .A1(G[6]), .A2(n158), .B1(H[6]), .B2(n155), .ZN(n27) );
  AOI22_X1 U47 ( .A1(G[7]), .A2(n158), .B1(H[7]), .B2(n155), .ZN(n23) );
  AOI22_X1 U48 ( .A1(G[8]), .A2(n158), .B1(H[8]), .B2(n155), .ZN(n19) );
  AOI22_X1 U49 ( .A1(G[9]), .A2(n158), .B1(H[9]), .B2(n155), .ZN(n7) );
  AOI22_X1 U50 ( .A1(G[10]), .A2(n156), .B1(H[10]), .B2(n153), .ZN(n135) );
  AOI22_X1 U51 ( .A1(G[11]), .A2(n156), .B1(H[11]), .B2(n153), .ZN(n131) );
  AOI22_X1 U52 ( .A1(G[12]), .A2(n156), .B1(H[12]), .B2(n153), .ZN(n127) );
  AOI22_X1 U53 ( .A1(G[13]), .A2(n156), .B1(H[13]), .B2(n153), .ZN(n123) );
  AOI22_X1 U54 ( .A1(G[14]), .A2(n156), .B1(H[14]), .B2(n153), .ZN(n119) );
  AOI22_X1 U55 ( .A1(G[15]), .A2(n156), .B1(H[15]), .B2(n153), .ZN(n115) );
  AOI22_X1 U56 ( .A1(G[16]), .A2(n156), .B1(H[16]), .B2(n153), .ZN(n111) );
  AOI22_X1 U57 ( .A1(G[17]), .A2(n156), .B1(H[17]), .B2(n153), .ZN(n107) );
  AOI22_X1 U58 ( .A1(G[18]), .A2(n156), .B1(H[18]), .B2(n153), .ZN(n103) );
  AOI22_X1 U59 ( .A1(G[19]), .A2(n156), .B1(H[19]), .B2(n153), .ZN(n99) );
  AOI22_X1 U60 ( .A1(G[20]), .A2(n157), .B1(H[20]), .B2(n153), .ZN(n91) );
  AOI22_X1 U61 ( .A1(G[21]), .A2(n157), .B1(H[21]), .B2(n154), .ZN(n87) );
  AOI22_X1 U62 ( .A1(G[22]), .A2(n157), .B1(H[22]), .B2(n154), .ZN(n83) );
  AOI22_X1 U63 ( .A1(G[23]), .A2(n157), .B1(H[23]), .B2(n154), .ZN(n79) );
  AOI22_X1 U64 ( .A1(G[24]), .A2(n157), .B1(H[24]), .B2(n154), .ZN(n75) );
  AOI22_X1 U65 ( .A1(G[0]), .A2(n156), .B1(H[0]), .B2(n153), .ZN(n139) );
  AOI22_X1 U66 ( .A1(G[31]), .A2(n157), .B1(H[31]), .B2(n154), .ZN(n43) );
  INV_X1 U67 ( .A(SEL[1]), .ZN(n142) );
  INV_X1 U68 ( .A(SEL[2]), .ZN(n143) );
  INV_X1 U69 ( .A(SEL[0]), .ZN(n144) );
  AOI22_X1 U70 ( .A1(B[6]), .A2(n162), .B1(E[6]), .B2(n159), .ZN(n28) );
  AOI22_X1 U71 ( .A1(B[7]), .A2(n162), .B1(E[7]), .B2(n159), .ZN(n24) );
  AOI22_X1 U72 ( .A1(B[8]), .A2(n162), .B1(E[8]), .B2(n159), .ZN(n20) );
  AOI22_X1 U73 ( .A1(B[9]), .A2(n162), .B1(E[9]), .B2(n159), .ZN(n8) );
  AOI22_X1 U74 ( .A1(B[10]), .A2(n164), .B1(E[10]), .B2(n161), .ZN(n136) );
  AOI22_X1 U75 ( .A1(B[11]), .A2(n164), .B1(E[11]), .B2(n161), .ZN(n132) );
  AOI22_X1 U76 ( .A1(B[12]), .A2(n164), .B1(E[12]), .B2(n161), .ZN(n128) );
  AOI22_X1 U77 ( .A1(B[13]), .A2(n164), .B1(E[13]), .B2(n161), .ZN(n124) );
  AOI22_X1 U78 ( .A1(B[14]), .A2(n164), .B1(E[14]), .B2(n161), .ZN(n120) );
  AOI22_X1 U79 ( .A1(B[15]), .A2(n163), .B1(E[15]), .B2(n160), .ZN(n116) );
  AOI22_X1 U80 ( .A1(B[16]), .A2(n163), .B1(E[16]), .B2(n160), .ZN(n112) );
  AOI22_X1 U81 ( .A1(B[17]), .A2(n163), .B1(E[17]), .B2(n160), .ZN(n108) );
  AOI22_X1 U82 ( .A1(B[18]), .A2(n163), .B1(E[18]), .B2(n160), .ZN(n104) );
  AOI22_X1 U83 ( .A1(B[19]), .A2(n163), .B1(E[19]), .B2(n160), .ZN(n100) );
  AOI22_X1 U84 ( .A1(B[20]), .A2(n163), .B1(E[20]), .B2(n160), .ZN(n92) );
  AOI22_X1 U85 ( .A1(B[21]), .A2(n163), .B1(E[21]), .B2(n160), .ZN(n88) );
  AOI22_X1 U86 ( .A1(B[22]), .A2(n163), .B1(E[22]), .B2(n160), .ZN(n84) );
  AOI22_X1 U87 ( .A1(B[23]), .A2(n163), .B1(E[23]), .B2(n160), .ZN(n80) );
  AOI22_X1 U88 ( .A1(B[24]), .A2(n163), .B1(E[24]), .B2(n160), .ZN(n76) );
  AOI22_X1 U89 ( .A1(B[25]), .A2(n163), .B1(E[25]), .B2(n160), .ZN(n72) );
  AOI22_X1 U90 ( .A1(B[26]), .A2(n163), .B1(E[26]), .B2(n160), .ZN(n68) );
  AOI22_X1 U91 ( .A1(B[27]), .A2(n162), .B1(E[27]), .B2(n159), .ZN(n64) );
  AOI22_X1 U92 ( .A1(B[28]), .A2(n162), .B1(E[28]), .B2(n159), .ZN(n60) );
  AOI22_X1 U93 ( .A1(B[29]), .A2(n162), .B1(E[29]), .B2(n159), .ZN(n56) );
  AOI22_X1 U94 ( .A1(B[0]), .A2(n164), .B1(E[0]), .B2(n161), .ZN(n140) );
  AOI22_X1 U95 ( .A1(B[3]), .A2(n162), .B1(E[3]), .B2(n159), .ZN(n40) );
  AOI22_X1 U96 ( .A1(B[4]), .A2(n162), .B1(E[4]), .B2(n159), .ZN(n36) );
  AOI22_X1 U97 ( .A1(B[5]), .A2(n162), .B1(E[5]), .B2(n159), .ZN(n32) );
  AOI22_X1 U98 ( .A1(C[10]), .A2(n152), .B1(F[10]), .B2(n149), .ZN(n134) );
  AOI22_X1 U99 ( .A1(C[11]), .A2(n152), .B1(F[11]), .B2(n149), .ZN(n130) );
  AOI22_X1 U100 ( .A1(C[12]), .A2(n152), .B1(F[12]), .B2(n149), .ZN(n126) );
  AOI22_X1 U101 ( .A1(C[13]), .A2(n152), .B1(F[13]), .B2(n149), .ZN(n122) );
  AOI22_X1 U102 ( .A1(C[14]), .A2(n152), .B1(F[14]), .B2(n149), .ZN(n118) );
  AOI22_X1 U103 ( .A1(C[15]), .A2(n152), .B1(F[15]), .B2(n149), .ZN(n114) );
  AOI22_X1 U104 ( .A1(C[16]), .A2(n151), .B1(F[16]), .B2(n148), .ZN(n110) );
  AOI22_X1 U105 ( .A1(C[17]), .A2(n151), .B1(F[17]), .B2(n148), .ZN(n106) );
  AOI22_X1 U106 ( .A1(C[18]), .A2(n151), .B1(F[18]), .B2(n148), .ZN(n102) );
  AOI22_X1 U107 ( .A1(C[19]), .A2(n151), .B1(F[19]), .B2(n148), .ZN(n98) );
  AOI22_X1 U108 ( .A1(C[20]), .A2(n151), .B1(F[20]), .B2(n148), .ZN(n90) );
  AOI22_X1 U109 ( .A1(C[21]), .A2(n151), .B1(F[21]), .B2(n148), .ZN(n86) );
  AOI22_X1 U110 ( .A1(C[22]), .A2(n151), .B1(F[22]), .B2(n148), .ZN(n82) );
  AOI22_X1 U111 ( .A1(C[23]), .A2(n151), .B1(F[23]), .B2(n148), .ZN(n78) );
  AOI22_X1 U112 ( .A1(C[24]), .A2(n151), .B1(F[24]), .B2(n148), .ZN(n74) );
  AOI22_X1 U113 ( .A1(C[25]), .A2(n151), .B1(F[25]), .B2(n148), .ZN(n70) );
  AOI22_X1 U114 ( .A1(C[26]), .A2(n151), .B1(F[26]), .B2(n148), .ZN(n66) );
  AOI22_X1 U115 ( .A1(D[27]), .A2(n4), .B1(A[27]), .B2(n1), .ZN(n61) );
  AOI22_X1 U116 ( .A1(D[28]), .A2(n4), .B1(A[28]), .B2(n1), .ZN(n57) );
  AOI22_X1 U117 ( .A1(C[0]), .A2(n150), .B1(F[0]), .B2(n147), .ZN(n138) );
  AOI22_X1 U118 ( .A1(C[1]), .A2(n151), .B1(F[1]), .B2(n148), .ZN(n94) );
  AOI22_X1 U119 ( .A1(C[2]), .A2(n150), .B1(F[2]), .B2(n147), .ZN(n50) );
  AOI22_X1 U120 ( .A1(D[29]), .A2(n4), .B1(A[29]), .B2(n1), .ZN(n53) );
  AOI22_X1 U121 ( .A1(D[30]), .A2(n4), .B1(A[30]), .B2(n1), .ZN(n45) );
  NAND4_X1 U122 ( .A1(n37), .A2(n38), .A3(n39), .A4(n40), .ZN(Y[3]) );
  AOI22_X1 U123 ( .A1(D[3]), .A2(n4), .B1(A[3]), .B2(n1), .ZN(n37) );
  AOI22_X1 U124 ( .A1(C[3]), .A2(n150), .B1(F[3]), .B2(n147), .ZN(n38) );
  NAND4_X1 U125 ( .A1(n33), .A2(n34), .A3(n35), .A4(n36), .ZN(Y[4]) );
  AOI22_X1 U126 ( .A1(D[4]), .A2(n4), .B1(A[4]), .B2(n1), .ZN(n33) );
  AOI22_X1 U127 ( .A1(C[4]), .A2(n150), .B1(F[4]), .B2(n147), .ZN(n34) );
  NAND4_X1 U128 ( .A1(n29), .A2(n30), .A3(n31), .A4(n32), .ZN(Y[5]) );
  AOI22_X1 U129 ( .A1(D[5]), .A2(n4), .B1(A[5]), .B2(n1), .ZN(n29) );
  AOI22_X1 U130 ( .A1(C[5]), .A2(n150), .B1(F[5]), .B2(n147), .ZN(n30) );
  NAND4_X1 U131 ( .A1(n25), .A2(n26), .A3(n27), .A4(n28), .ZN(Y[6]) );
  AOI22_X1 U132 ( .A1(D[6]), .A2(n4), .B1(A[6]), .B2(n1), .ZN(n25) );
  AOI22_X1 U133 ( .A1(C[6]), .A2(n150), .B1(F[6]), .B2(n147), .ZN(n26) );
  NAND4_X1 U134 ( .A1(n21), .A2(n22), .A3(n23), .A4(n24), .ZN(Y[7]) );
  AOI22_X1 U135 ( .A1(D[7]), .A2(n4), .B1(A[7]), .B2(n1), .ZN(n21) );
  AOI22_X1 U136 ( .A1(C[7]), .A2(n150), .B1(F[7]), .B2(n147), .ZN(n22) );
  NAND4_X1 U137 ( .A1(n17), .A2(n18), .A3(n19), .A4(n20), .ZN(Y[8]) );
  AOI22_X1 U138 ( .A1(D[8]), .A2(n4), .B1(A[8]), .B2(n1), .ZN(n17) );
  AOI22_X1 U139 ( .A1(C[8]), .A2(n150), .B1(F[8]), .B2(n147), .ZN(n18) );
  NAND4_X1 U140 ( .A1(n5), .A2(n6), .A3(n7), .A4(n8), .ZN(Y[9]) );
  AOI22_X1 U141 ( .A1(D[9]), .A2(n145), .B1(A[9]), .B2(n2), .ZN(n5) );
  AOI22_X1 U142 ( .A1(C[9]), .A2(n151), .B1(F[9]), .B2(n148), .ZN(n6) );
  NAND4_X1 U143 ( .A1(n137), .A2(n138), .A3(n139), .A4(n140), .ZN(Y[0]) );
  AOI22_X1 U144 ( .A1(D[0]), .A2(n4), .B1(A[0]), .B2(n1), .ZN(n137) );
  NAND4_X1 U145 ( .A1(n53), .A2(n54), .A3(n55), .A4(n56), .ZN(Y[29]) );
  AOI22_X1 U146 ( .A1(C[29]), .A2(n150), .B1(F[29]), .B2(n147), .ZN(n54) );
  NAND4_X1 U147 ( .A1(n45), .A2(n46), .A3(n47), .A4(n48), .ZN(Y[30]) );
  AOI22_X1 U148 ( .A1(C[30]), .A2(n150), .B1(F[30]), .B2(n147), .ZN(n46) );
  AOI22_X1 U149 ( .A1(B[30]), .A2(n162), .B1(E[30]), .B2(n159), .ZN(n48) );
  NAND4_X1 U150 ( .A1(n41), .A2(n42), .A3(n43), .A4(n44), .ZN(Y[31]) );
  AOI22_X1 U151 ( .A1(C[31]), .A2(n150), .B1(F[31]), .B2(n147), .ZN(n42) );
  AOI22_X1 U152 ( .A1(B[31]), .A2(n162), .B1(E[31]), .B2(n159), .ZN(n44) );
  NAND4_X1 U153 ( .A1(n93), .A2(n94), .A3(n95), .A4(n96), .ZN(Y[1]) );
  AOI22_X1 U154 ( .A1(D[1]), .A2(n145), .B1(A[1]), .B2(n2), .ZN(n93) );
  AOI22_X1 U155 ( .A1(B[1]), .A2(n163), .B1(E[1]), .B2(n160), .ZN(n96) );
  NAND4_X1 U156 ( .A1(n49), .A2(n50), .A3(n51), .A4(n52), .ZN(Y[2]) );
  AOI22_X1 U157 ( .A1(D[2]), .A2(n4), .B1(A[2]), .B2(n1), .ZN(n49) );
  AOI22_X1 U158 ( .A1(B[2]), .A2(n162), .B1(E[2]), .B2(n159), .ZN(n52) );
  NAND4_X1 U159 ( .A1(n133), .A2(n134), .A3(n135), .A4(n136), .ZN(Y[10]) );
  AOI22_X1 U160 ( .A1(D[10]), .A2(n146), .B1(A[10]), .B2(n3), .ZN(n133) );
  NAND4_X1 U161 ( .A1(n129), .A2(n130), .A3(n131), .A4(n132), .ZN(Y[11]) );
  AOI22_X1 U162 ( .A1(D[11]), .A2(n146), .B1(A[11]), .B2(n3), .ZN(n129) );
  NAND4_X1 U163 ( .A1(n125), .A2(n126), .A3(n127), .A4(n128), .ZN(Y[12]) );
  AOI22_X1 U164 ( .A1(D[12]), .A2(n146), .B1(A[12]), .B2(n3), .ZN(n125) );
  NAND4_X1 U165 ( .A1(n121), .A2(n122), .A3(n123), .A4(n124), .ZN(Y[13]) );
  AOI22_X1 U166 ( .A1(D[13]), .A2(n146), .B1(A[13]), .B2(n3), .ZN(n121) );
  NAND4_X1 U167 ( .A1(n117), .A2(n118), .A3(n119), .A4(n120), .ZN(Y[14]) );
  AOI22_X1 U168 ( .A1(D[14]), .A2(n146), .B1(A[14]), .B2(n3), .ZN(n117) );
  NAND4_X1 U169 ( .A1(n105), .A2(n106), .A3(n107), .A4(n108), .ZN(Y[17]) );
  AOI22_X1 U170 ( .A1(D[17]), .A2(n145), .B1(A[17]), .B2(n2), .ZN(n105) );
  NAND4_X1 U171 ( .A1(n97), .A2(n98), .A3(n99), .A4(n100), .ZN(Y[19]) );
  AOI22_X1 U172 ( .A1(D[19]), .A2(n145), .B1(A[19]), .B2(n2), .ZN(n97) );
  NAND4_X1 U173 ( .A1(n85), .A2(n86), .A3(n87), .A4(n88), .ZN(Y[21]) );
  AOI22_X1 U174 ( .A1(D[21]), .A2(n145), .B1(A[21]), .B2(n2), .ZN(n85) );
  NAND4_X1 U175 ( .A1(n81), .A2(n82), .A3(n83), .A4(n84), .ZN(Y[22]) );
  AOI22_X1 U176 ( .A1(D[22]), .A2(n145), .B1(A[22]), .B2(n2), .ZN(n81) );
  NAND4_X1 U177 ( .A1(n77), .A2(n78), .A3(n79), .A4(n80), .ZN(Y[23]) );
  AOI22_X1 U178 ( .A1(D[23]), .A2(n145), .B1(A[23]), .B2(n2), .ZN(n77) );
  NAND4_X1 U179 ( .A1(n65), .A2(n66), .A3(n67), .A4(n68), .ZN(Y[26]) );
  AOI22_X1 U180 ( .A1(D[26]), .A2(n145), .B1(A[26]), .B2(n2), .ZN(n65) );
  NAND4_X1 U181 ( .A1(n109), .A2(n110), .A3(n111), .A4(n112), .ZN(Y[16]) );
  AOI22_X1 U182 ( .A1(D[16]), .A2(n145), .B1(A[16]), .B2(n2), .ZN(n109) );
  NAND4_X1 U183 ( .A1(n61), .A2(n62), .A3(n63), .A4(n64), .ZN(Y[27]) );
  AOI22_X1 U184 ( .A1(C[27]), .A2(n150), .B1(F[27]), .B2(n147), .ZN(n62) );
  NAND4_X1 U185 ( .A1(n57), .A2(n58), .A3(n59), .A4(n60), .ZN(Y[28]) );
  AOI22_X1 U186 ( .A1(C[28]), .A2(n150), .B1(F[28]), .B2(n147), .ZN(n58) );
  NAND4_X1 U187 ( .A1(n113), .A2(n114), .A3(n115), .A4(n116), .ZN(Y[15]) );
  AOI22_X1 U188 ( .A1(D[15]), .A2(n146), .B1(A[15]), .B2(n3), .ZN(n113) );
  NAND4_X1 U189 ( .A1(n101), .A2(n102), .A3(n103), .A4(n104), .ZN(Y[18]) );
  AOI22_X1 U190 ( .A1(D[18]), .A2(n145), .B1(A[18]), .B2(n2), .ZN(n101) );
  NAND4_X1 U191 ( .A1(n89), .A2(n90), .A3(n91), .A4(n92), .ZN(Y[20]) );
  AOI22_X1 U192 ( .A1(D[20]), .A2(n145), .B1(A[20]), .B2(n2), .ZN(n89) );
  NAND4_X1 U193 ( .A1(n73), .A2(n74), .A3(n75), .A4(n76), .ZN(Y[24]) );
  AOI22_X1 U194 ( .A1(D[24]), .A2(n145), .B1(A[24]), .B2(n2), .ZN(n73) );
  NAND4_X1 U195 ( .A1(n69), .A2(n70), .A3(n71), .A4(n72), .ZN(Y[25]) );
  AOI22_X1 U196 ( .A1(D[25]), .A2(n145), .B1(A[25]), .B2(n2), .ZN(n69) );
endmodule


module MUX41_GEN_N39 ( A, B, C, D, SEL, Y );
  input [38:0] A;
  input [38:0] B;
  input [38:0] C;
  input [38:0] D;
  input [1:0] SEL;
  output [38:0] Y;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n1, n2,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98;

  NAND2_X1 U84 ( .A1(n3), .A2(n4), .ZN(Y[9]) );
  NAND2_X1 U85 ( .A1(n9), .A2(n10), .ZN(Y[8]) );
  NAND2_X1 U86 ( .A1(n11), .A2(n12), .ZN(Y[7]) );
  NAND2_X1 U87 ( .A1(n13), .A2(n14), .ZN(Y[6]) );
  NAND2_X1 U88 ( .A1(n15), .A2(n16), .ZN(Y[5]) );
  NAND2_X1 U89 ( .A1(n17), .A2(n18), .ZN(Y[4]) );
  NAND2_X1 U90 ( .A1(n19), .A2(n20), .ZN(Y[3]) );
  NAND2_X1 U91 ( .A1(n21), .A2(n22), .ZN(Y[38]) );
  NAND2_X1 U92 ( .A1(n23), .A2(n24), .ZN(Y[37]) );
  NAND2_X1 U93 ( .A1(n25), .A2(n26), .ZN(Y[36]) );
  NAND2_X1 U94 ( .A1(n27), .A2(n28), .ZN(Y[35]) );
  NAND2_X1 U95 ( .A1(n29), .A2(n30), .ZN(Y[34]) );
  NAND2_X1 U96 ( .A1(n31), .A2(n32), .ZN(Y[33]) );
  NAND2_X1 U97 ( .A1(n33), .A2(n34), .ZN(Y[32]) );
  NAND2_X1 U98 ( .A1(n35), .A2(n36), .ZN(Y[31]) );
  NAND2_X1 U99 ( .A1(n37), .A2(n38), .ZN(Y[30]) );
  NAND2_X1 U100 ( .A1(n39), .A2(n40), .ZN(Y[2]) );
  NAND2_X1 U101 ( .A1(n41), .A2(n42), .ZN(Y[29]) );
  NAND2_X1 U102 ( .A1(n43), .A2(n44), .ZN(Y[28]) );
  NAND2_X1 U103 ( .A1(n45), .A2(n46), .ZN(Y[27]) );
  NAND2_X1 U104 ( .A1(n47), .A2(n48), .ZN(Y[26]) );
  NAND2_X1 U105 ( .A1(n49), .A2(n50), .ZN(Y[25]) );
  NAND2_X1 U106 ( .A1(n51), .A2(n52), .ZN(Y[24]) );
  NAND2_X1 U107 ( .A1(n53), .A2(n54), .ZN(Y[23]) );
  NAND2_X1 U108 ( .A1(n55), .A2(n56), .ZN(Y[22]) );
  NAND2_X1 U109 ( .A1(n57), .A2(n58), .ZN(Y[21]) );
  NAND2_X1 U110 ( .A1(n59), .A2(n60), .ZN(Y[20]) );
  NAND2_X1 U111 ( .A1(n61), .A2(n62), .ZN(Y[1]) );
  NAND2_X1 U112 ( .A1(n63), .A2(n64), .ZN(Y[19]) );
  NAND2_X1 U113 ( .A1(n65), .A2(n66), .ZN(Y[18]) );
  NAND2_X1 U114 ( .A1(n67), .A2(n68), .ZN(Y[17]) );
  NAND2_X1 U115 ( .A1(n69), .A2(n70), .ZN(Y[16]) );
  NAND2_X1 U116 ( .A1(n71), .A2(n72), .ZN(Y[15]) );
  NAND2_X1 U117 ( .A1(n73), .A2(n74), .ZN(Y[14]) );
  NAND2_X1 U118 ( .A1(n75), .A2(n76), .ZN(Y[13]) );
  NAND2_X1 U119 ( .A1(n77), .A2(n78), .ZN(Y[12]) );
  NAND2_X1 U120 ( .A1(n79), .A2(n80), .ZN(Y[11]) );
  NAND2_X1 U121 ( .A1(n81), .A2(n82), .ZN(Y[10]) );
  NAND2_X1 U122 ( .A1(n83), .A2(n84), .ZN(Y[0]) );
  BUF_X1 U1 ( .A(n7), .Z(n90) );
  BUF_X1 U2 ( .A(n7), .Z(n91) );
  BUF_X1 U3 ( .A(n7), .Z(n92) );
  AOI22_X1 U4 ( .A1(B[38]), .A2(n96), .B1(C[38]), .B2(n93), .ZN(n22) );
  AOI22_X1 U5 ( .A1(D[38]), .A2(n92), .B1(A[38]), .B2(n87), .ZN(n21) );
  AOI22_X1 U6 ( .A1(B[31]), .A2(n97), .B1(C[31]), .B2(n94), .ZN(n36) );
  AOI22_X1 U7 ( .A1(D[31]), .A2(n91), .B1(A[31]), .B2(n88), .ZN(n35) );
  AOI22_X1 U8 ( .A1(B[32]), .A2(n97), .B1(C[32]), .B2(n94), .ZN(n34) );
  AOI22_X1 U9 ( .A1(D[32]), .A2(n91), .B1(A[32]), .B2(n88), .ZN(n33) );
  AND3_X1 U10 ( .A1(n1), .A2(n2), .A3(n86), .ZN(n7) );
  INV_X1 U11 ( .A(n6), .ZN(n1) );
  INV_X1 U12 ( .A(n8), .ZN(n2) );
  INV_X1 U13 ( .A(n5), .ZN(n86) );
  AOI22_X1 U14 ( .A1(B[33]), .A2(n96), .B1(C[33]), .B2(n93), .ZN(n32) );
  AOI22_X1 U15 ( .A1(D[33]), .A2(n92), .B1(A[33]), .B2(n87), .ZN(n31) );
  AOI22_X1 U16 ( .A1(B[34]), .A2(n96), .B1(C[34]), .B2(n93), .ZN(n30) );
  AOI22_X1 U17 ( .A1(D[34]), .A2(n92), .B1(A[34]), .B2(n87), .ZN(n29) );
  AOI22_X1 U18 ( .A1(B[35]), .A2(n96), .B1(C[35]), .B2(n93), .ZN(n28) );
  AOI22_X1 U19 ( .A1(D[35]), .A2(n92), .B1(A[35]), .B2(n87), .ZN(n27) );
  AOI22_X1 U20 ( .A1(B[36]), .A2(n96), .B1(C[36]), .B2(n93), .ZN(n26) );
  AOI22_X1 U21 ( .A1(D[36]), .A2(n92), .B1(A[36]), .B2(n87), .ZN(n25) );
  AOI22_X1 U22 ( .A1(B[37]), .A2(n96), .B1(C[37]), .B2(n93), .ZN(n24) );
  AOI22_X1 U23 ( .A1(D[37]), .A2(n92), .B1(A[37]), .B2(n87), .ZN(n23) );
  BUF_X1 U24 ( .A(n6), .Z(n95) );
  BUF_X1 U25 ( .A(n6), .Z(n94) );
  BUF_X1 U26 ( .A(n6), .Z(n93) );
  BUF_X1 U27 ( .A(n5), .Z(n98) );
  BUF_X1 U28 ( .A(n5), .Z(n97) );
  BUF_X1 U29 ( .A(n5), .Z(n96) );
  BUF_X1 U30 ( .A(n8), .Z(n89) );
  BUF_X1 U31 ( .A(n8), .Z(n88) );
  BUF_X1 U32 ( .A(n8), .Z(n87) );
  AOI22_X1 U33 ( .A1(B[7]), .A2(n96), .B1(C[7]), .B2(n93), .ZN(n12) );
  AOI22_X1 U34 ( .A1(D[7]), .A2(n92), .B1(A[7]), .B2(n87), .ZN(n11) );
  AOI22_X1 U35 ( .A1(B[8]), .A2(n96), .B1(C[8]), .B2(n93), .ZN(n10) );
  AOI22_X1 U36 ( .A1(D[8]), .A2(n92), .B1(A[8]), .B2(n87), .ZN(n9) );
  AOI22_X1 U37 ( .A1(B[9]), .A2(n96), .B1(C[9]), .B2(n93), .ZN(n4) );
  AOI22_X1 U38 ( .A1(D[9]), .A2(n92), .B1(A[9]), .B2(n87), .ZN(n3) );
  AOI22_X1 U39 ( .A1(B[10]), .A2(n98), .B1(C[10]), .B2(n95), .ZN(n82) );
  AOI22_X1 U40 ( .A1(D[10]), .A2(n90), .B1(A[10]), .B2(n89), .ZN(n81) );
  AOI22_X1 U41 ( .A1(B[11]), .A2(n98), .B1(C[11]), .B2(n95), .ZN(n80) );
  AOI22_X1 U42 ( .A1(D[11]), .A2(n90), .B1(A[11]), .B2(n89), .ZN(n79) );
  AOI22_X1 U43 ( .A1(B[12]), .A2(n98), .B1(C[12]), .B2(n95), .ZN(n78) );
  AOI22_X1 U44 ( .A1(D[12]), .A2(n90), .B1(A[12]), .B2(n89), .ZN(n77) );
  AOI22_X1 U45 ( .A1(B[13]), .A2(n98), .B1(C[13]), .B2(n95), .ZN(n76) );
  AOI22_X1 U46 ( .A1(D[13]), .A2(n90), .B1(A[13]), .B2(n89), .ZN(n75) );
  AOI22_X1 U47 ( .A1(B[14]), .A2(n98), .B1(C[14]), .B2(n95), .ZN(n74) );
  AOI22_X1 U48 ( .A1(D[14]), .A2(n90), .B1(A[14]), .B2(n89), .ZN(n73) );
  AOI22_X1 U49 ( .A1(B[15]), .A2(n98), .B1(C[15]), .B2(n95), .ZN(n72) );
  AOI22_X1 U50 ( .A1(D[15]), .A2(n90), .B1(A[15]), .B2(n89), .ZN(n71) );
  AOI22_X1 U51 ( .A1(B[16]), .A2(n98), .B1(C[16]), .B2(n95), .ZN(n70) );
  AOI22_X1 U52 ( .A1(D[16]), .A2(n90), .B1(A[16]), .B2(n89), .ZN(n69) );
  AOI22_X1 U53 ( .A1(B[17]), .A2(n98), .B1(C[17]), .B2(n95), .ZN(n68) );
  AOI22_X1 U54 ( .A1(D[17]), .A2(n90), .B1(A[17]), .B2(n89), .ZN(n67) );
  AOI22_X1 U55 ( .A1(B[18]), .A2(n98), .B1(C[18]), .B2(n95), .ZN(n66) );
  AOI22_X1 U56 ( .A1(D[18]), .A2(n90), .B1(A[18]), .B2(n89), .ZN(n65) );
  AOI22_X1 U57 ( .A1(B[19]), .A2(n98), .B1(C[19]), .B2(n95), .ZN(n64) );
  AOI22_X1 U58 ( .A1(D[19]), .A2(n90), .B1(A[19]), .B2(n89), .ZN(n63) );
  AOI22_X1 U59 ( .A1(B[20]), .A2(n98), .B1(C[20]), .B2(n95), .ZN(n60) );
  AOI22_X1 U60 ( .A1(D[20]), .A2(n90), .B1(A[20]), .B2(n89), .ZN(n59) );
  AOI22_X1 U61 ( .A1(B[21]), .A2(n97), .B1(C[21]), .B2(n94), .ZN(n58) );
  AOI22_X1 U62 ( .A1(D[21]), .A2(n91), .B1(A[21]), .B2(n88), .ZN(n57) );
  AOI22_X1 U63 ( .A1(B[22]), .A2(n97), .B1(C[22]), .B2(n94), .ZN(n56) );
  AOI22_X1 U64 ( .A1(D[22]), .A2(n91), .B1(A[22]), .B2(n88), .ZN(n55) );
  AOI22_X1 U65 ( .A1(B[23]), .A2(n97), .B1(C[23]), .B2(n94), .ZN(n54) );
  AOI22_X1 U66 ( .A1(D[23]), .A2(n91), .B1(A[23]), .B2(n88), .ZN(n53) );
  AOI22_X1 U67 ( .A1(B[24]), .A2(n97), .B1(C[24]), .B2(n94), .ZN(n52) );
  AOI22_X1 U68 ( .A1(D[24]), .A2(n91), .B1(A[24]), .B2(n88), .ZN(n51) );
  AOI22_X1 U69 ( .A1(B[25]), .A2(n97), .B1(C[25]), .B2(n94), .ZN(n50) );
  AOI22_X1 U70 ( .A1(D[25]), .A2(n91), .B1(A[25]), .B2(n88), .ZN(n49) );
  AOI22_X1 U71 ( .A1(B[26]), .A2(n97), .B1(C[26]), .B2(n94), .ZN(n48) );
  AOI22_X1 U72 ( .A1(D[26]), .A2(n91), .B1(A[26]), .B2(n88), .ZN(n47) );
  AOI22_X1 U73 ( .A1(B[27]), .A2(n97), .B1(C[27]), .B2(n94), .ZN(n46) );
  AOI22_X1 U74 ( .A1(D[27]), .A2(n91), .B1(A[27]), .B2(n88), .ZN(n45) );
  AOI22_X1 U75 ( .A1(B[28]), .A2(n97), .B1(C[28]), .B2(n94), .ZN(n44) );
  AOI22_X1 U76 ( .A1(D[28]), .A2(n91), .B1(A[28]), .B2(n88), .ZN(n43) );
  AOI22_X1 U77 ( .A1(B[29]), .A2(n97), .B1(C[29]), .B2(n94), .ZN(n42) );
  AOI22_X1 U78 ( .A1(D[29]), .A2(n91), .B1(A[29]), .B2(n88), .ZN(n41) );
  AOI22_X1 U79 ( .A1(B[30]), .A2(n97), .B1(C[30]), .B2(n94), .ZN(n38) );
  AOI22_X1 U80 ( .A1(D[30]), .A2(n91), .B1(A[30]), .B2(n88), .ZN(n37) );
  NOR2_X1 U81 ( .A1(n85), .A2(SEL[1]), .ZN(n6) );
  AOI22_X1 U82 ( .A1(B[6]), .A2(n96), .B1(C[6]), .B2(n93), .ZN(n14) );
  AOI22_X1 U83 ( .A1(D[6]), .A2(n92), .B1(A[6]), .B2(n87), .ZN(n13) );
  AOI22_X1 U123 ( .A1(B[5]), .A2(n96), .B1(C[5]), .B2(n93), .ZN(n16) );
  AOI22_X1 U124 ( .A1(D[5]), .A2(n92), .B1(A[5]), .B2(n87), .ZN(n15) );
  AOI22_X1 U125 ( .A1(B[4]), .A2(n96), .B1(C[4]), .B2(n93), .ZN(n18) );
  AOI22_X1 U126 ( .A1(D[4]), .A2(n92), .B1(A[4]), .B2(n87), .ZN(n17) );
  AOI22_X1 U127 ( .A1(B[3]), .A2(n96), .B1(C[3]), .B2(n93), .ZN(n20) );
  AOI22_X1 U128 ( .A1(D[3]), .A2(n92), .B1(A[3]), .B2(n87), .ZN(n19) );
  AND2_X1 U129 ( .A1(SEL[0]), .A2(SEL[1]), .ZN(n8) );
  AND2_X1 U130 ( .A1(SEL[1]), .A2(n85), .ZN(n5) );
  AOI22_X1 U131 ( .A1(B[2]), .A2(n97), .B1(C[2]), .B2(n94), .ZN(n40) );
  AOI22_X1 U132 ( .A1(D[2]), .A2(n91), .B1(A[2]), .B2(n88), .ZN(n39) );
  INV_X1 U133 ( .A(SEL[0]), .ZN(n85) );
  AOI22_X1 U134 ( .A1(B[1]), .A2(n98), .B1(C[1]), .B2(n95), .ZN(n62) );
  AOI22_X1 U135 ( .A1(D[1]), .A2(n90), .B1(A[1]), .B2(n89), .ZN(n61) );
  AOI22_X1 U136 ( .A1(B[0]), .A2(n98), .B1(C[0]), .B2(n95), .ZN(n84) );
  AOI22_X1 U137 ( .A1(D[0]), .A2(n90), .B1(A[0]), .B2(n89), .ZN(n83) );
endmodule


module MUX21_GEN_N7_0 ( A, B, SEL, Y );
  input [6:0] A;
  input [6:0] B;
  output [6:0] Y;
  input SEL;
  wire   SB;
  wire   [6:0] Y1;
  wire   [6:0] Y2;

  INV_1_27 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_612 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_611 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_610 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_609 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_608 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_607 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_606 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_605 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_604 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_603 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_602 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_601 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_600 UND1_4 ( .A(A[4]), .B(SEL), .Y(Y1[4]) );
  NAND_GATE_599 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  NAND_GATE_598 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_597 UND1_5 ( .A(A[5]), .B(SEL), .Y(Y1[5]) );
  NAND_GATE_596 UND2_5 ( .A(B[5]), .B(SB), .Y(Y2[5]) );
  NAND_GATE_595 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_594 UND1_6 ( .A(A[6]), .B(SEL), .Y(Y1[6]) );
  NAND_GATE_593 UND2_6 ( .A(B[6]), .B(SB), .Y(Y2[6]) );
  NAND_GATE_592 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
endmodule


module MUX21_GEN_N8_0 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;
  wire   SB;
  wire   [7:0] Y1;
  wire   [7:0] Y2;

  INV_1_31 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_708 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_707 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_706 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_705 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_704 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_703 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_702 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_701 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_700 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_699 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_698 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_697 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_696 UND1_4 ( .A(A[4]), .B(SEL), .Y(Y1[4]) );
  NAND_GATE_695 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  NAND_GATE_694 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_693 UND1_5 ( .A(A[5]), .B(SEL), .Y(Y1[5]) );
  NAND_GATE_692 UND2_5 ( .A(B[5]), .B(SB), .Y(Y2[5]) );
  NAND_GATE_691 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_690 UND1_6 ( .A(A[6]), .B(SEL), .Y(Y1[6]) );
  NAND_GATE_689 UND2_6 ( .A(B[6]), .B(SB), .Y(Y2[6]) );
  NAND_GATE_688 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_687 UND1_7 ( .A(A[7]), .B(SEL), .Y(Y1[7]) );
  NAND_GATE_686 UND2_7 ( .A(B[7]), .B(SB), .Y(Y2[7]) );
  NAND_GATE_685 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
endmodule


module N_NAND_N4_0 ( A, Y );
  input [3:0] A;
  output Y;


  NAND4_X1 U1 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module N_NAND_N3_0 ( A, Y );
  input [2:0] A;
  output Y;


  NAND3_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(Y) );
endmodule


module MUX61 ( A, B, C, D, E, F, SEL, Y );
  input [2:0] SEL;
  input A, B, C, D, E, F;
  output Y;
  wire   n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19;

  NAND2_X1 U12 ( .A1(A), .A2(n6), .ZN(n8) );
  NAND2_X1 U13 ( .A1(SEL[2]), .A2(SEL[1]), .ZN(n10) );
  NAND2_X1 U14 ( .A1(C), .A2(n12), .ZN(n14) );
  NAND2_X1 U15 ( .A1(SEL[1]), .A2(SEL[0]), .ZN(n19) );
  AOI22_X1 U1 ( .A1(n15), .A2(n16), .B1(D), .B2(SEL[2]), .ZN(n13) );
  AND2_X1 U2 ( .A1(SEL[2]), .A2(SEL[0]), .ZN(n12) );
  AOI22_X1 U3 ( .A1(n9), .A2(n10), .B1(B), .B2(n11), .ZN(n7) );
  INV_X1 U4 ( .A(n10), .ZN(n11) );
  INV_X1 U5 ( .A(n17), .ZN(n15) );
  INV_X1 U6 ( .A(n19), .ZN(n18) );
  INV_X1 U7 ( .A(SEL[2]), .ZN(n16) );
  AND3_X1 U8 ( .A1(SEL[1]), .A2(SEL[0]), .A3(SEL[2]), .ZN(n6) );
  OAI21_X1 U9 ( .B1(n6), .B2(n7), .A(n8), .ZN(Y) );
  OAI21_X1 U10 ( .B1(n12), .B2(n13), .A(n14), .ZN(n9) );
  AOI22_X1 U11 ( .A1(E), .A2(n18), .B1(F), .B2(n19), .ZN(n17) );
endmodule


module N_NOR_N32 ( A, Y );
  input [31:0] A;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  NOR4_X1 U1 ( .A1(A[9]), .A2(A[8]), .A3(A[7]), .A4(A[6]), .ZN(n10) );
  NOR4_X1 U2 ( .A1(A[5]), .A2(A[4]), .A3(A[3]), .A4(A[31]), .ZN(n9) );
  NOR4_X1 U3 ( .A1(A[30]), .A2(A[2]), .A3(A[29]), .A4(A[28]), .ZN(n8) );
  NOR4_X1 U4 ( .A1(A[27]), .A2(A[26]), .A3(A[25]), .A4(A[24]), .ZN(n7) );
  NOR4_X1 U5 ( .A1(A[23]), .A2(A[22]), .A3(A[21]), .A4(A[20]), .ZN(n6) );
  NOR4_X1 U6 ( .A1(A[1]), .A2(A[19]), .A3(A[18]), .A4(A[17]), .ZN(n5) );
  NOR4_X1 U7 ( .A1(A[16]), .A2(A[15]), .A3(A[14]), .A4(A[13]), .ZN(n4) );
  NOR2_X1 U8 ( .A1(n1), .A2(n2), .ZN(Y) );
  NAND4_X1 U9 ( .A1(n7), .A2(n8), .A3(n9), .A4(n10), .ZN(n1) );
  NOR4_X1 U10 ( .A1(A[12]), .A2(A[11]), .A3(A[10]), .A4(A[0]), .ZN(n3) );
  NAND4_X1 U11 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(n2) );
endmodule


module SUM_GENERATOR_N32 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  CSA_N4_8 DO_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0]) );
  CSA_N4_7 DO_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4]) );
  CSA_N4_6 DO_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  CSA_N4_5 DO_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(S[15:12]) );
  CSA_N4_4 DO_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(S[19:16]) );
  CSA_N4_3 DO_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(S[23:20]) );
  CSA_N4_2 DO_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(S[27:24]) );
  CSA_N4_1 DO_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(S[31:28]) );
endmodule


module CARRY_GENERATOR_N32 ( A, B, Ci, Co );
  input [31:0] A;
  input [31:0] B;
  output [7:0] Co;
  input Ci;
  wire   \pro_signal[4][7] , \pro_signal[4][6] , \pro_signal[3][7] ,
         \pro_signal[3][5] , \pro_signal[3][3] , \pro_signal[3][2] ,
         \pro_signal[2][7] , \pro_signal[2][6] , \pro_signal[2][5] ,
         \pro_signal[2][4] , \pro_signal[2][3] , \pro_signal[2][1] ,
         \pro_signal[1][15] , \pro_signal[1][14] , \pro_signal[1][13] ,
         \pro_signal[1][12] , \pro_signal[1][11] , \pro_signal[1][10] ,
         \pro_signal[1][9] , \pro_signal[1][8] , \pro_signal[1][7] ,
         \pro_signal[1][6] , \pro_signal[1][5] , \pro_signal[1][4] ,
         \pro_signal[1][3] , \pro_signal[1][2] , \pro_signal[1][1] ,
         \pro_signal[0][31] , \pro_signal[0][30] , \pro_signal[0][29] ,
         \pro_signal[0][28] , \pro_signal[0][27] , \pro_signal[0][26] ,
         \pro_signal[0][25] , \pro_signal[0][24] , \pro_signal[0][23] ,
         \pro_signal[0][22] , \pro_signal[0][21] , \pro_signal[0][20] ,
         \pro_signal[0][19] , \pro_signal[0][18] , \pro_signal[0][17] ,
         \pro_signal[0][16] , \pro_signal[0][15] , \pro_signal[0][14] ,
         \pro_signal[0][13] , \pro_signal[0][12] , \pro_signal[0][11] ,
         \pro_signal[0][10] , \pro_signal[0][9] , \pro_signal[0][8] ,
         \pro_signal[0][7] , \pro_signal[0][6] , \pro_signal[0][5] ,
         \pro_signal[0][4] , \pro_signal[0][3] , \pro_signal[0][2] ,
         \pro_signal[0][1] , \gen_signal[4][7] , \gen_signal[4][6] ,
         \gen_signal[3][7] , \gen_signal[3][5] , \gen_signal[3][3] ,
         \gen_signal[2][7] , \gen_signal[2][6] , \gen_signal[2][5] ,
         \gen_signal[2][4] , \gen_signal[2][3] , \gen_signal[2][2] ,
         \gen_signal[2][1] , \gen_signal[1][15] , \gen_signal[1][14] ,
         \gen_signal[1][13] , \gen_signal[1][12] , \gen_signal[1][11] ,
         \gen_signal[1][10] , \gen_signal[1][9] , \gen_signal[1][8] ,
         \gen_signal[1][7] , \gen_signal[1][6] , \gen_signal[1][5] ,
         \gen_signal[1][4] , \gen_signal[1][3] , \gen_signal[1][2] ,
         \gen_signal[1][1] , \gen_signal[1][0] , \gen_signal[0][31] ,
         \gen_signal[0][30] , \gen_signal[0][29] , \gen_signal[0][28] ,
         \gen_signal[0][27] , \gen_signal[0][26] , \gen_signal[0][25] ,
         \gen_signal[0][24] , \gen_signal[0][23] , \gen_signal[0][22] ,
         \gen_signal[0][21] , \gen_signal[0][20] , \gen_signal[0][19] ,
         \gen_signal[0][18] , \gen_signal[0][17] , \gen_signal[0][16] ,
         \gen_signal[0][15] , \gen_signal[0][14] , \gen_signal[0][13] ,
         \gen_signal[0][12] , \gen_signal[0][11] , \gen_signal[0][10] ,
         \gen_signal[0][9] , \gen_signal[0][8] , \gen_signal[0][7] ,
         \gen_signal[0][6] , \gen_signal[0][5] , \gen_signal[0][4] ,
         \gen_signal[0][3] , \gen_signal[0][2] , \gen_signal[0][1] ,
         \gen_signal[0][0] ;
  wire   SYNOPSYS_UNCONNECTED__0;

  PG_NETWORK_N32 PG_NETWORK_INST ( .A(A), .B(B), .Ci(Ci), .G({
        \gen_signal[0][31] , \gen_signal[0][30] , \gen_signal[0][29] , 
        \gen_signal[0][28] , \gen_signal[0][27] , \gen_signal[0][26] , 
        \gen_signal[0][25] , \gen_signal[0][24] , \gen_signal[0][23] , 
        \gen_signal[0][22] , \gen_signal[0][21] , \gen_signal[0][20] , 
        \gen_signal[0][19] , \gen_signal[0][18] , \gen_signal[0][17] , 
        \gen_signal[0][16] , \gen_signal[0][15] , \gen_signal[0][14] , 
        \gen_signal[0][13] , \gen_signal[0][12] , \gen_signal[0][11] , 
        \gen_signal[0][10] , \gen_signal[0][9] , \gen_signal[0][8] , 
        \gen_signal[0][7] , \gen_signal[0][6] , \gen_signal[0][5] , 
        \gen_signal[0][4] , \gen_signal[0][3] , \gen_signal[0][2] , 
        \gen_signal[0][1] , \gen_signal[0][0] }), .P({\pro_signal[0][31] , 
        \pro_signal[0][30] , \pro_signal[0][29] , \pro_signal[0][28] , 
        \pro_signal[0][27] , \pro_signal[0][26] , \pro_signal[0][25] , 
        \pro_signal[0][24] , \pro_signal[0][23] , \pro_signal[0][22] , 
        \pro_signal[0][21] , \pro_signal[0][20] , \pro_signal[0][19] , 
        \pro_signal[0][18] , \pro_signal[0][17] , \pro_signal[0][16] , 
        \pro_signal[0][15] , \pro_signal[0][14] , \pro_signal[0][13] , 
        \pro_signal[0][12] , \pro_signal[0][11] , \pro_signal[0][10] , 
        \pro_signal[0][9] , \pro_signal[0][8] , \pro_signal[0][7] , 
        \pro_signal[0][6] , \pro_signal[0][5] , \pro_signal[0][4] , 
        \pro_signal[0][3] , \pro_signal[0][2] , \pro_signal[0][1] , 
        SYNOPSYS_UNCONNECTED__0}) );
  GENERAL_GENERATE_0 G_INST_1_0_0 ( .Gi_0(\gen_signal[0][0] ), .Gi_1(
        \gen_signal[0][1] ), .Pi(\pro_signal[0][1] ), .Go(\gen_signal[1][0] )
         );
  PG_BLOCK_0 PG_INST_1_0_1 ( .Gi_0(\gen_signal[0][2] ), .Gi_1(
        \gen_signal[0][3] ), .Pi_0(\pro_signal[0][2] ), .Pi_1(
        \pro_signal[0][3] ), .Po(\pro_signal[1][1] ), .Go(\gen_signal[1][1] )
         );
  PG_BLOCK_26 PG_INST_1_0_2 ( .Gi_0(\gen_signal[0][4] ), .Gi_1(
        \gen_signal[0][5] ), .Pi_0(\pro_signal[0][4] ), .Pi_1(
        \pro_signal[0][5] ), .Po(\pro_signal[1][2] ), .Go(\gen_signal[1][2] )
         );
  PG_BLOCK_25 PG_INST_1_0_3 ( .Gi_0(\gen_signal[0][6] ), .Gi_1(
        \gen_signal[0][7] ), .Pi_0(\pro_signal[0][6] ), .Pi_1(
        \pro_signal[0][7] ), .Po(\pro_signal[1][3] ), .Go(\gen_signal[1][3] )
         );
  PG_BLOCK_24 PG_INST_1_0_4 ( .Gi_0(\gen_signal[0][8] ), .Gi_1(
        \gen_signal[0][9] ), .Pi_0(\pro_signal[0][8] ), .Pi_1(
        \pro_signal[0][9] ), .Po(\pro_signal[1][4] ), .Go(\gen_signal[1][4] )
         );
  PG_BLOCK_23 PG_INST_1_0_5 ( .Gi_0(\gen_signal[0][10] ), .Gi_1(
        \gen_signal[0][11] ), .Pi_0(\pro_signal[0][10] ), .Pi_1(
        \pro_signal[0][11] ), .Po(\pro_signal[1][5] ), .Go(\gen_signal[1][5] )
         );
  PG_BLOCK_22 PG_INST_1_0_6 ( .Gi_0(\gen_signal[0][12] ), .Gi_1(
        \gen_signal[0][13] ), .Pi_0(\pro_signal[0][12] ), .Pi_1(
        \pro_signal[0][13] ), .Po(\pro_signal[1][6] ), .Go(\gen_signal[1][6] )
         );
  PG_BLOCK_21 PG_INST_1_0_7 ( .Gi_0(\gen_signal[0][14] ), .Gi_1(
        \gen_signal[0][15] ), .Pi_0(\pro_signal[0][14] ), .Pi_1(
        \pro_signal[0][15] ), .Po(\pro_signal[1][7] ), .Go(\gen_signal[1][7] )
         );
  PG_BLOCK_20 PG_INST_1_0_8 ( .Gi_0(\gen_signal[0][16] ), .Gi_1(
        \gen_signal[0][17] ), .Pi_0(\pro_signal[0][16] ), .Pi_1(
        \pro_signal[0][17] ), .Po(\pro_signal[1][8] ), .Go(\gen_signal[1][8] )
         );
  PG_BLOCK_19 PG_INST_1_0_9 ( .Gi_0(\gen_signal[0][18] ), .Gi_1(
        \gen_signal[0][19] ), .Pi_0(\pro_signal[0][18] ), .Pi_1(
        \pro_signal[0][19] ), .Po(\pro_signal[1][9] ), .Go(\gen_signal[1][9] )
         );
  PG_BLOCK_18 PG_INST_1_0_10 ( .Gi_0(\gen_signal[0][20] ), .Gi_1(
        \gen_signal[0][21] ), .Pi_0(\pro_signal[0][20] ), .Pi_1(
        \pro_signal[0][21] ), .Po(\pro_signal[1][10] ), .Go(
        \gen_signal[1][10] ) );
  PG_BLOCK_17 PG_INST_1_0_11 ( .Gi_0(\gen_signal[0][22] ), .Gi_1(
        \gen_signal[0][23] ), .Pi_0(\pro_signal[0][22] ), .Pi_1(
        \pro_signal[0][23] ), .Po(\pro_signal[1][11] ), .Go(
        \gen_signal[1][11] ) );
  PG_BLOCK_16 PG_INST_1_0_12 ( .Gi_0(\gen_signal[0][24] ), .Gi_1(
        \gen_signal[0][25] ), .Pi_0(\pro_signal[0][24] ), .Pi_1(
        \pro_signal[0][25] ), .Po(\pro_signal[1][12] ), .Go(
        \gen_signal[1][12] ) );
  PG_BLOCK_15 PG_INST_1_0_13 ( .Gi_0(\gen_signal[0][26] ), .Gi_1(
        \gen_signal[0][27] ), .Pi_0(\pro_signal[0][26] ), .Pi_1(
        \pro_signal[0][27] ), .Po(\pro_signal[1][13] ), .Go(
        \gen_signal[1][13] ) );
  PG_BLOCK_14 PG_INST_1_0_14 ( .Gi_0(\gen_signal[0][28] ), .Gi_1(
        \gen_signal[0][29] ), .Pi_0(\pro_signal[0][28] ), .Pi_1(
        \pro_signal[0][29] ), .Po(\pro_signal[1][14] ), .Go(
        \gen_signal[1][14] ) );
  PG_BLOCK_13 PG_INST_1_0_15 ( .Gi_0(\gen_signal[0][30] ), .Gi_1(
        \gen_signal[0][31] ), .Pi_0(\pro_signal[0][30] ), .Pi_1(
        \pro_signal[0][31] ), .Po(\pro_signal[1][15] ), .Go(
        \gen_signal[1][15] ) );
  GENERAL_GENERATE_36 G_INST_1_1_0 ( .Gi_0(\gen_signal[1][0] ), .Gi_1(
        \gen_signal[1][1] ), .Pi(\pro_signal[1][1] ), .Go(Co[0]) );
  PG_BLOCK_12 PG_INST_1_1_1 ( .Gi_0(\gen_signal[1][2] ), .Gi_1(
        \gen_signal[1][3] ), .Pi_0(\pro_signal[1][2] ), .Pi_1(
        \pro_signal[1][3] ), .Po(\pro_signal[2][1] ), .Go(\gen_signal[2][1] )
         );
  PG_BLOCK_11 PG_INST_1_1_2 ( .Gi_0(\gen_signal[1][4] ), .Gi_1(
        \gen_signal[1][5] ), .Pi_0(\pro_signal[1][4] ), .Pi_1(
        \pro_signal[1][5] ), .Po(\pro_signal[3][2] ), .Go(\gen_signal[2][2] )
         );
  PG_BLOCK_10 PG_INST_1_1_3 ( .Gi_0(\gen_signal[1][6] ), .Gi_1(
        \gen_signal[1][7] ), .Pi_0(\pro_signal[1][6] ), .Pi_1(
        \pro_signal[1][7] ), .Po(\pro_signal[2][3] ), .Go(\gen_signal[2][3] )
         );
  PG_BLOCK_9 PG_INST_1_1_4 ( .Gi_0(\gen_signal[1][8] ), .Gi_1(
        \gen_signal[1][9] ), .Pi_0(\pro_signal[1][8] ), .Pi_1(
        \pro_signal[1][9] ), .Po(\pro_signal[2][4] ), .Go(\gen_signal[2][4] )
         );
  PG_BLOCK_8 PG_INST_1_1_5 ( .Gi_0(\gen_signal[1][10] ), .Gi_1(
        \gen_signal[1][11] ), .Pi_0(\pro_signal[1][10] ), .Pi_1(
        \pro_signal[1][11] ), .Po(\pro_signal[2][5] ), .Go(\gen_signal[2][5] )
         );
  PG_BLOCK_7 PG_INST_1_1_6 ( .Gi_0(\gen_signal[1][12] ), .Gi_1(
        \gen_signal[1][13] ), .Pi_0(\pro_signal[1][12] ), .Pi_1(
        \pro_signal[1][13] ), .Po(\pro_signal[2][6] ), .Go(\gen_signal[2][6] )
         );
  PG_BLOCK_6 PG_INST_1_1_7 ( .Gi_0(\gen_signal[1][14] ), .Gi_1(
        \gen_signal[1][15] ), .Pi_0(\pro_signal[1][14] ), .Pi_1(
        \pro_signal[1][15] ), .Po(\pro_signal[2][7] ), .Go(\gen_signal[2][7] )
         );
  GENERAL_GENERATE_35 G_INST_2_2_0_1 ( .Gi_0(Co[0]), .Gi_1(\gen_signal[2][1] ), 
        .Pi(\pro_signal[2][1] ), .Go(Co[1]) );
  PG_BLOCK_5 PG_INST_2_2_1_1 ( .Gi_0(\gen_signal[2][2] ), .Gi_1(
        \gen_signal[2][3] ), .Pi_0(\pro_signal[3][2] ), .Pi_1(
        \pro_signal[2][3] ), .Po(\pro_signal[3][3] ), .Go(\gen_signal[3][3] )
         );
  PG_BLOCK_4 PG_INST_2_2_2_1 ( .Gi_0(\gen_signal[2][4] ), .Gi_1(
        \gen_signal[2][5] ), .Pi_0(\pro_signal[2][4] ), .Pi_1(
        \pro_signal[2][5] ), .Po(\pro_signal[3][5] ), .Go(\gen_signal[3][5] )
         );
  PG_BLOCK_3 PG_INST_2_2_3_1 ( .Gi_0(\gen_signal[2][6] ), .Gi_1(
        \gen_signal[2][7] ), .Pi_0(\pro_signal[2][6] ), .Pi_1(
        \pro_signal[2][7] ), .Po(\pro_signal[3][7] ), .Go(\gen_signal[3][7] )
         );
  GENERAL_GENERATE_34 G_INST_2_3_0_2 ( .Gi_0(Co[1]), .Gi_1(\gen_signal[2][2] ), 
        .Pi(\pro_signal[3][2] ), .Go(Co[2]) );
  GENERAL_GENERATE_33 G_INST_2_3_0_3 ( .Gi_0(Co[1]), .Gi_1(\gen_signal[3][3] ), 
        .Pi(\pro_signal[3][3] ), .Go(Co[3]) );
  PG_BLOCK_2 PG_INST_2_3_1_2 ( .Gi_0(\gen_signal[3][5] ), .Gi_1(
        \gen_signal[2][6] ), .Pi_0(\pro_signal[3][5] ), .Pi_1(
        \pro_signal[2][6] ), .Po(\pro_signal[4][6] ), .Go(\gen_signal[4][6] )
         );
  PG_BLOCK_1 PG_INST_2_3_1_3 ( .Gi_0(\gen_signal[3][5] ), .Gi_1(
        \gen_signal[3][7] ), .Pi_0(\pro_signal[3][5] ), .Pi_1(
        \pro_signal[3][7] ), .Po(\pro_signal[4][7] ), .Go(\gen_signal[4][7] )
         );
  GENERAL_GENERATE_32 G_INST_2_4_0_4 ( .Gi_0(Co[3]), .Gi_1(\gen_signal[2][4] ), 
        .Pi(\pro_signal[2][4] ), .Go(Co[4]) );
  GENERAL_GENERATE_31 G_INST_2_4_0_5 ( .Gi_0(Co[3]), .Gi_1(\gen_signal[3][5] ), 
        .Pi(\pro_signal[3][5] ), .Go(Co[5]) );
  GENERAL_GENERATE_30 G_INST_2_4_0_6 ( .Gi_0(Co[3]), .Gi_1(\gen_signal[4][6] ), 
        .Pi(\pro_signal[4][6] ), .Go(Co[6]) );
  GENERAL_GENERATE_29 G_INST_2_4_0_7 ( .Gi_0(Co[3]), .Gi_1(\gen_signal[4][7] ), 
        .Pi(\pro_signal[4][7] ), .Go(Co[7]) );
endmodule


module NOR_GATE_0 ( A, B, Y );
  input A, B;
  output Y;


  NOR2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module N_AND_N32_0 ( A, Y );
  input [31:0] A;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  NOR4_X1 U1 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(n2) );
  NAND4_X1 U2 ( .A1(A[12]), .A2(A[11]), .A3(A[10]), .A4(A[0]), .ZN(n3) );
  NAND4_X1 U3 ( .A1(A[16]), .A2(A[15]), .A3(A[14]), .A4(A[13]), .ZN(n4) );
  NAND4_X1 U4 ( .A1(A[1]), .A2(A[19]), .A3(A[18]), .A4(A[17]), .ZN(n5) );
  AND2_X1 U5 ( .A1(n1), .A2(n2), .ZN(Y) );
  NOR4_X1 U6 ( .A1(n7), .A2(n8), .A3(n9), .A4(n10), .ZN(n1) );
  NAND4_X1 U7 ( .A1(A[23]), .A2(A[22]), .A3(A[21]), .A4(A[20]), .ZN(n6) );
  NAND4_X1 U8 ( .A1(A[9]), .A2(A[8]), .A3(A[7]), .A4(A[6]), .ZN(n10) );
  NAND4_X1 U9 ( .A1(A[5]), .A2(A[4]), .A3(A[3]), .A4(A[31]), .ZN(n9) );
  NAND4_X1 U10 ( .A1(A[30]), .A2(A[2]), .A3(A[29]), .A4(A[28]), .ZN(n8) );
  NAND4_X1 U11 ( .A1(A[27]), .A2(A[26]), .A3(A[25]), .A4(A[24]), .ZN(n7) );
endmodule


module FFT_0 ( T, CLK, EN, RST, Q );
  input T, CLK, EN, RST;
  output Q;
  wire   n2, n3, n5;

  DFF_X1 TMP_reg ( .D(n5), .CK(CLK), .Q(Q) );
  XOR2_X1 U4 ( .A(n3), .B(Q), .Z(n2) );
  NAND2_X1 U5 ( .A1(T), .A2(EN), .ZN(n3) );
  NOR2_X1 U3 ( .A1(RST), .A2(n2), .ZN(n5) );
endmodule


module N_AND_N23 ( A, Y );
  input [22:0] A;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;

  NAND4_X1 U1 ( .A1(A[9]), .A2(A[8]), .A3(n5), .A4(A[7]), .ZN(n4) );
  NAND4_X1 U2 ( .A1(A[3]), .A2(A[2]), .A3(A[4]), .A4(n6), .ZN(n3) );
  NOR4_X1 U3 ( .A1(n1), .A2(n2), .A3(n3), .A4(n4), .ZN(Y) );
  NAND4_X1 U4 ( .A1(A[13]), .A2(A[12]), .A3(A[14]), .A4(n8), .ZN(n1) );
  NAND4_X1 U5 ( .A1(A[19]), .A2(A[18]), .A3(A[1]), .A4(n7), .ZN(n2) );
  AND3_X1 U6 ( .A1(A[16]), .A2(A[15]), .A3(A[17]), .ZN(n7) );
  AND3_X1 U7 ( .A1(A[10]), .A2(A[0]), .A3(A[11]), .ZN(n8) );
  AND3_X1 U8 ( .A1(A[21]), .A2(A[20]), .A3(A[22]), .ZN(n6) );
  AND2_X1 U9 ( .A1(A[6]), .A2(A[5]), .ZN(n5) );
endmodule


module N_AND_N5_0 ( A, Y );
  input [4:0] A;
  output Y;
  wire   n1;

  AND3_X1 U1 ( .A1(A[4]), .A2(A[3]), .A3(n1), .ZN(Y) );
  AND3_X1 U2 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .ZN(n1) );
endmodule


module XNOR_GATE_0 ( A, B, Y );
  input A, B;
  output Y;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(Y) );
endmodule


module MUX61_GEN_N32 ( A, B, C, D, E, F, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [31:0] F;
  input [2:0] SEL;
  output [31:0] Y;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n1, n2, n3, n4, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98;

  NAND2_X1 U75 ( .A1(n5), .A2(n6), .ZN(Y[9]) );
  NAND2_X1 U76 ( .A1(n13), .A2(n14), .ZN(Y[8]) );
  NAND2_X1 U77 ( .A1(n15), .A2(n16), .ZN(Y[7]) );
  NAND2_X1 U78 ( .A1(n17), .A2(n18), .ZN(Y[6]) );
  NAND2_X1 U79 ( .A1(n19), .A2(n20), .ZN(Y[5]) );
  NAND2_X1 U80 ( .A1(n21), .A2(n22), .ZN(Y[4]) );
  NAND2_X1 U81 ( .A1(n23), .A2(n24), .ZN(Y[3]) );
  NAND2_X1 U82 ( .A1(n25), .A2(n26), .ZN(Y[31]) );
  NAND2_X1 U83 ( .A1(n27), .A2(n28), .ZN(Y[30]) );
  NAND2_X1 U84 ( .A1(n29), .A2(n30), .ZN(Y[2]) );
  NAND2_X1 U85 ( .A1(n31), .A2(n32), .ZN(Y[29]) );
  NAND2_X1 U86 ( .A1(n33), .A2(n34), .ZN(Y[28]) );
  NAND2_X1 U87 ( .A1(n35), .A2(n36), .ZN(Y[27]) );
  NAND2_X1 U88 ( .A1(n37), .A2(n38), .ZN(Y[26]) );
  NAND2_X1 U89 ( .A1(n39), .A2(n40), .ZN(Y[25]) );
  NAND2_X1 U90 ( .A1(n41), .A2(n42), .ZN(Y[24]) );
  NAND2_X1 U91 ( .A1(n43), .A2(n44), .ZN(Y[23]) );
  NAND2_X1 U92 ( .A1(n45), .A2(n46), .ZN(Y[22]) );
  NAND2_X1 U93 ( .A1(n47), .A2(n48), .ZN(Y[21]) );
  NAND2_X1 U94 ( .A1(n49), .A2(n50), .ZN(Y[20]) );
  NAND2_X1 U95 ( .A1(n51), .A2(n52), .ZN(Y[1]) );
  NAND2_X1 U96 ( .A1(n53), .A2(n54), .ZN(Y[19]) );
  NAND2_X1 U97 ( .A1(n55), .A2(n56), .ZN(Y[18]) );
  NAND2_X1 U98 ( .A1(n57), .A2(n58), .ZN(Y[17]) );
  NAND2_X1 U99 ( .A1(n59), .A2(n60), .ZN(Y[16]) );
  NAND2_X1 U100 ( .A1(n61), .A2(n62), .ZN(Y[15]) );
  NAND2_X1 U101 ( .A1(n63), .A2(n64), .ZN(Y[14]) );
  NAND2_X1 U102 ( .A1(n65), .A2(n66), .ZN(Y[13]) );
  NAND2_X1 U103 ( .A1(n67), .A2(n68), .ZN(Y[12]) );
  NAND2_X1 U104 ( .A1(n69), .A2(n70), .ZN(Y[11]) );
  NAND2_X1 U105 ( .A1(n71), .A2(n72), .ZN(Y[10]) );
  NAND2_X1 U106 ( .A1(n73), .A2(n74), .ZN(Y[0]) );
  BUF_X1 U1 ( .A(n7), .Z(n96) );
  AOI222_X1 U2 ( .A1(E[0]), .A2(n98), .B1(B[0]), .B2(n93), .C1(D[0]), .C2(n92), 
        .ZN(n74) );
  AND3_X1 U3 ( .A1(n4), .A2(n79), .A3(n80), .ZN(n28) );
  AND3_X1 U4 ( .A1(n1), .A2(n2), .A3(n3), .ZN(n26) );
  NAND2_X1 U5 ( .A1(E[31]), .A2(n96), .ZN(n1) );
  NAND2_X1 U6 ( .A1(B[31]), .A2(n94), .ZN(n2) );
  NAND2_X1 U7 ( .A1(D[31]), .A2(n90), .ZN(n3) );
  NAND2_X1 U8 ( .A1(E[30]), .A2(n96), .ZN(n4) );
  NAND2_X1 U9 ( .A1(B[30]), .A2(n94), .ZN(n79) );
  NAND2_X1 U10 ( .A1(D[30]), .A2(n90), .ZN(n80) );
  BUF_X1 U11 ( .A(n11), .Z(n84) );
  BUF_X1 U12 ( .A(n11), .Z(n85) );
  BUF_X1 U13 ( .A(n11), .Z(n86) );
  NOR4_X1 U14 ( .A1(n81), .A2(n87), .A3(n93), .A4(n75), .ZN(n11) );
  OR2_X1 U15 ( .A1(n98), .A2(n92), .ZN(n75) );
  BUF_X1 U16 ( .A(n12), .Z(n81) );
  BUF_X1 U17 ( .A(n12), .Z(n82) );
  BUF_X1 U18 ( .A(n10), .Z(n87) );
  BUF_X1 U19 ( .A(n10), .Z(n88) );
  BUF_X1 U20 ( .A(n12), .Z(n83) );
  BUF_X1 U21 ( .A(n10), .Z(n89) );
  NOR3_X1 U22 ( .A1(n76), .A2(SEL[1]), .A3(n78), .ZN(n12) );
  NOR3_X1 U23 ( .A1(n76), .A2(n77), .A3(n78), .ZN(n10) );
  BUF_X1 U24 ( .A(n8), .Z(n93) );
  BUF_X1 U25 ( .A(n8), .Z(n94) );
  BUF_X1 U26 ( .A(n9), .Z(n91) );
  BUF_X1 U27 ( .A(n9), .Z(n90) );
  BUF_X1 U28 ( .A(n7), .Z(n97) );
  BUF_X1 U29 ( .A(n8), .Z(n95) );
  BUF_X1 U30 ( .A(n9), .Z(n92) );
  BUF_X1 U31 ( .A(n7), .Z(n98) );
  INV_X1 U32 ( .A(SEL[1]), .ZN(n77) );
  NOR3_X1 U33 ( .A1(n77), .A2(SEL[0]), .A3(n76), .ZN(n8) );
  NOR3_X1 U34 ( .A1(n77), .A2(SEL[2]), .A3(n78), .ZN(n7) );
  NOR3_X1 U35 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n76), .ZN(n9) );
  INV_X1 U36 ( .A(SEL[2]), .ZN(n76) );
  INV_X1 U37 ( .A(SEL[0]), .ZN(n78) );
  AOI222_X1 U38 ( .A1(E[3]), .A2(n96), .B1(B[3]), .B2(n95), .C1(D[3]), .C2(n90), .ZN(n24) );
  AOI222_X1 U39 ( .A1(E[4]), .A2(n96), .B1(B[4]), .B2(n95), .C1(D[4]), .C2(n90), .ZN(n22) );
  AOI222_X1 U40 ( .A1(E[5]), .A2(n96), .B1(B[5]), .B2(n95), .C1(D[5]), .C2(n90), .ZN(n20) );
  AOI222_X1 U41 ( .A1(E[6]), .A2(n96), .B1(B[6]), .B2(n95), .C1(D[6]), .C2(n90), .ZN(n18) );
  AOI222_X1 U42 ( .A1(E[7]), .A2(n96), .B1(B[7]), .B2(n95), .C1(D[7]), .C2(n90), .ZN(n16) );
  AOI222_X1 U43 ( .A1(E[8]), .A2(n96), .B1(B[8]), .B2(n95), .C1(D[8]), .C2(n90), .ZN(n14) );
  AOI222_X1 U44 ( .A1(E[9]), .A2(n96), .B1(B[9]), .B2(n95), .C1(D[9]), .C2(n90), .ZN(n6) );
  AOI222_X1 U45 ( .A1(E[29]), .A2(n96), .B1(B[29]), .B2(n94), .C1(D[29]), .C2(
        n90), .ZN(n32) );
  AOI222_X1 U46 ( .A1(E[1]), .A2(n97), .B1(B[1]), .B2(n93), .C1(D[1]), .C2(n91), .ZN(n52) );
  AOI222_X1 U47 ( .A1(E[2]), .A2(n96), .B1(B[2]), .B2(n94), .C1(D[2]), .C2(n90), .ZN(n30) );
  AOI222_X1 U48 ( .A1(E[10]), .A2(n98), .B1(B[10]), .B2(n93), .C1(D[10]), .C2(
        n92), .ZN(n72) );
  AOI222_X1 U49 ( .A1(E[11]), .A2(n98), .B1(B[11]), .B2(n93), .C1(D[11]), .C2(
        n92), .ZN(n70) );
  AOI222_X1 U50 ( .A1(E[12]), .A2(n98), .B1(B[12]), .B2(n93), .C1(D[12]), .C2(
        n92), .ZN(n68) );
  AOI222_X1 U51 ( .A1(E[13]), .A2(n98), .B1(B[13]), .B2(n93), .C1(D[13]), .C2(
        n92), .ZN(n66) );
  AOI222_X1 U52 ( .A1(E[14]), .A2(n98), .B1(B[14]), .B2(n93), .C1(D[14]), .C2(
        n92), .ZN(n64) );
  AOI222_X1 U53 ( .A1(E[17]), .A2(n97), .B1(B[17]), .B2(n93), .C1(D[17]), .C2(
        n91), .ZN(n58) );
  AOI222_X1 U54 ( .A1(E[19]), .A2(n97), .B1(B[19]), .B2(n93), .C1(D[19]), .C2(
        n91), .ZN(n54) );
  AOI222_X1 U55 ( .A1(E[21]), .A2(n97), .B1(B[21]), .B2(n94), .C1(D[21]), .C2(
        n91), .ZN(n48) );
  AOI222_X1 U56 ( .A1(E[22]), .A2(n97), .B1(B[22]), .B2(n94), .C1(D[22]), .C2(
        n91), .ZN(n46) );
  AOI222_X1 U57 ( .A1(E[23]), .A2(n97), .B1(B[23]), .B2(n94), .C1(D[23]), .C2(
        n91), .ZN(n44) );
  AOI222_X1 U58 ( .A1(E[26]), .A2(n97), .B1(B[26]), .B2(n94), .C1(D[26]), .C2(
        n91), .ZN(n38) );
  AOI222_X1 U59 ( .A1(A[0]), .A2(n87), .B1(F[0]), .B2(n84), .C1(C[0]), .C2(n81), .ZN(n73) );
  AOI222_X1 U60 ( .A1(A[1]), .A2(n87), .B1(F[1]), .B2(n84), .C1(C[1]), .C2(n81), .ZN(n51) );
  AOI222_X1 U61 ( .A1(A[2]), .A2(n88), .B1(F[2]), .B2(n85), .C1(C[2]), .C2(n82), .ZN(n29) );
  AOI222_X1 U62 ( .A1(A[3]), .A2(n89), .B1(F[3]), .B2(n85), .C1(C[3]), .C2(n83), .ZN(n23) );
  AOI222_X1 U63 ( .A1(A[4]), .A2(n89), .B1(F[4]), .B2(n86), .C1(C[4]), .C2(n83), .ZN(n21) );
  AOI222_X1 U64 ( .A1(A[5]), .A2(n89), .B1(F[5]), .B2(n86), .C1(C[5]), .C2(n83), .ZN(n19) );
  AOI222_X1 U65 ( .A1(A[6]), .A2(n89), .B1(F[6]), .B2(n86), .C1(C[6]), .C2(n83), .ZN(n17) );
  AOI222_X1 U66 ( .A1(A[7]), .A2(n89), .B1(F[7]), .B2(n86), .C1(C[7]), .C2(n83), .ZN(n15) );
  AOI222_X1 U67 ( .A1(A[8]), .A2(n89), .B1(F[8]), .B2(n86), .C1(C[8]), .C2(n83), .ZN(n13) );
  AOI222_X1 U68 ( .A1(A[9]), .A2(n89), .B1(F[9]), .B2(n86), .C1(C[9]), .C2(n83), .ZN(n5) );
  AOI222_X1 U69 ( .A1(A[10]), .A2(n87), .B1(F[10]), .B2(n84), .C1(C[10]), .C2(
        n81), .ZN(n71) );
  AOI222_X1 U70 ( .A1(A[11]), .A2(n87), .B1(F[11]), .B2(n84), .C1(C[11]), .C2(
        n81), .ZN(n69) );
  AOI222_X1 U71 ( .A1(A[12]), .A2(n87), .B1(F[12]), .B2(n84), .C1(C[12]), .C2(
        n81), .ZN(n67) );
  AOI222_X1 U72 ( .A1(A[13]), .A2(n87), .B1(F[13]), .B2(n84), .C1(C[13]), .C2(
        n81), .ZN(n65) );
  AOI222_X1 U73 ( .A1(A[14]), .A2(n87), .B1(F[14]), .B2(n84), .C1(C[14]), .C2(
        n81), .ZN(n63) );
  AOI222_X1 U74 ( .A1(A[15]), .A2(n87), .B1(F[15]), .B2(n84), .C1(C[15]), .C2(
        n81), .ZN(n61) );
  AOI222_X1 U107 ( .A1(A[16]), .A2(n87), .B1(F[16]), .B2(n84), .C1(C[16]), 
        .C2(n81), .ZN(n59) );
  AOI222_X1 U108 ( .A1(A[17]), .A2(n87), .B1(F[17]), .B2(n84), .C1(C[17]), 
        .C2(n81), .ZN(n57) );
  AOI222_X1 U109 ( .A1(A[18]), .A2(n87), .B1(F[18]), .B2(n84), .C1(C[18]), 
        .C2(n81), .ZN(n55) );
  AOI222_X1 U110 ( .A1(A[19]), .A2(n87), .B1(F[19]), .B2(n84), .C1(C[19]), 
        .C2(n81), .ZN(n53) );
  AOI222_X1 U111 ( .A1(A[20]), .A2(n88), .B1(F[20]), .B2(n84), .C1(C[20]), 
        .C2(n82), .ZN(n49) );
  AOI222_X1 U112 ( .A1(A[21]), .A2(n88), .B1(F[21]), .B2(n85), .C1(C[21]), 
        .C2(n82), .ZN(n47) );
  AOI222_X1 U113 ( .A1(A[22]), .A2(n88), .B1(F[22]), .B2(n85), .C1(C[22]), 
        .C2(n82), .ZN(n45) );
  AOI222_X1 U114 ( .A1(A[23]), .A2(n88), .B1(F[23]), .B2(n85), .C1(C[23]), 
        .C2(n82), .ZN(n43) );
  AOI222_X1 U115 ( .A1(A[24]), .A2(n88), .B1(F[24]), .B2(n85), .C1(C[24]), 
        .C2(n82), .ZN(n41) );
  AOI222_X1 U116 ( .A1(A[25]), .A2(n88), .B1(F[25]), .B2(n85), .C1(C[25]), 
        .C2(n82), .ZN(n39) );
  AOI222_X1 U117 ( .A1(A[26]), .A2(n88), .B1(F[26]), .B2(n85), .C1(C[26]), 
        .C2(n82), .ZN(n37) );
  AOI222_X1 U118 ( .A1(A[27]), .A2(n88), .B1(F[27]), .B2(n85), .C1(C[27]), 
        .C2(n82), .ZN(n35) );
  AOI222_X1 U119 ( .A1(A[28]), .A2(n88), .B1(F[28]), .B2(n85), .C1(C[28]), 
        .C2(n82), .ZN(n33) );
  AOI222_X1 U120 ( .A1(A[29]), .A2(n88), .B1(F[29]), .B2(n85), .C1(C[29]), 
        .C2(n82), .ZN(n31) );
  AOI222_X1 U121 ( .A1(A[30]), .A2(n88), .B1(F[30]), .B2(n85), .C1(C[30]), 
        .C2(n82), .ZN(n27) );
  AOI222_X1 U122 ( .A1(A[31]), .A2(n88), .B1(F[31]), .B2(n85), .C1(C[31]), 
        .C2(n82), .ZN(n25) );
  AOI222_X1 U123 ( .A1(E[16]), .A2(n97), .B1(B[16]), .B2(n93), .C1(D[16]), 
        .C2(n91), .ZN(n60) );
  AOI222_X1 U124 ( .A1(E[27]), .A2(n96), .B1(B[27]), .B2(n94), .C1(D[27]), 
        .C2(n90), .ZN(n36) );
  AOI222_X1 U125 ( .A1(E[28]), .A2(n96), .B1(B[28]), .B2(n94), .C1(D[28]), 
        .C2(n90), .ZN(n34) );
  AOI222_X1 U126 ( .A1(E[15]), .A2(n97), .B1(B[15]), .B2(n93), .C1(D[15]), 
        .C2(n91), .ZN(n62) );
  AOI222_X1 U127 ( .A1(E[18]), .A2(n97), .B1(B[18]), .B2(n93), .C1(D[18]), 
        .C2(n91), .ZN(n56) );
  AOI222_X1 U128 ( .A1(E[20]), .A2(n97), .B1(B[20]), .B2(n94), .C1(D[20]), 
        .C2(n91), .ZN(n50) );
  AOI222_X1 U129 ( .A1(E[24]), .A2(n97), .B1(B[24]), .B2(n94), .C1(D[24]), 
        .C2(n91), .ZN(n42) );
  AOI222_X1 U130 ( .A1(E[25]), .A2(n97), .B1(B[25]), .B2(n94), .C1(D[25]), 
        .C2(n91), .ZN(n40) );
endmodule


module NR_DIVISOR ( CLK, RST, EN, Z, D, Q, R, ADD_IN_D, ADD_IN_R, SIGN, 
        ADD_OUT );
  input [15:0] Z;
  input [15:0] D;
  output [15:0] Q;
  output [15:0] R;
  output [15:0] ADD_IN_D;
  output [15:0] ADD_IN_R;
  input [15:0] ADD_OUT;
  input CLK, RST, EN;
  output SIGN;
  wire   MSB_REM, SEL_R_MUX_IN, SEL_Q_MUX_IN, SEL_D_MUX, EN_D, EN_Z, EN_Q,
         EN_R, EN_SIGN;
  wire   [1:0] SEL_ADD_IN_D_MUX;
  wire   [1:0] SEL_ADD_IN_R_MUX;
  wire   [1:0] SEL_SIGN_MUX;

  NR_DIVISOR_DATAPATH INST_DATAPATH ( .CLK(CLK), .RST(RST), .Z(Z), .D(D), .Q(Q), .R(R), .MSB_REM(MSB_REM), .ADD_IN_D(ADD_IN_D), .ADD_IN_R(ADD_IN_R), .SIGN(
        SIGN), .ADD_OUT(ADD_OUT), .SEL_R_MUX_IN(SEL_R_MUX_IN), .SEL_Q_MUX_IN(
        SEL_Q_MUX_IN), .SEL_D_MUX(SEL_D_MUX), .SEL_ADD_IN_D_MUX(
        SEL_ADD_IN_D_MUX), .SEL_ADD_IN_R_MUX(SEL_ADD_IN_R_MUX), .SEL_SIGN_MUX(
        SEL_SIGN_MUX), .EN_D(EN_D), .EN_Z(EN_Z), .EN_Q(EN_Q), .EN_R(EN_R), 
        .EN_SIGN(EN_SIGN) );
  FSM_DIVISOR INST_FSM ( .CLK(CLK), .RST(RST), .EN(EN), .SEL_R_MUX_IN(
        SEL_R_MUX_IN), .SEL_Q_MUX_IN(SEL_Q_MUX_IN), .SEL_D_MUX(SEL_D_MUX), 
        .SEL_ADD_IN_D_MUX(SEL_ADD_IN_D_MUX), .SEL_ADD_IN_R_MUX(
        SEL_ADD_IN_R_MUX), .SEL_SIGN_MUX(SEL_SIGN_MUX), .EN_D(EN_D), .EN_Z(
        EN_Z), .EN_Q(EN_Q), .EN_R(EN_R), .EN_SIGN(EN_SIGN), .MSB_REM(MSB_REM)
         );
endmodule


module BOOTHMUL ( A, B, CLK, EN, RST, P );
  input [15:0] A;
  input [15:0] B;
  output [31:0] P;
  input CLK, EN, RST;
  wire   P_31, n1, n2, n3, n4, n5, n6;
  wire   [15:0] NOT_A;
  wire   [15:0] NEG_A;
  wire   [20:0] OUT_1;
  wire   [3:0] P_1;
  wire   [16:0] IN_COMP_2;
  wire   [15:0] A_1;
  wire   [15:0] B_1;
  wire   [15:0] NEG_A_1;
  wire   [22:0] OUT_2;
  wire   [16:0] IN_COMP_3;
  wire   [15:0] A_2;
  wire   [15:0] B_2;
  wire   [15:0] NEG_A_2;
  assign P[31] = P_31;
  assign P[30] = P_31;

  RCA_GEN_NO_C_N16 NEG_A_GEN ( .A({n3, NOT_A[14:0]}), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b1}), .S(NEG_A) );
  BOOTHMUL_COMP_1 COMP_1 ( .A(A), .NEG_A(NEG_A), .B(B), .P(OUT_1) );
  REG_N4 PIPE_1_0 ( .D(OUT_1[3:0]), .Q(P_1), .EN(EN), .RST(n6), .CLK(CLK) );
  REG_N17_0 PIPE_1_1 ( .D(OUT_1[20:4]), .Q(IN_COMP_2), .EN(EN), .RST(n6), 
        .CLK(CLK) );
  REG_N16_0 PIPE_1_2 ( .D(A), .Q(A_1), .EN(EN), .RST(n4), .CLK(CLK) );
  REG_N16_5 PIPE_1_3 ( .D(B), .Q(B_1), .EN(EN), .RST(n5), .CLK(CLK) );
  REG_N16_4 PIPE_1_4 ( .D(NEG_A), .Q(NEG_A_1), .EN(EN), .RST(n6), .CLK(CLK) );
  BOOTHMUL_COMP_2 COMP_2 ( .PREVIOUS(IN_COMP_2), .A(A_1), .NEG_A(NEG_A_1), .B(
        B_1), .P(OUT_2) );
  REG_N10 PIPE_2_0 ( .D({OUT_2[5:0], P_1}), .Q(P[9:0]), .EN(EN), .RST(n6), 
        .CLK(CLK) );
  REG_N17_1 PIPE_2_1 ( .D(OUT_2[22:6]), .Q(IN_COMP_3), .EN(EN), .RST(n4), 
        .CLK(CLK) );
  REG_N16_3 PIPE_2_2 ( .D(A_1), .Q(A_2), .EN(EN), .RST(n5), .CLK(CLK) );
  REG_N16_2 PIPE_2_3 ( .D({B_1[15:8], n1, n2, B_1[5:0]}), .Q(B_2), .EN(EN), 
        .RST(n5), .CLK(CLK) );
  REG_N16_1 PIPE_2_4 ( .D(NEG_A_1), .Q(NEG_A_2), .EN(EN), .RST(n4), .CLK(CLK)
         );
  BOOTHMUL_COMP_3 COMP_3 ( .PREVIOUS(IN_COMP_3), .A(A_2), .NEG_A(NEG_A_2), .B(
        B_2), .P({P_31, P[29:10]}) );
  CLKBUF_X1 U3 ( .A(B_1[7]), .Z(n1) );
  INV_X4 U4 ( .A(A[1]), .ZN(NOT_A[1]) );
  INV_X4 U5 ( .A(A[0]), .ZN(NOT_A[0]) );
  INV_X2 U6 ( .A(A[2]), .ZN(NOT_A[2]) );
  INV_X2 U7 ( .A(A[3]), .ZN(NOT_A[3]) );
  INV_X1 U8 ( .A(A[4]), .ZN(NOT_A[4]) );
  CLKBUF_X1 U9 ( .A(B_1[6]), .Z(n2) );
  INV_X1 U10 ( .A(A[6]), .ZN(NOT_A[6]) );
  INV_X1 U11 ( .A(A[7]), .ZN(NOT_A[7]) );
  INV_X1 U12 ( .A(A[8]), .ZN(NOT_A[8]) );
  INV_X1 U13 ( .A(A[9]), .ZN(NOT_A[9]) );
  INV_X1 U14 ( .A(A[10]), .ZN(NOT_A[10]) );
  INV_X1 U15 ( .A(A[11]), .ZN(NOT_A[11]) );
  INV_X1 U16 ( .A(A[12]), .ZN(NOT_A[12]) );
  INV_X1 U17 ( .A(A[13]), .ZN(NOT_A[13]) );
  INV_X1 U18 ( .A(A[14]), .ZN(NOT_A[14]) );
  INV_X1 U19 ( .A(A[5]), .ZN(NOT_A[5]) );
  BUF_X1 U20 ( .A(RST), .Z(n6) );
  BUF_X1 U21 ( .A(RST), .Z(n5) );
  BUF_X1 U22 ( .A(RST), .Z(n4) );
  INV_X1 U23 ( .A(A[15]), .ZN(n3) );
endmodule


module T2_SHIFTER_N32 ( A, B, ARITH_LOG, RIGHT_LEFT, Y );
  input [31:0] A;
  input [4:0] B;
  output [31:0] Y;
  input ARITH_LOG, RIGHT_LEFT;
  wire   \SIGN[6] , n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [38:0] MASK_00;
  wire   [38:0] MASK_08;
  wire   [38:0] MASK_16;
  wire   [38:0] MASK_24;
  wire   [38:0] SEL_MASK;
  wire   [2:0] SEL;

  XOR2_X1 U2 ( .A(n7), .B(B[2]), .Z(SEL[2]) );
  XOR2_X1 U3 ( .A(n8), .B(B[1]), .Z(SEL[1]) );
  XOR2_X1 U4 ( .A(n9), .B(B[0]), .Z(SEL[0]) );
  MUX21_1 ARITH_MUX ( .A(A[31]), .B(1'b0), .S(ARITH_LOG), .Y(\SIGN[6] ) );
  MUX21_GEN_N8_0 MUXS_00_1_0 ( .A(A[7:0]), .B({A[0], 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .SEL(n7), .Y(MASK_00[7:0]) );
  MUX21_GEN_N8_15 MUXS_00_2_1 ( .A(A[15:8]), .B(A[8:1]), .SEL(n7), .Y(
        MASK_00[15:8]) );
  MUX21_GEN_N8_14 MUXS_00_2_2 ( .A(A[23:16]), .B(A[16:9]), .SEL(n7), .Y(
        MASK_00[23:16]) );
  MUX21_GEN_N8_13 MUXS_00_2_3 ( .A(A[31:24]), .B(A[24:17]), .SEL(n7), .Y(
        MASK_00[31:24]) );
  MUX21_GEN_N7_0 MUXS_00_3_4 ( .A({n6, n6, n6, n6, n6, n6, n6}), .B(A[31:25]), 
        .SEL(n9), .Y(MASK_00[38:32]) );
  MUX21_GEN_N8_12 MUXS_08_1_0 ( .A(A[15:8]), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .SEL(n7), .Y(MASK_08[7:0]) );
  MUX21_GEN_N8_11 MUXS_08_2_1_1 ( .A(A[23:16]), .B({A[0], 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .SEL(n7), .Y(MASK_08[15:8]) );
  MUX21_GEN_N8_10 MUXS_08_2_2_2 ( .A(A[31:24]), .B(A[8:1]), .SEL(n8), .Y(
        MASK_08[23:16]) );
  MUX21_GEN_N8_9 MUXS_08_2_3_3 ( .A({n3, n3, n3, n2, n2, n2, n2, n2}), .B(
        A[16:9]), .SEL(n8), .Y(MASK_08[31:24]) );
  MUX21_GEN_N7_3 MUXS_08_3_4 ( .A({n1, n1, n1, n1, n1, n1, n1}), .B(A[31:25]), 
        .SEL(n9), .Y(MASK_08[38:32]) );
  MUX21_GEN_N8_8 MUXS_16_1_0 ( .A(A[23:16]), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .SEL(n7), .Y(MASK_16[7:0]) );
  MUX21_GEN_N8_7 MUXS_16_1_1 ( .A(A[31:24]), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .SEL(n8), .Y(MASK_16[15:8]) );
  MUX21_GEN_N8_6 MUXS_16_2_2 ( .A({n3, n3, n3, n3, n3, n3, n3, n3}), .B({A[0], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL(n8), .Y(
        MASK_16[23:16]) );
  MUX21_GEN_N8_5 MUXS_16_3_3 ( .A({n4, n4, n4, n4, n4, n4, n3, n3}), .B(A[8:1]), .SEL(n8), .Y(MASK_16[31:24]) );
  MUX21_GEN_N7_2 MUXS_16_3_4 ( .A({n2, n1, n1, n1, n1, n1, n1}), .B(A[15:9]), 
        .SEL(n9), .Y(MASK_16[38:32]) );
  MUX21_GEN_N8_4 MUXS_24_1_0 ( .A(A[31:24]), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .SEL(n8), .Y(MASK_24[7:0]) );
  MUX21_GEN_N8_3 MUXS_24_2_1 ( .A({n5, n4, n4, n4, n4, n4, n4, n4}), .B({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL(n8), .Y(MASK_24[15:8]) );
  MUX21_GEN_N8_2 MUXS_24_2_2 ( .A({n5, n5, n5, n5, n5, n5, n5, n5}), .B({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL(n8), .Y(
        MASK_24[23:16]) );
  MUX21_GEN_N8_1 MUXS_24_3_3 ( .A({n6, n6, n6, n6, n5, n5, n5, n5}), .B({A[0], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL(n7), .Y(
        MASK_24[31:24]) );
  MUX21_GEN_N7_1 MUXS_24_4_4 ( .A({n2, n2, n2, n2, n2, n2, n2}), .B(A[7:1]), 
        .SEL(n9), .Y(MASK_24[38:32]) );
  MUX41_GEN_N39 COARSE_GRAIN ( .A(MASK_24), .B(MASK_16), .C(MASK_08), .D(
        MASK_00), .SEL(B[4:3]), .Y(SEL_MASK) );
  MUX81_GEN_N32 FINE_GRAIN ( .A(SEL_MASK[31:0]), .B(SEL_MASK[32:1]), .C(
        SEL_MASK[33:2]), .D(SEL_MASK[34:3]), .E(SEL_MASK[35:4]), .F(
        SEL_MASK[36:5]), .G(SEL_MASK[37:6]), .H(SEL_MASK[38:7]), .SEL(SEL), 
        .Y(Y) );
  BUF_X1 U5 ( .A(RIGHT_LEFT), .Z(n9) );
  BUF_X2 U6 ( .A(RIGHT_LEFT), .Z(n8) );
  BUF_X2 U7 ( .A(RIGHT_LEFT), .Z(n7) );
  BUF_X1 U8 ( .A(\SIGN[6] ), .Z(n5) );
  BUF_X1 U9 ( .A(\SIGN[6] ), .Z(n4) );
  BUF_X1 U10 ( .A(\SIGN[6] ), .Z(n3) );
  BUF_X1 U11 ( .A(\SIGN[6] ), .Z(n2) );
  BUF_X1 U12 ( .A(\SIGN[6] ), .Z(n1) );
  BUF_X1 U13 ( .A(\SIGN[6] ), .Z(n6) );
endmodule


module T2_LOGICALS_N32 ( OP, A, B, Y );
  input [3:0] OP;
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  wire   \NAND_IN_1[31][1] , \NAND_IN_1[31][0] , \NAND_IN_1[30][1] ,
         \NAND_IN_1[30][0] , \NAND_IN_1[29][1] , \NAND_IN_1[29][0] ,
         \NAND_IN_1[28][1] , \NAND_IN_1[28][0] , \NAND_IN_1[27][1] ,
         \NAND_IN_1[27][0] , \NAND_IN_1[26][1] , \NAND_IN_1[26][0] ,
         \NAND_IN_1[25][1] , \NAND_IN_1[25][0] , \NAND_IN_1[24][1] ,
         \NAND_IN_1[24][0] , \NAND_IN_1[23][1] , \NAND_IN_1[23][0] ,
         \NAND_IN_1[22][1] , \NAND_IN_1[22][0] , \NAND_IN_1[21][1] ,
         \NAND_IN_1[21][0] , \NAND_IN_1[20][1] , \NAND_IN_1[20][0] ,
         \NAND_IN_1[19][1] , \NAND_IN_1[19][0] , \NAND_IN_1[18][1] ,
         \NAND_IN_1[18][0] , \NAND_IN_1[17][1] , \NAND_IN_1[17][0] ,
         \NAND_IN_1[16][1] , \NAND_IN_1[16][0] , \NAND_IN_1[15][1] ,
         \NAND_IN_1[15][0] , \NAND_IN_1[14][1] , \NAND_IN_1[14][0] ,
         \NAND_IN_1[13][1] , \NAND_IN_1[13][0] , \NAND_IN_1[12][1] ,
         \NAND_IN_1[12][0] , \NAND_IN_1[11][1] , \NAND_IN_1[11][0] ,
         \NAND_IN_1[10][1] , \NAND_IN_1[10][0] , \NAND_IN_1[9][1] ,
         \NAND_IN_1[9][0] , \NAND_IN_1[8][1] , \NAND_IN_1[8][0] ,
         \NAND_IN_1[7][1] , \NAND_IN_1[7][0] , \NAND_IN_1[6][1] ,
         \NAND_IN_1[6][0] , \NAND_IN_1[5][1] , \NAND_IN_1[5][0] ,
         \NAND_IN_1[4][1] , \NAND_IN_1[4][0] , \NAND_IN_1[3][1] ,
         \NAND_IN_1[3][0] , \NAND_IN_1[2][1] , \NAND_IN_1[2][0] ,
         \NAND_IN_1[1][1] , \NAND_IN_1[1][0] , \NAND_IN_1[0][1] ,
         \NAND_IN_1[0][0] , \NAND_IN_5[31][3] , \NAND_IN_5[31][2] ,
         \NAND_IN_5[31][1] , \NAND_IN_5[31][0] , \NAND_IN_5[30][3] ,
         \NAND_IN_5[30][2] , \NAND_IN_5[30][1] , \NAND_IN_5[30][0] ,
         \NAND_IN_5[29][3] , \NAND_IN_5[29][2] , \NAND_IN_5[29][1] ,
         \NAND_IN_5[29][0] , \NAND_IN_5[28][3] , \NAND_IN_5[28][2] ,
         \NAND_IN_5[28][1] , \NAND_IN_5[28][0] , \NAND_IN_5[27][3] ,
         \NAND_IN_5[27][2] , \NAND_IN_5[27][1] , \NAND_IN_5[27][0] ,
         \NAND_IN_5[26][3] , \NAND_IN_5[26][2] , \NAND_IN_5[26][1] ,
         \NAND_IN_5[26][0] , \NAND_IN_5[25][3] , \NAND_IN_5[25][2] ,
         \NAND_IN_5[25][1] , \NAND_IN_5[25][0] , \NAND_IN_5[24][3] ,
         \NAND_IN_5[24][2] , \NAND_IN_5[24][1] , \NAND_IN_5[24][0] ,
         \NAND_IN_5[23][3] , \NAND_IN_5[23][2] , \NAND_IN_5[23][1] ,
         \NAND_IN_5[23][0] , \NAND_IN_5[22][3] , \NAND_IN_5[22][2] ,
         \NAND_IN_5[22][1] , \NAND_IN_5[22][0] , \NAND_IN_5[21][3] ,
         \NAND_IN_5[21][2] , \NAND_IN_5[21][1] , \NAND_IN_5[21][0] ,
         \NAND_IN_5[20][3] , \NAND_IN_5[20][2] , \NAND_IN_5[20][1] ,
         \NAND_IN_5[20][0] , \NAND_IN_5[19][3] , \NAND_IN_5[19][2] ,
         \NAND_IN_5[19][1] , \NAND_IN_5[19][0] , \NAND_IN_5[18][3] ,
         \NAND_IN_5[18][2] , \NAND_IN_5[18][1] , \NAND_IN_5[18][0] ,
         \NAND_IN_5[17][3] , \NAND_IN_5[17][2] , \NAND_IN_5[17][1] ,
         \NAND_IN_5[17][0] , \NAND_IN_5[16][3] , \NAND_IN_5[16][2] ,
         \NAND_IN_5[16][1] , \NAND_IN_5[16][0] , \NAND_IN_5[15][3] ,
         \NAND_IN_5[15][2] , \NAND_IN_5[15][1] , \NAND_IN_5[15][0] ,
         \NAND_IN_5[14][3] , \NAND_IN_5[14][2] , \NAND_IN_5[14][1] ,
         \NAND_IN_5[14][0] , \NAND_IN_5[13][3] , \NAND_IN_5[13][2] ,
         \NAND_IN_5[13][1] , \NAND_IN_5[13][0] , \NAND_IN_5[12][3] ,
         \NAND_IN_5[12][2] , \NAND_IN_5[12][1] , \NAND_IN_5[12][0] ,
         \NAND_IN_5[11][3] , \NAND_IN_5[11][2] , \NAND_IN_5[11][1] ,
         \NAND_IN_5[11][0] , \NAND_IN_5[10][3] , \NAND_IN_5[10][2] ,
         \NAND_IN_5[10][1] , \NAND_IN_5[10][0] , \NAND_IN_5[9][3] ,
         \NAND_IN_5[9][2] , \NAND_IN_5[9][1] , \NAND_IN_5[9][0] ,
         \NAND_IN_5[8][3] , \NAND_IN_5[8][2] , \NAND_IN_5[8][1] ,
         \NAND_IN_5[8][0] , \NAND_IN_5[7][3] , \NAND_IN_5[7][2] ,
         \NAND_IN_5[7][1] , \NAND_IN_5[7][0] , \NAND_IN_5[6][3] ,
         \NAND_IN_5[6][2] , \NAND_IN_5[6][1] , \NAND_IN_5[6][0] ,
         \NAND_IN_5[5][3] , \NAND_IN_5[5][2] , \NAND_IN_5[5][1] ,
         \NAND_IN_5[5][0] , \NAND_IN_5[4][3] , \NAND_IN_5[4][2] ,
         \NAND_IN_5[4][1] , \NAND_IN_5[4][0] , \NAND_IN_5[3][3] ,
         \NAND_IN_5[3][2] , \NAND_IN_5[3][1] , \NAND_IN_5[3][0] ,
         \NAND_IN_5[2][3] , \NAND_IN_5[2][2] , \NAND_IN_5[2][1] ,
         \NAND_IN_5[2][0] , \NAND_IN_5[1][3] , \NAND_IN_5[1][2] ,
         \NAND_IN_5[1][1] , \NAND_IN_5[1][0] , \NAND_IN_5[0][3] ,
         \NAND_IN_5[0][2] , \NAND_IN_5[0][1] , \NAND_IN_5[0][0] , n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12;

  INV_1_103 INVERTING_1_0 ( .A(A[0]), .Y(\NAND_IN_1[0][1] ) );
  INV_1_102 INVERTING_1_1 ( .A(A[1]), .Y(\NAND_IN_1[1][1] ) );
  INV_1_101 INVERTING_1_2 ( .A(A[2]), .Y(\NAND_IN_1[2][1] ) );
  INV_1_100 INVERTING_1_3 ( .A(A[3]), .Y(\NAND_IN_1[3][1] ) );
  INV_1_99 INVERTING_1_4 ( .A(A[4]), .Y(\NAND_IN_1[4][1] ) );
  INV_1_98 INVERTING_1_5 ( .A(A[5]), .Y(\NAND_IN_1[5][1] ) );
  INV_1_97 INVERTING_1_6 ( .A(A[6]), .Y(\NAND_IN_1[6][1] ) );
  INV_1_96 INVERTING_1_7 ( .A(A[7]), .Y(\NAND_IN_1[7][1] ) );
  INV_1_95 INVERTING_1_8 ( .A(A[8]), .Y(\NAND_IN_1[8][1] ) );
  INV_1_94 INVERTING_1_9 ( .A(A[9]), .Y(\NAND_IN_1[9][1] ) );
  INV_1_93 INVERTING_1_10 ( .A(A[10]), .Y(\NAND_IN_1[10][1] ) );
  INV_1_92 INVERTING_1_11 ( .A(A[11]), .Y(\NAND_IN_1[11][1] ) );
  INV_1_91 INVERTING_1_12 ( .A(A[12]), .Y(\NAND_IN_1[12][1] ) );
  INV_1_90 INVERTING_1_13 ( .A(A[13]), .Y(\NAND_IN_1[13][1] ) );
  INV_1_89 INVERTING_1_14 ( .A(A[14]), .Y(\NAND_IN_1[14][1] ) );
  INV_1_88 INVERTING_1_15 ( .A(A[15]), .Y(\NAND_IN_1[15][1] ) );
  INV_1_87 INVERTING_1_16 ( .A(A[16]), .Y(\NAND_IN_1[16][1] ) );
  INV_1_86 INVERTING_1_17 ( .A(A[17]), .Y(\NAND_IN_1[17][1] ) );
  INV_1_85 INVERTING_1_18 ( .A(A[18]), .Y(\NAND_IN_1[18][1] ) );
  INV_1_84 INVERTING_1_19 ( .A(A[19]), .Y(\NAND_IN_1[19][1] ) );
  INV_1_83 INVERTING_1_20 ( .A(A[20]), .Y(\NAND_IN_1[20][1] ) );
  INV_1_82 INVERTING_1_21 ( .A(A[21]), .Y(\NAND_IN_1[21][1] ) );
  INV_1_81 INVERTING_1_22 ( .A(A[22]), .Y(\NAND_IN_1[22][1] ) );
  INV_1_80 INVERTING_1_23 ( .A(A[23]), .Y(\NAND_IN_1[23][1] ) );
  INV_1_79 INVERTING_1_24 ( .A(A[24]), .Y(\NAND_IN_1[24][1] ) );
  INV_1_78 INVERTING_1_25 ( .A(A[25]), .Y(\NAND_IN_1[25][1] ) );
  INV_1_77 INVERTING_1_26 ( .A(A[26]), .Y(\NAND_IN_1[26][1] ) );
  INV_1_76 INVERTING_1_27 ( .A(A[27]), .Y(\NAND_IN_1[27][1] ) );
  INV_1_75 INVERTING_1_28 ( .A(A[28]), .Y(\NAND_IN_1[28][1] ) );
  INV_1_74 INVERTING_1_29 ( .A(A[29]), .Y(\NAND_IN_1[29][1] ) );
  INV_1_73 INVERTING_1_30 ( .A(A[30]), .Y(\NAND_IN_1[30][1] ) );
  INV_1_72 INVERTING_1_31 ( .A(A[31]), .Y(\NAND_IN_1[31][1] ) );
  INV_1_71 INVERTING_2_0 ( .A(B[0]), .Y(\NAND_IN_1[0][0] ) );
  INV_1_70 INVERTING_2_1 ( .A(B[1]), .Y(\NAND_IN_1[1][0] ) );
  INV_1_69 INVERTING_2_2 ( .A(B[2]), .Y(\NAND_IN_1[2][0] ) );
  INV_1_68 INVERTING_2_3 ( .A(B[3]), .Y(\NAND_IN_1[3][0] ) );
  INV_1_67 INVERTING_2_4 ( .A(B[4]), .Y(\NAND_IN_1[4][0] ) );
  INV_1_66 INVERTING_2_5 ( .A(B[5]), .Y(\NAND_IN_1[5][0] ) );
  INV_1_65 INVERTING_2_6 ( .A(B[6]), .Y(\NAND_IN_1[6][0] ) );
  INV_1_64 INVERTING_2_7 ( .A(B[7]), .Y(\NAND_IN_1[7][0] ) );
  INV_1_63 INVERTING_2_8 ( .A(B[8]), .Y(\NAND_IN_1[8][0] ) );
  INV_1_62 INVERTING_2_9 ( .A(B[9]), .Y(\NAND_IN_1[9][0] ) );
  INV_1_61 INVERTING_2_10 ( .A(B[10]), .Y(\NAND_IN_1[10][0] ) );
  INV_1_60 INVERTING_2_11 ( .A(B[11]), .Y(\NAND_IN_1[11][0] ) );
  INV_1_59 INVERTING_2_12 ( .A(B[12]), .Y(\NAND_IN_1[12][0] ) );
  INV_1_58 INVERTING_2_13 ( .A(B[13]), .Y(\NAND_IN_1[13][0] ) );
  INV_1_57 INVERTING_2_14 ( .A(B[14]), .Y(\NAND_IN_1[14][0] ) );
  INV_1_56 INVERTING_2_15 ( .A(B[15]), .Y(\NAND_IN_1[15][0] ) );
  INV_1_55 INVERTING_2_16 ( .A(B[16]), .Y(\NAND_IN_1[16][0] ) );
  INV_1_54 INVERTING_2_17 ( .A(B[17]), .Y(\NAND_IN_1[17][0] ) );
  INV_1_53 INVERTING_2_18 ( .A(B[18]), .Y(\NAND_IN_1[18][0] ) );
  INV_1_52 INVERTING_2_19 ( .A(B[19]), .Y(\NAND_IN_1[19][0] ) );
  INV_1_51 INVERTING_2_20 ( .A(B[20]), .Y(\NAND_IN_1[20][0] ) );
  INV_1_50 INVERTING_2_21 ( .A(B[21]), .Y(\NAND_IN_1[21][0] ) );
  INV_1_49 INVERTING_2_22 ( .A(B[22]), .Y(\NAND_IN_1[22][0] ) );
  INV_1_48 INVERTING_2_23 ( .A(B[23]), .Y(\NAND_IN_1[23][0] ) );
  INV_1_47 INVERTING_2_24 ( .A(B[24]), .Y(\NAND_IN_1[24][0] ) );
  INV_1_46 INVERTING_2_25 ( .A(B[25]), .Y(\NAND_IN_1[25][0] ) );
  INV_1_45 INVERTING_2_26 ( .A(B[26]), .Y(\NAND_IN_1[26][0] ) );
  INV_1_44 INVERTING_2_27 ( .A(B[27]), .Y(\NAND_IN_1[27][0] ) );
  INV_1_43 INVERTING_2_28 ( .A(B[28]), .Y(\NAND_IN_1[28][0] ) );
  INV_1_42 INVERTING_2_29 ( .A(B[29]), .Y(\NAND_IN_1[29][0] ) );
  INV_1_41 INVERTING_2_30 ( .A(B[30]), .Y(\NAND_IN_1[30][0] ) );
  INV_1_40 INVERTING_2_31 ( .A(B[31]), .Y(\NAND_IN_1[31][0] ) );
  N_NAND_N3_0 NANDS_1_0 ( .A({n10, \NAND_IN_1[0][1] , \NAND_IN_1[0][0] }), .Y(
        \NAND_IN_5[0][0] ) );
  N_NAND_N3_127 NANDS_1_1 ( .A({n12, \NAND_IN_1[1][1] , \NAND_IN_1[1][0] }), 
        .Y(\NAND_IN_5[1][0] ) );
  N_NAND_N3_126 NANDS_1_2 ( .A({n12, \NAND_IN_1[2][1] , \NAND_IN_1[2][0] }), 
        .Y(\NAND_IN_5[2][0] ) );
  N_NAND_N3_125 NANDS_1_3 ( .A({n12, \NAND_IN_1[3][1] , \NAND_IN_1[3][0] }), 
        .Y(\NAND_IN_5[3][0] ) );
  N_NAND_N3_124 NANDS_1_4 ( .A({n12, \NAND_IN_1[4][1] , \NAND_IN_1[4][0] }), 
        .Y(\NAND_IN_5[4][0] ) );
  N_NAND_N3_123 NANDS_1_5 ( .A({n12, \NAND_IN_1[5][1] , \NAND_IN_1[5][0] }), 
        .Y(\NAND_IN_5[5][0] ) );
  N_NAND_N3_122 NANDS_1_6 ( .A({n12, \NAND_IN_1[6][1] , \NAND_IN_1[6][0] }), 
        .Y(\NAND_IN_5[6][0] ) );
  N_NAND_N3_121 NANDS_1_7 ( .A({n11, \NAND_IN_1[7][1] , \NAND_IN_1[7][0] }), 
        .Y(\NAND_IN_5[7][0] ) );
  N_NAND_N3_120 NANDS_1_8 ( .A({n11, \NAND_IN_1[8][1] , \NAND_IN_1[8][0] }), 
        .Y(\NAND_IN_5[8][0] ) );
  N_NAND_N3_119 NANDS_1_9 ( .A({n11, \NAND_IN_1[9][1] , \NAND_IN_1[9][0] }), 
        .Y(\NAND_IN_5[9][0] ) );
  N_NAND_N3_118 NANDS_1_10 ( .A({n11, \NAND_IN_1[10][1] , \NAND_IN_1[10][0] }), 
        .Y(\NAND_IN_5[10][0] ) );
  N_NAND_N3_117 NANDS_1_11 ( .A({n11, \NAND_IN_1[11][1] , \NAND_IN_1[11][0] }), 
        .Y(\NAND_IN_5[11][0] ) );
  N_NAND_N3_116 NANDS_1_12 ( .A({n11, \NAND_IN_1[12][1] , \NAND_IN_1[12][0] }), 
        .Y(\NAND_IN_5[12][0] ) );
  N_NAND_N3_115 NANDS_1_13 ( .A({n11, \NAND_IN_1[13][1] , \NAND_IN_1[13][0] }), 
        .Y(\NAND_IN_5[13][0] ) );
  N_NAND_N3_114 NANDS_1_14 ( .A({n11, \NAND_IN_1[14][1] , \NAND_IN_1[14][0] }), 
        .Y(\NAND_IN_5[14][0] ) );
  N_NAND_N3_113 NANDS_1_15 ( .A({n11, \NAND_IN_1[15][1] , \NAND_IN_1[15][0] }), 
        .Y(\NAND_IN_5[15][0] ) );
  N_NAND_N3_112 NANDS_1_16 ( .A({n11, \NAND_IN_1[16][1] , \NAND_IN_1[16][0] }), 
        .Y(\NAND_IN_5[16][0] ) );
  N_NAND_N3_111 NANDS_1_17 ( .A({n11, \NAND_IN_1[17][1] , \NAND_IN_1[17][0] }), 
        .Y(\NAND_IN_5[17][0] ) );
  N_NAND_N3_110 NANDS_1_18 ( .A({n11, \NAND_IN_1[18][1] , \NAND_IN_1[18][0] }), 
        .Y(\NAND_IN_5[18][0] ) );
  N_NAND_N3_109 NANDS_1_19 ( .A({n11, \NAND_IN_1[19][1] , \NAND_IN_1[19][0] }), 
        .Y(\NAND_IN_5[19][0] ) );
  N_NAND_N3_108 NANDS_1_20 ( .A({n10, \NAND_IN_1[20][1] , \NAND_IN_1[20][0] }), 
        .Y(\NAND_IN_5[20][0] ) );
  N_NAND_N3_107 NANDS_1_21 ( .A({n10, \NAND_IN_1[21][1] , \NAND_IN_1[21][0] }), 
        .Y(\NAND_IN_5[21][0] ) );
  N_NAND_N3_106 NANDS_1_22 ( .A({n10, \NAND_IN_1[22][1] , \NAND_IN_1[22][0] }), 
        .Y(\NAND_IN_5[22][0] ) );
  N_NAND_N3_105 NANDS_1_23 ( .A({n10, \NAND_IN_1[23][1] , \NAND_IN_1[23][0] }), 
        .Y(\NAND_IN_5[23][0] ) );
  N_NAND_N3_104 NANDS_1_24 ( .A({n10, \NAND_IN_1[24][1] , \NAND_IN_1[24][0] }), 
        .Y(\NAND_IN_5[24][0] ) );
  N_NAND_N3_103 NANDS_1_25 ( .A({n10, \NAND_IN_1[25][1] , \NAND_IN_1[25][0] }), 
        .Y(\NAND_IN_5[25][0] ) );
  N_NAND_N3_102 NANDS_1_26 ( .A({n10, \NAND_IN_1[26][1] , \NAND_IN_1[26][0] }), 
        .Y(\NAND_IN_5[26][0] ) );
  N_NAND_N3_101 NANDS_1_27 ( .A({n10, \NAND_IN_1[27][1] , \NAND_IN_1[27][0] }), 
        .Y(\NAND_IN_5[27][0] ) );
  N_NAND_N3_100 NANDS_1_28 ( .A({n10, \NAND_IN_1[28][1] , \NAND_IN_1[28][0] }), 
        .Y(\NAND_IN_5[28][0] ) );
  N_NAND_N3_99 NANDS_1_29 ( .A({n10, \NAND_IN_1[29][1] , \NAND_IN_1[29][0] }), 
        .Y(\NAND_IN_5[29][0] ) );
  N_NAND_N3_98 NANDS_1_30 ( .A({n10, \NAND_IN_1[30][1] , \NAND_IN_1[30][0] }), 
        .Y(\NAND_IN_5[30][0] ) );
  N_NAND_N3_97 NANDS_1_31 ( .A({n10, \NAND_IN_1[31][1] , \NAND_IN_1[31][0] }), 
        .Y(\NAND_IN_5[31][0] ) );
  N_NAND_N3_96 NANDS_2_0 ( .A({n9, \NAND_IN_1[0][1] , B[0]}), .Y(
        \NAND_IN_5[0][1] ) );
  N_NAND_N3_95 NANDS_2_1 ( .A({n9, \NAND_IN_1[1][1] , B[1]}), .Y(
        \NAND_IN_5[1][1] ) );
  N_NAND_N3_94 NANDS_2_2 ( .A({n9, \NAND_IN_1[2][1] , B[2]}), .Y(
        \NAND_IN_5[2][1] ) );
  N_NAND_N3_93 NANDS_2_3 ( .A({n9, \NAND_IN_1[3][1] , B[3]}), .Y(
        \NAND_IN_5[3][1] ) );
  N_NAND_N3_92 NANDS_2_4 ( .A({n9, \NAND_IN_1[4][1] , B[4]}), .Y(
        \NAND_IN_5[4][1] ) );
  N_NAND_N3_91 NANDS_2_5 ( .A({n9, \NAND_IN_1[5][1] , B[5]}), .Y(
        \NAND_IN_5[5][1] ) );
  N_NAND_N3_90 NANDS_2_6 ( .A({n8, \NAND_IN_1[6][1] , B[6]}), .Y(
        \NAND_IN_5[6][1] ) );
  N_NAND_N3_89 NANDS_2_7 ( .A({n8, \NAND_IN_1[7][1] , B[7]}), .Y(
        \NAND_IN_5[7][1] ) );
  N_NAND_N3_88 NANDS_2_8 ( .A({n8, \NAND_IN_1[8][1] , B[8]}), .Y(
        \NAND_IN_5[8][1] ) );
  N_NAND_N3_87 NANDS_2_9 ( .A({n8, \NAND_IN_1[9][1] , B[9]}), .Y(
        \NAND_IN_5[9][1] ) );
  N_NAND_N3_86 NANDS_2_10 ( .A({n8, \NAND_IN_1[10][1] , B[10]}), .Y(
        \NAND_IN_5[10][1] ) );
  N_NAND_N3_85 NANDS_2_11 ( .A({n8, \NAND_IN_1[11][1] , B[11]}), .Y(
        \NAND_IN_5[11][1] ) );
  N_NAND_N3_84 NANDS_2_12 ( .A({n8, \NAND_IN_1[12][1] , B[12]}), .Y(
        \NAND_IN_5[12][1] ) );
  N_NAND_N3_83 NANDS_2_13 ( .A({n8, \NAND_IN_1[13][1] , B[13]}), .Y(
        \NAND_IN_5[13][1] ) );
  N_NAND_N3_82 NANDS_2_14 ( .A({n8, \NAND_IN_1[14][1] , B[14]}), .Y(
        \NAND_IN_5[14][1] ) );
  N_NAND_N3_81 NANDS_2_15 ( .A({n8, \NAND_IN_1[15][1] , B[15]}), .Y(
        \NAND_IN_5[15][1] ) );
  N_NAND_N3_80 NANDS_2_16 ( .A({n8, \NAND_IN_1[16][1] , B[16]}), .Y(
        \NAND_IN_5[16][1] ) );
  N_NAND_N3_79 NANDS_2_17 ( .A({n8, \NAND_IN_1[17][1] , B[17]}), .Y(
        \NAND_IN_5[17][1] ) );
  N_NAND_N3_78 NANDS_2_18 ( .A({n8, \NAND_IN_1[18][1] , B[18]}), .Y(
        \NAND_IN_5[18][1] ) );
  N_NAND_N3_77 NANDS_2_19 ( .A({n7, \NAND_IN_1[19][1] , B[19]}), .Y(
        \NAND_IN_5[19][1] ) );
  N_NAND_N3_76 NANDS_2_20 ( .A({n7, \NAND_IN_1[20][1] , B[20]}), .Y(
        \NAND_IN_5[20][1] ) );
  N_NAND_N3_75 NANDS_2_21 ( .A({n7, \NAND_IN_1[21][1] , B[21]}), .Y(
        \NAND_IN_5[21][1] ) );
  N_NAND_N3_74 NANDS_2_22 ( .A({n7, \NAND_IN_1[22][1] , B[22]}), .Y(
        \NAND_IN_5[22][1] ) );
  N_NAND_N3_73 NANDS_2_23 ( .A({n7, \NAND_IN_1[23][1] , B[23]}), .Y(
        \NAND_IN_5[23][1] ) );
  N_NAND_N3_72 NANDS_2_24 ( .A({n7, \NAND_IN_1[24][1] , B[24]}), .Y(
        \NAND_IN_5[24][1] ) );
  N_NAND_N3_71 NANDS_2_25 ( .A({n7, \NAND_IN_1[25][1] , B[25]}), .Y(
        \NAND_IN_5[25][1] ) );
  N_NAND_N3_70 NANDS_2_26 ( .A({n7, \NAND_IN_1[26][1] , B[26]}), .Y(
        \NAND_IN_5[26][1] ) );
  N_NAND_N3_69 NANDS_2_27 ( .A({n7, \NAND_IN_1[27][1] , B[27]}), .Y(
        \NAND_IN_5[27][1] ) );
  N_NAND_N3_68 NANDS_2_28 ( .A({n7, \NAND_IN_1[28][1] , B[28]}), .Y(
        \NAND_IN_5[28][1] ) );
  N_NAND_N3_67 NANDS_2_29 ( .A({n7, \NAND_IN_1[29][1] , B[29]}), .Y(
        \NAND_IN_5[29][1] ) );
  N_NAND_N3_66 NANDS_2_30 ( .A({n7, \NAND_IN_1[30][1] , B[30]}), .Y(
        \NAND_IN_5[30][1] ) );
  N_NAND_N3_65 NANDS_2_31 ( .A({n7, \NAND_IN_1[31][1] , B[31]}), .Y(
        \NAND_IN_5[31][1] ) );
  N_NAND_N3_64 NANDS_3_0 ( .A({n6, A[0], \NAND_IN_1[0][0] }), .Y(
        \NAND_IN_5[0][2] ) );
  N_NAND_N3_63 NANDS_3_1 ( .A({n6, A[1], \NAND_IN_1[1][0] }), .Y(
        \NAND_IN_5[1][2] ) );
  N_NAND_N3_62 NANDS_3_2 ( .A({n6, A[2], \NAND_IN_1[2][0] }), .Y(
        \NAND_IN_5[2][2] ) );
  N_NAND_N3_61 NANDS_3_3 ( .A({n6, A[3], \NAND_IN_1[3][0] }), .Y(
        \NAND_IN_5[3][2] ) );
  N_NAND_N3_60 NANDS_3_4 ( .A({n6, A[4], \NAND_IN_1[4][0] }), .Y(
        \NAND_IN_5[4][2] ) );
  N_NAND_N3_59 NANDS_3_5 ( .A({n6, A[5], \NAND_IN_1[5][0] }), .Y(
        \NAND_IN_5[5][2] ) );
  N_NAND_N3_58 NANDS_3_6 ( .A({n5, A[6], \NAND_IN_1[6][0] }), .Y(
        \NAND_IN_5[6][2] ) );
  N_NAND_N3_57 NANDS_3_7 ( .A({n5, A[7], \NAND_IN_1[7][0] }), .Y(
        \NAND_IN_5[7][2] ) );
  N_NAND_N3_56 NANDS_3_8 ( .A({n5, A[8], \NAND_IN_1[8][0] }), .Y(
        \NAND_IN_5[8][2] ) );
  N_NAND_N3_55 NANDS_3_9 ( .A({n5, A[9], \NAND_IN_1[9][0] }), .Y(
        \NAND_IN_5[9][2] ) );
  N_NAND_N3_54 NANDS_3_10 ( .A({n5, A[10], \NAND_IN_1[10][0] }), .Y(
        \NAND_IN_5[10][2] ) );
  N_NAND_N3_53 NANDS_3_11 ( .A({n5, A[11], \NAND_IN_1[11][0] }), .Y(
        \NAND_IN_5[11][2] ) );
  N_NAND_N3_52 NANDS_3_12 ( .A({n5, A[12], \NAND_IN_1[12][0] }), .Y(
        \NAND_IN_5[12][2] ) );
  N_NAND_N3_51 NANDS_3_13 ( .A({n5, A[13], \NAND_IN_1[13][0] }), .Y(
        \NAND_IN_5[13][2] ) );
  N_NAND_N3_50 NANDS_3_14 ( .A({n5, A[14], \NAND_IN_1[14][0] }), .Y(
        \NAND_IN_5[14][2] ) );
  N_NAND_N3_49 NANDS_3_15 ( .A({n5, A[15], \NAND_IN_1[15][0] }), .Y(
        \NAND_IN_5[15][2] ) );
  N_NAND_N3_48 NANDS_3_16 ( .A({n5, A[16], \NAND_IN_1[16][0] }), .Y(
        \NAND_IN_5[16][2] ) );
  N_NAND_N3_47 NANDS_3_17 ( .A({n5, A[17], \NAND_IN_1[17][0] }), .Y(
        \NAND_IN_5[17][2] ) );
  N_NAND_N3_46 NANDS_3_18 ( .A({n5, A[18], \NAND_IN_1[18][0] }), .Y(
        \NAND_IN_5[18][2] ) );
  N_NAND_N3_45 NANDS_3_19 ( .A({n4, A[19], \NAND_IN_1[19][0] }), .Y(
        \NAND_IN_5[19][2] ) );
  N_NAND_N3_44 NANDS_3_20 ( .A({n4, A[20], \NAND_IN_1[20][0] }), .Y(
        \NAND_IN_5[20][2] ) );
  N_NAND_N3_43 NANDS_3_21 ( .A({n4, A[21], \NAND_IN_1[21][0] }), .Y(
        \NAND_IN_5[21][2] ) );
  N_NAND_N3_42 NANDS_3_22 ( .A({n4, A[22], \NAND_IN_1[22][0] }), .Y(
        \NAND_IN_5[22][2] ) );
  N_NAND_N3_41 NANDS_3_23 ( .A({n4, A[23], \NAND_IN_1[23][0] }), .Y(
        \NAND_IN_5[23][2] ) );
  N_NAND_N3_40 NANDS_3_24 ( .A({n4, A[24], \NAND_IN_1[24][0] }), .Y(
        \NAND_IN_5[24][2] ) );
  N_NAND_N3_39 NANDS_3_25 ( .A({n4, A[25], \NAND_IN_1[25][0] }), .Y(
        \NAND_IN_5[25][2] ) );
  N_NAND_N3_38 NANDS_3_26 ( .A({n4, A[26], \NAND_IN_1[26][0] }), .Y(
        \NAND_IN_5[26][2] ) );
  N_NAND_N3_37 NANDS_3_27 ( .A({n4, A[27], \NAND_IN_1[27][0] }), .Y(
        \NAND_IN_5[27][2] ) );
  N_NAND_N3_36 NANDS_3_28 ( .A({n4, A[28], \NAND_IN_1[28][0] }), .Y(
        \NAND_IN_5[28][2] ) );
  N_NAND_N3_35 NANDS_3_29 ( .A({n4, A[29], \NAND_IN_1[29][0] }), .Y(
        \NAND_IN_5[29][2] ) );
  N_NAND_N3_34 NANDS_3_30 ( .A({n4, A[30], \NAND_IN_1[30][0] }), .Y(
        \NAND_IN_5[30][2] ) );
  N_NAND_N3_33 NANDS_3_31 ( .A({n4, A[31], \NAND_IN_1[31][0] }), .Y(
        \NAND_IN_5[31][2] ) );
  N_NAND_N3_32 NANDS_4_0 ( .A({n3, A[0], B[0]}), .Y(\NAND_IN_5[0][3] ) );
  N_NAND_N3_31 NANDS_4_1 ( .A({n3, A[1], B[1]}), .Y(\NAND_IN_5[1][3] ) );
  N_NAND_N3_30 NANDS_4_2 ( .A({n3, A[2], B[2]}), .Y(\NAND_IN_5[2][3] ) );
  N_NAND_N3_29 NANDS_4_3 ( .A({n3, A[3], B[3]}), .Y(\NAND_IN_5[3][3] ) );
  N_NAND_N3_28 NANDS_4_4 ( .A({n3, A[4], B[4]}), .Y(\NAND_IN_5[4][3] ) );
  N_NAND_N3_27 NANDS_4_5 ( .A({n3, A[5], B[5]}), .Y(\NAND_IN_5[5][3] ) );
  N_NAND_N3_26 NANDS_4_6 ( .A({n2, A[6], B[6]}), .Y(\NAND_IN_5[6][3] ) );
  N_NAND_N3_25 NANDS_4_7 ( .A({n2, A[7], B[7]}), .Y(\NAND_IN_5[7][3] ) );
  N_NAND_N3_24 NANDS_4_8 ( .A({n2, A[8], B[8]}), .Y(\NAND_IN_5[8][3] ) );
  N_NAND_N3_23 NANDS_4_9 ( .A({n2, A[9], B[9]}), .Y(\NAND_IN_5[9][3] ) );
  N_NAND_N3_22 NANDS_4_10 ( .A({n2, A[10], B[10]}), .Y(\NAND_IN_5[10][3] ) );
  N_NAND_N3_21 NANDS_4_11 ( .A({n2, A[11], B[11]}), .Y(\NAND_IN_5[11][3] ) );
  N_NAND_N3_20 NANDS_4_12 ( .A({n2, A[12], B[12]}), .Y(\NAND_IN_5[12][3] ) );
  N_NAND_N3_19 NANDS_4_13 ( .A({n2, A[13], B[13]}), .Y(\NAND_IN_5[13][3] ) );
  N_NAND_N3_18 NANDS_4_14 ( .A({n2, A[14], B[14]}), .Y(\NAND_IN_5[14][3] ) );
  N_NAND_N3_17 NANDS_4_15 ( .A({n2, A[15], B[15]}), .Y(\NAND_IN_5[15][3] ) );
  N_NAND_N3_16 NANDS_4_16 ( .A({n2, A[16], B[16]}), .Y(\NAND_IN_5[16][3] ) );
  N_NAND_N3_15 NANDS_4_17 ( .A({n2, A[17], B[17]}), .Y(\NAND_IN_5[17][3] ) );
  N_NAND_N3_14 NANDS_4_18 ( .A({n2, A[18], B[18]}), .Y(\NAND_IN_5[18][3] ) );
  N_NAND_N3_13 NANDS_4_19 ( .A({n1, A[19], B[19]}), .Y(\NAND_IN_5[19][3] ) );
  N_NAND_N3_12 NANDS_4_20 ( .A({n1, A[20], B[20]}), .Y(\NAND_IN_5[20][3] ) );
  N_NAND_N3_11 NANDS_4_21 ( .A({n1, A[21], B[21]}), .Y(\NAND_IN_5[21][3] ) );
  N_NAND_N3_10 NANDS_4_22 ( .A({n1, A[22], B[22]}), .Y(\NAND_IN_5[22][3] ) );
  N_NAND_N3_9 NANDS_4_23 ( .A({n1, A[23], B[23]}), .Y(\NAND_IN_5[23][3] ) );
  N_NAND_N3_8 NANDS_4_24 ( .A({n1, A[24], B[24]}), .Y(\NAND_IN_5[24][3] ) );
  N_NAND_N3_7 NANDS_4_25 ( .A({n1, A[25], B[25]}), .Y(\NAND_IN_5[25][3] ) );
  N_NAND_N3_6 NANDS_4_26 ( .A({n1, A[26], B[26]}), .Y(\NAND_IN_5[26][3] ) );
  N_NAND_N3_5 NANDS_4_27 ( .A({n1, A[27], B[27]}), .Y(\NAND_IN_5[27][3] ) );
  N_NAND_N3_4 NANDS_4_28 ( .A({n1, A[28], B[28]}), .Y(\NAND_IN_5[28][3] ) );
  N_NAND_N3_3 NANDS_4_29 ( .A({n1, A[29], B[29]}), .Y(\NAND_IN_5[29][3] ) );
  N_NAND_N3_2 NANDS_4_30 ( .A({n1, A[30], B[30]}), .Y(\NAND_IN_5[30][3] ) );
  N_NAND_N3_1 NANDS_4_31 ( .A({n1, A[31], B[31]}), .Y(\NAND_IN_5[31][3] ) );
  N_NAND_N4_0 NANDS_5_0 ( .A({\NAND_IN_5[0][3] , \NAND_IN_5[0][2] , 
        \NAND_IN_5[0][1] , \NAND_IN_5[0][0] }), .Y(Y[0]) );
  N_NAND_N4_31 NANDS_5_1 ( .A({\NAND_IN_5[1][3] , \NAND_IN_5[1][2] , 
        \NAND_IN_5[1][1] , \NAND_IN_5[1][0] }), .Y(Y[1]) );
  N_NAND_N4_30 NANDS_5_2 ( .A({\NAND_IN_5[2][3] , \NAND_IN_5[2][2] , 
        \NAND_IN_5[2][1] , \NAND_IN_5[2][0] }), .Y(Y[2]) );
  N_NAND_N4_29 NANDS_5_3 ( .A({\NAND_IN_5[3][3] , \NAND_IN_5[3][2] , 
        \NAND_IN_5[3][1] , \NAND_IN_5[3][0] }), .Y(Y[3]) );
  N_NAND_N4_28 NANDS_5_4 ( .A({\NAND_IN_5[4][3] , \NAND_IN_5[4][2] , 
        \NAND_IN_5[4][1] , \NAND_IN_5[4][0] }), .Y(Y[4]) );
  N_NAND_N4_27 NANDS_5_5 ( .A({\NAND_IN_5[5][3] , \NAND_IN_5[5][2] , 
        \NAND_IN_5[5][1] , \NAND_IN_5[5][0] }), .Y(Y[5]) );
  N_NAND_N4_26 NANDS_5_6 ( .A({\NAND_IN_5[6][3] , \NAND_IN_5[6][2] , 
        \NAND_IN_5[6][1] , \NAND_IN_5[6][0] }), .Y(Y[6]) );
  N_NAND_N4_25 NANDS_5_7 ( .A({\NAND_IN_5[7][3] , \NAND_IN_5[7][2] , 
        \NAND_IN_5[7][1] , \NAND_IN_5[7][0] }), .Y(Y[7]) );
  N_NAND_N4_24 NANDS_5_8 ( .A({\NAND_IN_5[8][3] , \NAND_IN_5[8][2] , 
        \NAND_IN_5[8][1] , \NAND_IN_5[8][0] }), .Y(Y[8]) );
  N_NAND_N4_23 NANDS_5_9 ( .A({\NAND_IN_5[9][3] , \NAND_IN_5[9][2] , 
        \NAND_IN_5[9][1] , \NAND_IN_5[9][0] }), .Y(Y[9]) );
  N_NAND_N4_22 NANDS_5_10 ( .A({\NAND_IN_5[10][3] , \NAND_IN_5[10][2] , 
        \NAND_IN_5[10][1] , \NAND_IN_5[10][0] }), .Y(Y[10]) );
  N_NAND_N4_21 NANDS_5_11 ( .A({\NAND_IN_5[11][3] , \NAND_IN_5[11][2] , 
        \NAND_IN_5[11][1] , \NAND_IN_5[11][0] }), .Y(Y[11]) );
  N_NAND_N4_20 NANDS_5_12 ( .A({\NAND_IN_5[12][3] , \NAND_IN_5[12][2] , 
        \NAND_IN_5[12][1] , \NAND_IN_5[12][0] }), .Y(Y[12]) );
  N_NAND_N4_19 NANDS_5_13 ( .A({\NAND_IN_5[13][3] , \NAND_IN_5[13][2] , 
        \NAND_IN_5[13][1] , \NAND_IN_5[13][0] }), .Y(Y[13]) );
  N_NAND_N4_18 NANDS_5_14 ( .A({\NAND_IN_5[14][3] , \NAND_IN_5[14][2] , 
        \NAND_IN_5[14][1] , \NAND_IN_5[14][0] }), .Y(Y[14]) );
  N_NAND_N4_17 NANDS_5_15 ( .A({\NAND_IN_5[15][3] , \NAND_IN_5[15][2] , 
        \NAND_IN_5[15][1] , \NAND_IN_5[15][0] }), .Y(Y[15]) );
  N_NAND_N4_16 NANDS_5_16 ( .A({\NAND_IN_5[16][3] , \NAND_IN_5[16][2] , 
        \NAND_IN_5[16][1] , \NAND_IN_5[16][0] }), .Y(Y[16]) );
  N_NAND_N4_15 NANDS_5_17 ( .A({\NAND_IN_5[17][3] , \NAND_IN_5[17][2] , 
        \NAND_IN_5[17][1] , \NAND_IN_5[17][0] }), .Y(Y[17]) );
  N_NAND_N4_14 NANDS_5_18 ( .A({\NAND_IN_5[18][3] , \NAND_IN_5[18][2] , 
        \NAND_IN_5[18][1] , \NAND_IN_5[18][0] }), .Y(Y[18]) );
  N_NAND_N4_13 NANDS_5_19 ( .A({\NAND_IN_5[19][3] , \NAND_IN_5[19][2] , 
        \NAND_IN_5[19][1] , \NAND_IN_5[19][0] }), .Y(Y[19]) );
  N_NAND_N4_12 NANDS_5_20 ( .A({\NAND_IN_5[20][3] , \NAND_IN_5[20][2] , 
        \NAND_IN_5[20][1] , \NAND_IN_5[20][0] }), .Y(Y[20]) );
  N_NAND_N4_11 NANDS_5_21 ( .A({\NAND_IN_5[21][3] , \NAND_IN_5[21][2] , 
        \NAND_IN_5[21][1] , \NAND_IN_5[21][0] }), .Y(Y[21]) );
  N_NAND_N4_10 NANDS_5_22 ( .A({\NAND_IN_5[22][3] , \NAND_IN_5[22][2] , 
        \NAND_IN_5[22][1] , \NAND_IN_5[22][0] }), .Y(Y[22]) );
  N_NAND_N4_9 NANDS_5_23 ( .A({\NAND_IN_5[23][3] , \NAND_IN_5[23][2] , 
        \NAND_IN_5[23][1] , \NAND_IN_5[23][0] }), .Y(Y[23]) );
  N_NAND_N4_8 NANDS_5_24 ( .A({\NAND_IN_5[24][3] , \NAND_IN_5[24][2] , 
        \NAND_IN_5[24][1] , \NAND_IN_5[24][0] }), .Y(Y[24]) );
  N_NAND_N4_7 NANDS_5_25 ( .A({\NAND_IN_5[25][3] , \NAND_IN_5[25][2] , 
        \NAND_IN_5[25][1] , \NAND_IN_5[25][0] }), .Y(Y[25]) );
  N_NAND_N4_6 NANDS_5_26 ( .A({\NAND_IN_5[26][3] , \NAND_IN_5[26][2] , 
        \NAND_IN_5[26][1] , \NAND_IN_5[26][0] }), .Y(Y[26]) );
  N_NAND_N4_5 NANDS_5_27 ( .A({\NAND_IN_5[27][3] , \NAND_IN_5[27][2] , 
        \NAND_IN_5[27][1] , \NAND_IN_5[27][0] }), .Y(Y[27]) );
  N_NAND_N4_4 NANDS_5_28 ( .A({\NAND_IN_5[28][3] , \NAND_IN_5[28][2] , 
        \NAND_IN_5[28][1] , \NAND_IN_5[28][0] }), .Y(Y[28]) );
  N_NAND_N4_3 NANDS_5_29 ( .A({\NAND_IN_5[29][3] , \NAND_IN_5[29][2] , 
        \NAND_IN_5[29][1] , \NAND_IN_5[29][0] }), .Y(Y[29]) );
  N_NAND_N4_2 NANDS_5_30 ( .A({\NAND_IN_5[30][3] , \NAND_IN_5[30][2] , 
        \NAND_IN_5[30][1] , \NAND_IN_5[30][0] }), .Y(Y[30]) );
  N_NAND_N4_1 NANDS_5_31 ( .A({\NAND_IN_5[31][3] , \NAND_IN_5[31][2] , 
        \NAND_IN_5[31][1] , \NAND_IN_5[31][0] }), .Y(Y[31]) );
  BUF_X1 U1 ( .A(OP[2]), .Z(n8) );
  BUF_X1 U2 ( .A(OP[1]), .Z(n5) );
  BUF_X1 U3 ( .A(OP[0]), .Z(n2) );
  BUF_X1 U4 ( .A(OP[3]), .Z(n11) );
  BUF_X1 U5 ( .A(OP[3]), .Z(n10) );
  BUF_X1 U6 ( .A(OP[2]), .Z(n7) );
  BUF_X1 U7 ( .A(OP[1]), .Z(n4) );
  BUF_X1 U8 ( .A(OP[0]), .Z(n1) );
  BUF_X1 U9 ( .A(OP[2]), .Z(n9) );
  BUF_X1 U10 ( .A(OP[1]), .Z(n6) );
  BUF_X1 U11 ( .A(OP[0]), .Z(n3) );
  BUF_X1 U12 ( .A(OP[3]), .Z(n12) );
endmodule


module CMP_N32 ( C, S, OP_SEL, UNSIGN, MSB_A, MSB_B, Y );
  input [31:0] S;
  input [2:0] OP_SEL;
  output [31:0] Y;
  input C, UNSIGN, MSB_A, MSB_B;
  wire   DIF, SIGN, MUX_SEL, NC, Z, NZ, G_UNSIGNED, G_SIGNED, OUT_MUX_G,
         GE_SIGNED, OUT_MUX_GE, LE_UNSIGNED, LE_SIGNED, OUT_MUX_LE, L_SIGNED,
         OUT_MUX_L;
  assign Y[31] = 1'b0;
  assign Y[30] = 1'b0;
  assign Y[29] = 1'b0;
  assign Y[28] = 1'b0;
  assign Y[27] = 1'b0;
  assign Y[26] = 1'b0;
  assign Y[25] = 1'b0;
  assign Y[24] = 1'b0;
  assign Y[23] = 1'b0;
  assign Y[22] = 1'b0;
  assign Y[21] = 1'b0;
  assign Y[20] = 1'b0;
  assign Y[19] = 1'b0;
  assign Y[18] = 1'b0;
  assign Y[17] = 1'b0;
  assign Y[16] = 1'b0;
  assign Y[15] = 1'b0;
  assign Y[14] = 1'b0;
  assign Y[13] = 1'b0;
  assign Y[12] = 1'b0;
  assign Y[11] = 1'b0;
  assign Y[10] = 1'b0;
  assign Y[9] = 1'b0;
  assign Y[8] = 1'b0;
  assign Y[7] = 1'b0;
  assign Y[6] = 1'b0;
  assign Y[5] = 1'b0;
  assign Y[4] = 1'b0;
  assign Y[3] = 1'b0;
  assign Y[2] = 1'b0;
  assign Y[1] = 1'b0;

  XOR_GATE_1 CHECK_SIGN ( .A(MSB_A), .B(MSB_B), .Y(DIF) );
  INV_1_110 INV_UNSIGN ( .A(UNSIGN), .Y(SIGN) );
  AND_GATE_1_644 GEN_SEL ( .A(DIF), .B(SIGN), .Y(MUX_SEL) );
  INV_1_109 INV_C ( .A(C), .Y(NC) );
  N_NOR_N32 N_NOR_INST ( .A(S), .Y(Z) );
  INV_1_108 INV_Z ( .A(Z), .Y(NZ) );
  AND_GATE_1_643 AND_INST ( .A(C), .B(NZ), .Y(G_UNSIGNED) );
  INV_1_107 INV_G ( .A(G_UNSIGNED), .Y(G_SIGNED) );
  MUX21_5 G_MUX ( .A(G_SIGNED), .B(G_UNSIGNED), .S(MUX_SEL), .Y(OUT_MUX_G) );
  INV_1_106 INV_GE ( .A(C), .Y(GE_SIGNED) );
  MUX21_4 GE_MUX ( .A(GE_SIGNED), .B(C), .S(MUX_SEL), .Y(OUT_MUX_GE) );
  OR_GATE_307 OR_INST ( .A(NC), .B(Z), .Y(LE_UNSIGNED) );
  INV_1_105 INV_LE ( .A(LE_UNSIGNED), .Y(LE_SIGNED) );
  MUX21_3 LE_MUX ( .A(LE_SIGNED), .B(LE_UNSIGNED), .S(MUX_SEL), .Y(OUT_MUX_LE)
         );
  INV_1_104 INV_L ( .A(NC), .Y(L_SIGNED) );
  MUX21_2 L_MUX ( .A(L_SIGNED), .B(NC), .S(MUX_SEL), .Y(OUT_MUX_L) );
  MUX61 MUX_INST ( .A(OUT_MUX_L), .B(OUT_MUX_LE), .C(Z), .D(NZ), .E(OUT_MUX_GE), .F(OUT_MUX_G), .SEL(OP_SEL), .Y(Y[0]) );
endmodule


module P4_ADDER_N32 ( A, B, Ci, Co, S );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;

  wire   [7:1] CARRY_VECTOR;

  CARRY_GENERATOR_N32 CARRY_GENERATION ( .A(A), .B(B), .Ci(Ci), .Co({Co, 
        CARRY_VECTOR}) );
  SUM_GENERATOR_N32 SUM_GENERATION ( .A(A), .B(B), .Ci({CARRY_VECTOR, Ci}), 
        .S(S) );
endmodule


module XOR_GATE_1_0 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module D_LATCH_0 ( D, EN, Q );
  input D, EN;
  output Q;
  wire   NOT_D, OUT_AND_1, OUT_AND_2, OUT_NOR_2;

  INV_169 INV_D ( .A(D), .Y(NOT_D) );
  AND_GATE_338 AND_1 ( .A(NOT_D), .B(EN), .Y(OUT_AND_1) );
  AND_GATE_337 AND_2 ( .A(D), .B(EN), .Y(OUT_AND_2) );
  NOR_GATE_0 NOR_1 ( .A(OUT_AND_1), .B(OUT_NOR_2), .Y(Q) );
  NOR_GATE_337 NOR_2 ( .A(OUT_AND_2), .B(Q), .Y(OUT_NOR_2) );
endmodule


module OR_GATE_0 ( A, B, Y );
  input A, B;
  output Y;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module MUX21_0 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  INV_1_111 UIV ( .A(S), .Y(SB) );
  NAND_GATE_921 UND1 ( .A(A), .B(S), .Y(Y1) );
  NAND_GATE_920 UND2 ( .A(B), .B(SB), .Y(Y2) );
  NAND_GATE_919 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GEN_N4_0 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   SB;
  wire   [3:0] Y1;
  wire   [3:0] Y2;

  INV_1_119 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_1017 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_1016 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_1015 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_1014 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_1013 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_1012 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_1011 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_1010 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_1009 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_1008 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_1007 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_1006 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
endmodule


module RCA_GEN_N4_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_269 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_268 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_267 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_266 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX41_0 ( A, B, C, D, SEL, Y );
  input [1:0] SEL;
  input A, B, C, D;
  output Y;
  wire   n5, n6, n7, n8, n9, n10, n11;

  NAND2_X1 U8 ( .A1(A), .A2(n5), .ZN(n7) );
  NOR2_X1 U1 ( .A1(n9), .A2(n11), .ZN(n5) );
  INV_X1 U2 ( .A(SEL[0]), .ZN(n11) );
  INV_X1 U3 ( .A(SEL[1]), .ZN(n9) );
  OAI21_X1 U4 ( .B1(n5), .B2(n6), .A(n7), .ZN(Y) );
  AOI22_X1 U5 ( .A1(n8), .A2(n9), .B1(B), .B2(SEL[1]), .ZN(n6) );
  INV_X1 U6 ( .A(n10), .ZN(n8) );
  AOI22_X1 U7 ( .A1(C), .A2(SEL[0]), .B1(D), .B2(n11), .ZN(n10) );
endmodule


module CACHE_DATA_BPU_N32_SET_BIT2 ( DATA_IN, DATA_OUT, ADDR, CLK, WE );
  input [31:0] DATA_IN;
  output [31:0] DATA_OUT;
  input [1:0] ADDR;
  input CLK, WE;
  wire   \CACHE_MEM[3][31] , \CACHE_MEM[3][30] , \CACHE_MEM[3][29] ,
         \CACHE_MEM[3][28] , \CACHE_MEM[3][27] , \CACHE_MEM[3][26] ,
         \CACHE_MEM[3][25] , \CACHE_MEM[3][24] , \CACHE_MEM[3][23] ,
         \CACHE_MEM[3][22] , \CACHE_MEM[3][21] , \CACHE_MEM[3][20] ,
         \CACHE_MEM[3][19] , \CACHE_MEM[3][18] , \CACHE_MEM[3][17] ,
         \CACHE_MEM[3][16] , \CACHE_MEM[3][15] , \CACHE_MEM[3][14] ,
         \CACHE_MEM[3][13] , \CACHE_MEM[3][12] , \CACHE_MEM[3][11] ,
         \CACHE_MEM[3][10] , \CACHE_MEM[3][9] , \CACHE_MEM[3][8] ,
         \CACHE_MEM[3][7] , \CACHE_MEM[3][6] , \CACHE_MEM[3][5] ,
         \CACHE_MEM[3][4] , \CACHE_MEM[3][3] , \CACHE_MEM[3][2] ,
         \CACHE_MEM[3][1] , \CACHE_MEM[3][0] , \CACHE_MEM[0][31] ,
         \CACHE_MEM[0][30] , \CACHE_MEM[0][29] , \CACHE_MEM[0][28] ,
         \CACHE_MEM[0][27] , \CACHE_MEM[0][26] , \CACHE_MEM[0][25] ,
         \CACHE_MEM[0][24] , \CACHE_MEM[0][23] , \CACHE_MEM[0][22] ,
         \CACHE_MEM[0][21] , \CACHE_MEM[0][20] , \CACHE_MEM[0][19] ,
         \CACHE_MEM[0][18] , \CACHE_MEM[0][17] , \CACHE_MEM[0][16] ,
         \CACHE_MEM[0][15] , \CACHE_MEM[0][14] , \CACHE_MEM[0][13] ,
         \CACHE_MEM[0][12] , \CACHE_MEM[0][11] , \CACHE_MEM[0][10] ,
         \CACHE_MEM[0][9] , \CACHE_MEM[0][8] , \CACHE_MEM[0][7] ,
         \CACHE_MEM[0][6] , \CACHE_MEM[0][5] , \CACHE_MEM[0][4] ,
         \CACHE_MEM[0][3] , \CACHE_MEM[0][2] , \CACHE_MEM[0][1] ,
         \CACHE_MEM[0][0] , n3, n4, n6, n8, n9, n10, n11, n12, n15, n18, n19,
         n21, n24, n25, n27, n30, n31, n33, n36, n37, n39, n42, n43, n45, n48,
         n49, n51, n54, n55, n57, n60, n61, n63, n66, n67, n69, n72, n73, n75,
         n78, n79, n81, n84, n85, n87, n90, n91, n93, n96, n97, n99, n102,
         n103, n105, n108, n109, n111, n114, n115, n117, n120, n121, n123,
         n126, n127, n129, n132, n133, n135, n138, n139, n141, n144, n145,
         n147, n150, n151, n153, n156, n157, n159, n162, n163, n165, n168,
         n169, n171, n174, n175, n177, n180, n181, n183, n186, n187, n189,
         n192, n193, n195, n198, n199, n202, n203, n205, n206, n369, n370,
         n372, n373, n374, n376, n377, n378, n380, n381, n382, n384, n385,
         n386, n388, n389, n390, n392, n393, n394, n396, n397, n398, n400,
         n401, n402, n404, n405, n406, n408, n409, n410, n412, n413, n414,
         n416, n417, n418, n420, n421, n422, n424, n425, n426, n428, n429,
         n430, n432, n433, n434, n436, n437, n438, n440, n441, n442, n444,
         n445, n446, n448, n449, n450, n452, n453, n454, n456, n457, n458,
         n460, n461, n462, n464, n465, n466, n468, n469, n470, n472, n473,
         n474, n476, n477, n478, n480, n481, n482, n484, n485, n486, n488,
         n489, n490, n492, n493, n494, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n1, n2, n5, n7, n13, n14, n16, n17, n20, n22, n23,
         n26, n28, n29, n32, n34, n35, n38, n40, n41, n44, n46, n47, n50, n52,
         n53, n56, n58, n59, n62, n64, n65, n68, n70, n71, n74, n76, n77, n80,
         n82, n83, n86, n88, n89, n92, n94, n95, n98, n100, n101, n104, n106,
         n107, n110, n112, n113, n116, n118, n119, n122, n124, n125, n128,
         n130, n131, n134, n136, n137, n140, n142, n143, n146, n148, n149,
         n152, n154, n155, n158, n160, n161, n164, n166, n167, n170, n172,
         n173, n176, n178, n179, n182, n184, n185, n188, n190, n191, n194,
         n196, n197, n200, n201, n204, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300;

  DFF_X1 \CACHE_MEM_reg[3][31]  ( .D(n592), .CK(CLK), .Q(\CACHE_MEM[3][31] ), 
        .QN(n196) );
  DFF_X1 \CACHE_MEM_reg[3][30]  ( .D(n591), .CK(CLK), .Q(\CACHE_MEM[3][30] ), 
        .QN(n194) );
  DFF_X1 \CACHE_MEM_reg[3][29]  ( .D(n590), .CK(CLK), .Q(\CACHE_MEM[3][29] ), 
        .QN(n191) );
  DFF_X1 \CACHE_MEM_reg[3][28]  ( .D(n589), .CK(CLK), .Q(\CACHE_MEM[3][28] ), 
        .QN(n190) );
  DFF_X1 \CACHE_MEM_reg[3][27]  ( .D(n588), .CK(CLK), .Q(\CACHE_MEM[3][27] ), 
        .QN(n188) );
  DFF_X1 \CACHE_MEM_reg[3][26]  ( .D(n587), .CK(CLK), .Q(\CACHE_MEM[3][26] ), 
        .QN(n185) );
  DFF_X1 \CACHE_MEM_reg[3][25]  ( .D(n586), .CK(CLK), .Q(\CACHE_MEM[3][25] ), 
        .QN(n184) );
  DFF_X1 \CACHE_MEM_reg[3][24]  ( .D(n585), .CK(CLK), .Q(\CACHE_MEM[3][24] ), 
        .QN(n182) );
  DFF_X1 \CACHE_MEM_reg[3][23]  ( .D(n584), .CK(CLK), .Q(\CACHE_MEM[3][23] ), 
        .QN(n179) );
  DFF_X1 \CACHE_MEM_reg[3][22]  ( .D(n583), .CK(CLK), .Q(\CACHE_MEM[3][22] ), 
        .QN(n178) );
  DFF_X1 \CACHE_MEM_reg[3][21]  ( .D(n582), .CK(CLK), .Q(\CACHE_MEM[3][21] ), 
        .QN(n176) );
  DFF_X1 \CACHE_MEM_reg[3][20]  ( .D(n581), .CK(CLK), .Q(\CACHE_MEM[3][20] ), 
        .QN(n173) );
  DFF_X1 \CACHE_MEM_reg[3][19]  ( .D(n580), .CK(CLK), .Q(\CACHE_MEM[3][19] ), 
        .QN(n172) );
  DFF_X1 \CACHE_MEM_reg[3][18]  ( .D(n579), .CK(CLK), .Q(\CACHE_MEM[3][18] ), 
        .QN(n170) );
  DFF_X1 \CACHE_MEM_reg[3][17]  ( .D(n578), .CK(CLK), .Q(\CACHE_MEM[3][17] ), 
        .QN(n167) );
  DFF_X1 \CACHE_MEM_reg[3][16]  ( .D(n577), .CK(CLK), .Q(\CACHE_MEM[3][16] ), 
        .QN(n166) );
  DFF_X1 \CACHE_MEM_reg[3][15]  ( .D(n576), .CK(CLK), .Q(\CACHE_MEM[3][15] ), 
        .QN(n164) );
  DFF_X1 \CACHE_MEM_reg[3][14]  ( .D(n575), .CK(CLK), .Q(\CACHE_MEM[3][14] ), 
        .QN(n161) );
  DFF_X1 \CACHE_MEM_reg[3][13]  ( .D(n574), .CK(CLK), .Q(\CACHE_MEM[3][13] ), 
        .QN(n160) );
  DFF_X1 \CACHE_MEM_reg[3][12]  ( .D(n573), .CK(CLK), .Q(\CACHE_MEM[3][12] ), 
        .QN(n158) );
  DFF_X1 \CACHE_MEM_reg[3][11]  ( .D(n572), .CK(CLK), .Q(\CACHE_MEM[3][11] ), 
        .QN(n155) );
  DFF_X1 \CACHE_MEM_reg[3][10]  ( .D(n571), .CK(CLK), .Q(\CACHE_MEM[3][10] ), 
        .QN(n154) );
  DFF_X1 \CACHE_MEM_reg[3][9]  ( .D(n570), .CK(CLK), .Q(\CACHE_MEM[3][9] ), 
        .QN(n152) );
  DFF_X1 \CACHE_MEM_reg[3][8]  ( .D(n569), .CK(CLK), .Q(\CACHE_MEM[3][8] ), 
        .QN(n149) );
  DFF_X1 \CACHE_MEM_reg[3][7]  ( .D(n568), .CK(CLK), .Q(\CACHE_MEM[3][7] ), 
        .QN(n148) );
  DFF_X1 \CACHE_MEM_reg[3][6]  ( .D(n567), .CK(CLK), .Q(\CACHE_MEM[3][6] ), 
        .QN(n146) );
  DFF_X1 \CACHE_MEM_reg[3][5]  ( .D(n566), .CK(CLK), .Q(\CACHE_MEM[3][5] ), 
        .QN(n143) );
  DFF_X1 \CACHE_MEM_reg[3][4]  ( .D(n565), .CK(CLK), .Q(\CACHE_MEM[3][4] ), 
        .QN(n142) );
  DFF_X1 \CACHE_MEM_reg[3][3]  ( .D(n564), .CK(CLK), .Q(\CACHE_MEM[3][3] ), 
        .QN(n140) );
  DFF_X1 \CACHE_MEM_reg[3][2]  ( .D(n563), .CK(CLK), .Q(\CACHE_MEM[3][2] ), 
        .QN(n137) );
  DFF_X1 \CACHE_MEM_reg[3][1]  ( .D(n562), .CK(CLK), .Q(\CACHE_MEM[3][1] ), 
        .QN(n136) );
  DFF_X1 \CACHE_MEM_reg[3][0]  ( .D(n561), .CK(CLK), .Q(\CACHE_MEM[3][0] ), 
        .QN(n134) );
  DFF_X1 \CACHE_MEM_reg[2][31]  ( .D(n560), .CK(CLK), .QN(n80) );
  DFF_X1 \CACHE_MEM_reg[2][30]  ( .D(n559), .CK(CLK), .QN(n77) );
  DFF_X1 \CACHE_MEM_reg[2][29]  ( .D(n558), .CK(CLK), .QN(n76) );
  DFF_X1 \CACHE_MEM_reg[2][28]  ( .D(n557), .CK(CLK), .QN(n74) );
  DFF_X1 \CACHE_MEM_reg[2][27]  ( .D(n556), .CK(CLK), .QN(n71) );
  DFF_X1 \CACHE_MEM_reg[2][26]  ( .D(n555), .CK(CLK), .QN(n70) );
  DFF_X1 \CACHE_MEM_reg[2][25]  ( .D(n554), .CK(CLK), .QN(n131) );
  DFF_X1 \CACHE_MEM_reg[2][24]  ( .D(n553), .CK(CLK), .QN(n130) );
  DFF_X1 \CACHE_MEM_reg[2][23]  ( .D(n552), .CK(CLK), .QN(n128) );
  DFF_X1 \CACHE_MEM_reg[2][22]  ( .D(n551), .CK(CLK), .QN(n125) );
  DFF_X1 \CACHE_MEM_reg[2][21]  ( .D(n550), .CK(CLK), .QN(n124) );
  DFF_X1 \CACHE_MEM_reg[2][20]  ( .D(n549), .CK(CLK), .QN(n122) );
  DFF_X1 \CACHE_MEM_reg[2][19]  ( .D(n548), .CK(CLK), .QN(n119) );
  DFF_X1 \CACHE_MEM_reg[2][18]  ( .D(n547), .CK(CLK), .QN(n118) );
  DFF_X1 \CACHE_MEM_reg[2][17]  ( .D(n546), .CK(CLK), .QN(n116) );
  DFF_X1 \CACHE_MEM_reg[2][16]  ( .D(n545), .CK(CLK), .QN(n113) );
  DFF_X1 \CACHE_MEM_reg[2][15]  ( .D(n544), .CK(CLK), .QN(n112) );
  DFF_X1 \CACHE_MEM_reg[2][14]  ( .D(n543), .CK(CLK), .QN(n110) );
  DFF_X1 \CACHE_MEM_reg[2][13]  ( .D(n542), .CK(CLK), .QN(n107) );
  DFF_X1 \CACHE_MEM_reg[2][12]  ( .D(n541), .CK(CLK), .QN(n106) );
  DFF_X1 \CACHE_MEM_reg[2][11]  ( .D(n540), .CK(CLK), .QN(n104) );
  DFF_X1 \CACHE_MEM_reg[2][10]  ( .D(n539), .CK(CLK), .QN(n101) );
  DFF_X1 \CACHE_MEM_reg[2][9]  ( .D(n538), .CK(CLK), .QN(n100) );
  DFF_X1 \CACHE_MEM_reg[2][8]  ( .D(n537), .CK(CLK), .QN(n98) );
  DFF_X1 \CACHE_MEM_reg[2][7]  ( .D(n536), .CK(CLK), .QN(n95) );
  DFF_X1 \CACHE_MEM_reg[2][6]  ( .D(n535), .CK(CLK), .QN(n94) );
  DFF_X1 \CACHE_MEM_reg[2][5]  ( .D(n534), .CK(CLK), .QN(n92) );
  DFF_X1 \CACHE_MEM_reg[2][4]  ( .D(n533), .CK(CLK), .QN(n89) );
  DFF_X1 \CACHE_MEM_reg[2][3]  ( .D(n532), .CK(CLK), .QN(n88) );
  DFF_X1 \CACHE_MEM_reg[2][2]  ( .D(n531), .CK(CLK), .QN(n86) );
  DFF_X1 \CACHE_MEM_reg[2][1]  ( .D(n530), .CK(CLK), .QN(n83) );
  DFF_X1 \CACHE_MEM_reg[2][0]  ( .D(n529), .CK(CLK), .QN(n82) );
  DFF_X1 \CACHE_MEM_reg[1][31]  ( .D(n528), .CK(CLK), .QN(n16) );
  DFF_X1 \CACHE_MEM_reg[1][30]  ( .D(n527), .CK(CLK), .QN(n14) );
  DFF_X1 \CACHE_MEM_reg[1][29]  ( .D(n526), .CK(CLK), .QN(n13) );
  DFF_X1 \CACHE_MEM_reg[1][28]  ( .D(n525), .CK(CLK), .QN(n7) );
  DFF_X1 \CACHE_MEM_reg[1][27]  ( .D(n524), .CK(CLK), .QN(n5) );
  DFF_X1 \CACHE_MEM_reg[1][26]  ( .D(n523), .CK(CLK), .QN(n2) );
  DFF_X1 \CACHE_MEM_reg[1][25]  ( .D(n522), .CK(CLK), .QN(n68) );
  DFF_X1 \CACHE_MEM_reg[1][24]  ( .D(n521), .CK(CLK), .QN(n65) );
  DFF_X1 \CACHE_MEM_reg[1][23]  ( .D(n520), .CK(CLK), .QN(n64) );
  DFF_X1 \CACHE_MEM_reg[1][22]  ( .D(n519), .CK(CLK), .QN(n62) );
  DFF_X1 \CACHE_MEM_reg[1][21]  ( .D(n518), .CK(CLK), .QN(n59) );
  DFF_X1 \CACHE_MEM_reg[1][20]  ( .D(n517), .CK(CLK), .QN(n58) );
  DFF_X1 \CACHE_MEM_reg[1][19]  ( .D(n516), .CK(CLK), .QN(n56) );
  DFF_X1 \CACHE_MEM_reg[1][18]  ( .D(n515), .CK(CLK), .QN(n53) );
  DFF_X1 \CACHE_MEM_reg[1][17]  ( .D(n514), .CK(CLK), .QN(n52) );
  DFF_X1 \CACHE_MEM_reg[1][16]  ( .D(n513), .CK(CLK), .QN(n50) );
  DFF_X1 \CACHE_MEM_reg[1][15]  ( .D(n512), .CK(CLK), .QN(n47) );
  DFF_X1 \CACHE_MEM_reg[1][14]  ( .D(n511), .CK(CLK), .QN(n46) );
  DFF_X1 \CACHE_MEM_reg[1][13]  ( .D(n510), .CK(CLK), .QN(n44) );
  DFF_X1 \CACHE_MEM_reg[1][12]  ( .D(n509), .CK(CLK), .QN(n41) );
  DFF_X1 \CACHE_MEM_reg[1][11]  ( .D(n508), .CK(CLK), .QN(n40) );
  DFF_X1 \CACHE_MEM_reg[1][10]  ( .D(n507), .CK(CLK), .QN(n38) );
  DFF_X1 \CACHE_MEM_reg[1][9]  ( .D(n506), .CK(CLK), .QN(n35) );
  DFF_X1 \CACHE_MEM_reg[1][8]  ( .D(n505), .CK(CLK), .QN(n34) );
  DFF_X1 \CACHE_MEM_reg[1][7]  ( .D(n504), .CK(CLK), .QN(n32) );
  DFF_X1 \CACHE_MEM_reg[1][6]  ( .D(n503), .CK(CLK), .QN(n29) );
  DFF_X1 \CACHE_MEM_reg[1][5]  ( .D(n502), .CK(CLK), .QN(n28) );
  DFF_X1 \CACHE_MEM_reg[1][4]  ( .D(n501), .CK(CLK), .QN(n26) );
  DFF_X1 \CACHE_MEM_reg[1][3]  ( .D(n500), .CK(CLK), .QN(n23) );
  DFF_X1 \CACHE_MEM_reg[1][2]  ( .D(n499), .CK(CLK), .QN(n22) );
  DFF_X1 \CACHE_MEM_reg[1][1]  ( .D(n498), .CK(CLK), .QN(n20) );
  DFF_X1 \CACHE_MEM_reg[1][0]  ( .D(n497), .CK(CLK), .QN(n17) );
  DFF_X1 \CACHE_MEM_reg[0][31]  ( .D(n496), .CK(CLK), .Q(\CACHE_MEM[0][31] ), 
        .QN(n208) );
  DFF_X1 \CACHE_MEM_reg[0][30]  ( .D(n492), .CK(CLK), .Q(\CACHE_MEM[0][30] ), 
        .QN(n207) );
  DFF_X1 \CACHE_MEM_reg[0][29]  ( .D(n488), .CK(CLK), .Q(\CACHE_MEM[0][29] ), 
        .QN(n204) );
  DFF_X1 \CACHE_MEM_reg[0][28]  ( .D(n484), .CK(CLK), .Q(\CACHE_MEM[0][28] ), 
        .QN(n201) );
  DFF_X1 \CACHE_MEM_reg[0][27]  ( .D(n480), .CK(CLK), .Q(\CACHE_MEM[0][27] ), 
        .QN(n200) );
  DFF_X1 \CACHE_MEM_reg[0][26]  ( .D(n476), .CK(CLK), .Q(\CACHE_MEM[0][26] ), 
        .QN(n197) );
  DFF_X1 \CACHE_MEM_reg[0][25]  ( .D(n472), .CK(CLK), .Q(\CACHE_MEM[0][25] ), 
        .QN(n234) );
  DFF_X1 \CACHE_MEM_reg[0][24]  ( .D(n468), .CK(CLK), .Q(\CACHE_MEM[0][24] ), 
        .QN(n233) );
  DFF_X1 \CACHE_MEM_reg[0][23]  ( .D(n464), .CK(CLK), .Q(\CACHE_MEM[0][23] ), 
        .QN(n232) );
  DFF_X1 \CACHE_MEM_reg[0][22]  ( .D(n460), .CK(CLK), .Q(\CACHE_MEM[0][22] ), 
        .QN(n231) );
  DFF_X1 \CACHE_MEM_reg[0][21]  ( .D(n456), .CK(CLK), .Q(\CACHE_MEM[0][21] ), 
        .QN(n230) );
  DFF_X1 \CACHE_MEM_reg[0][20]  ( .D(n452), .CK(CLK), .Q(\CACHE_MEM[0][20] ), 
        .QN(n229) );
  DFF_X1 \CACHE_MEM_reg[0][19]  ( .D(n448), .CK(CLK), .Q(\CACHE_MEM[0][19] ), 
        .QN(n228) );
  DFF_X1 \CACHE_MEM_reg[0][18]  ( .D(n444), .CK(CLK), .Q(\CACHE_MEM[0][18] ), 
        .QN(n227) );
  DFF_X1 \CACHE_MEM_reg[0][17]  ( .D(n440), .CK(CLK), .Q(\CACHE_MEM[0][17] ), 
        .QN(n226) );
  DFF_X1 \CACHE_MEM_reg[0][16]  ( .D(n436), .CK(CLK), .Q(\CACHE_MEM[0][16] ), 
        .QN(n225) );
  DFF_X1 \CACHE_MEM_reg[0][15]  ( .D(n432), .CK(CLK), .Q(\CACHE_MEM[0][15] ), 
        .QN(n224) );
  DFF_X1 \CACHE_MEM_reg[0][14]  ( .D(n428), .CK(CLK), .Q(\CACHE_MEM[0][14] ), 
        .QN(n223) );
  DFF_X1 \CACHE_MEM_reg[0][13]  ( .D(n424), .CK(CLK), .Q(\CACHE_MEM[0][13] ), 
        .QN(n222) );
  DFF_X1 \CACHE_MEM_reg[0][12]  ( .D(n420), .CK(CLK), .Q(\CACHE_MEM[0][12] ), 
        .QN(n221) );
  DFF_X1 \CACHE_MEM_reg[0][11]  ( .D(n416), .CK(CLK), .Q(\CACHE_MEM[0][11] ), 
        .QN(n220) );
  DFF_X1 \CACHE_MEM_reg[0][10]  ( .D(n412), .CK(CLK), .Q(\CACHE_MEM[0][10] ), 
        .QN(n219) );
  DFF_X1 \CACHE_MEM_reg[0][9]  ( .D(n408), .CK(CLK), .Q(\CACHE_MEM[0][9] ), 
        .QN(n218) );
  DFF_X1 \CACHE_MEM_reg[0][8]  ( .D(n404), .CK(CLK), .Q(\CACHE_MEM[0][8] ), 
        .QN(n217) );
  DFF_X1 \CACHE_MEM_reg[0][7]  ( .D(n400), .CK(CLK), .Q(\CACHE_MEM[0][7] ), 
        .QN(n216) );
  DFF_X1 \CACHE_MEM_reg[0][6]  ( .D(n396), .CK(CLK), .Q(\CACHE_MEM[0][6] ), 
        .QN(n215) );
  DFF_X1 \CACHE_MEM_reg[0][5]  ( .D(n392), .CK(CLK), .Q(\CACHE_MEM[0][5] ), 
        .QN(n214) );
  DFF_X1 \CACHE_MEM_reg[0][4]  ( .D(n388), .CK(CLK), .Q(\CACHE_MEM[0][4] ), 
        .QN(n213) );
  DFF_X1 \CACHE_MEM_reg[0][3]  ( .D(n384), .CK(CLK), .Q(\CACHE_MEM[0][3] ), 
        .QN(n212) );
  DFF_X1 \CACHE_MEM_reg[0][2]  ( .D(n380), .CK(CLK), .Q(\CACHE_MEM[0][2] ), 
        .QN(n211) );
  DFF_X1 \CACHE_MEM_reg[0][1]  ( .D(n376), .CK(CLK), .Q(\CACHE_MEM[0][1] ), 
        .QN(n210) );
  DFF_X1 \CACHE_MEM_reg[0][0]  ( .D(n372), .CK(CLK), .Q(\CACHE_MEM[0][0] ), 
        .QN(n209) );
  NAND2_X1 U3 ( .A1(n288), .A2(n3), .ZN(n370) );
  NAND2_X1 U9 ( .A1(n288), .A2(n15), .ZN(n374) );
  NAND2_X1 U15 ( .A1(n288), .A2(n21), .ZN(n378) );
  NAND2_X1 U21 ( .A1(n288), .A2(n27), .ZN(n382) );
  NAND2_X1 U27 ( .A1(n288), .A2(n33), .ZN(n386) );
  NAND2_X1 U33 ( .A1(n288), .A2(n39), .ZN(n390) );
  NAND2_X1 U39 ( .A1(n288), .A2(n45), .ZN(n394) );
  NAND2_X1 U45 ( .A1(n288), .A2(n51), .ZN(n398) );
  NAND2_X1 U51 ( .A1(n288), .A2(n57), .ZN(n402) );
  NAND2_X1 U57 ( .A1(n288), .A2(n63), .ZN(n406) );
  NAND2_X1 U63 ( .A1(n288), .A2(n69), .ZN(n410) );
  NAND2_X1 U69 ( .A1(n288), .A2(n75), .ZN(n414) );
  NAND2_X1 U75 ( .A1(n288), .A2(n81), .ZN(n418) );
  NAND2_X1 U81 ( .A1(n288), .A2(n87), .ZN(n422) );
  NAND2_X1 U87 ( .A1(n288), .A2(n93), .ZN(n426) );
  NAND2_X1 U93 ( .A1(n288), .A2(n99), .ZN(n430) );
  NAND2_X1 U99 ( .A1(n288), .A2(n105), .ZN(n434) );
  NAND2_X1 U105 ( .A1(n288), .A2(n111), .ZN(n438) );
  NAND2_X1 U111 ( .A1(n288), .A2(n117), .ZN(n442) );
  NAND2_X1 U117 ( .A1(n288), .A2(n123), .ZN(n446) );
  NAND2_X1 U123 ( .A1(n288), .A2(n129), .ZN(n450) );
  NAND2_X1 U129 ( .A1(n288), .A2(n135), .ZN(n454) );
  NAND2_X1 U135 ( .A1(n288), .A2(n141), .ZN(n458) );
  NAND2_X1 U141 ( .A1(n288), .A2(n147), .ZN(n462) );
  NAND2_X1 U147 ( .A1(n288), .A2(n153), .ZN(n466) );
  NAND2_X1 U153 ( .A1(n288), .A2(n159), .ZN(n470) );
  NAND2_X1 U159 ( .A1(n288), .A2(n165), .ZN(n474) );
  NAND2_X1 U165 ( .A1(n288), .A2(n171), .ZN(n478) );
  NAND2_X1 U171 ( .A1(n288), .A2(n177), .ZN(n482) );
  NAND2_X1 U177 ( .A1(n288), .A2(n183), .ZN(n486) );
  NAND2_X1 U183 ( .A1(n288), .A2(n189), .ZN(n490) );
  NAND2_X1 U189 ( .A1(n288), .A2(n195), .ZN(n494) );
  NAND2_X1 U264 ( .A1(ADDR[0]), .A2(n203), .ZN(n4) );
  NAND2_X1 U331 ( .A1(ADDR[1]), .A2(n206), .ZN(n6) );
  DFFRS_X1 \DATA_OUT_reg[31]  ( .D(1'b0), .CK(CLK), .RN(n493), .SN(n494), .Q(
        DATA_OUT[31]) );
  DFFRS_X1 \DATA_OUT_reg[30]  ( .D(1'b0), .CK(CLK), .RN(n489), .SN(n490), .Q(
        DATA_OUT[30]) );
  DFFRS_X1 \DATA_OUT_reg[29]  ( .D(1'b0), .CK(CLK), .RN(n485), .SN(n486), .Q(
        DATA_OUT[29]) );
  DFFRS_X1 \DATA_OUT_reg[28]  ( .D(1'b0), .CK(CLK), .RN(n481), .SN(n482), .Q(
        DATA_OUT[28]) );
  DFFRS_X1 \DATA_OUT_reg[27]  ( .D(1'b0), .CK(CLK), .RN(n477), .SN(n478), .Q(
        DATA_OUT[27]) );
  DFFRS_X1 \DATA_OUT_reg[26]  ( .D(1'b0), .CK(CLK), .RN(n473), .SN(n474), .Q(
        DATA_OUT[26]) );
  DFFRS_X1 \DATA_OUT_reg[25]  ( .D(1'b0), .CK(CLK), .RN(n469), .SN(n470), .Q(
        DATA_OUT[25]) );
  DFFRS_X1 \DATA_OUT_reg[24]  ( .D(1'b0), .CK(CLK), .RN(n465), .SN(n466), .Q(
        DATA_OUT[24]) );
  DFFRS_X1 \DATA_OUT_reg[23]  ( .D(1'b0), .CK(CLK), .RN(n461), .SN(n462), .Q(
        DATA_OUT[23]) );
  DFFRS_X1 \DATA_OUT_reg[22]  ( .D(1'b0), .CK(CLK), .RN(n457), .SN(n458), .Q(
        DATA_OUT[22]) );
  DFFRS_X1 \DATA_OUT_reg[21]  ( .D(1'b0), .CK(CLK), .RN(n453), .SN(n454), .Q(
        DATA_OUT[21]) );
  DFFRS_X1 \DATA_OUT_reg[20]  ( .D(1'b0), .CK(CLK), .RN(n449), .SN(n450), .Q(
        DATA_OUT[20]) );
  DFFRS_X1 \DATA_OUT_reg[19]  ( .D(1'b0), .CK(CLK), .RN(n445), .SN(n446), .Q(
        DATA_OUT[19]) );
  DFFRS_X1 \DATA_OUT_reg[18]  ( .D(1'b0), .CK(CLK), .RN(n441), .SN(n442), .Q(
        DATA_OUT[18]) );
  DFFRS_X1 \DATA_OUT_reg[17]  ( .D(1'b0), .CK(CLK), .RN(n437), .SN(n438), .Q(
        DATA_OUT[17]) );
  DFFRS_X1 \DATA_OUT_reg[16]  ( .D(1'b0), .CK(CLK), .RN(n433), .SN(n434), .Q(
        DATA_OUT[16]) );
  DFFRS_X1 \DATA_OUT_reg[15]  ( .D(1'b0), .CK(CLK), .RN(n429), .SN(n430), .Q(
        DATA_OUT[15]) );
  DFFRS_X1 \DATA_OUT_reg[14]  ( .D(1'b0), .CK(CLK), .RN(n425), .SN(n426), .Q(
        DATA_OUT[14]) );
  DFFRS_X1 \DATA_OUT_reg[13]  ( .D(1'b0), .CK(CLK), .RN(n421), .SN(n422), .Q(
        DATA_OUT[13]) );
  DFFRS_X1 \DATA_OUT_reg[12]  ( .D(1'b0), .CK(CLK), .RN(n417), .SN(n418), .Q(
        DATA_OUT[12]) );
  DFFRS_X1 \DATA_OUT_reg[11]  ( .D(1'b0), .CK(CLK), .RN(n413), .SN(n414), .Q(
        DATA_OUT[11]) );
  DFFRS_X1 \DATA_OUT_reg[10]  ( .D(1'b0), .CK(CLK), .RN(n409), .SN(n410), .Q(
        DATA_OUT[10]) );
  DFFRS_X1 \DATA_OUT_reg[9]  ( .D(1'b0), .CK(CLK), .RN(n405), .SN(n406), .Q(
        DATA_OUT[9]) );
  DFFRS_X1 \DATA_OUT_reg[8]  ( .D(1'b0), .CK(CLK), .RN(n401), .SN(n402), .Q(
        DATA_OUT[8]) );
  DFFRS_X1 \DATA_OUT_reg[7]  ( .D(1'b0), .CK(CLK), .RN(n397), .SN(n398), .Q(
        DATA_OUT[7]) );
  DFFRS_X1 \DATA_OUT_reg[6]  ( .D(1'b0), .CK(CLK), .RN(n393), .SN(n394), .Q(
        DATA_OUT[6]) );
  DFFRS_X1 \DATA_OUT_reg[5]  ( .D(1'b0), .CK(CLK), .RN(n389), .SN(n390), .Q(
        DATA_OUT[5]) );
  DFFRS_X1 \DATA_OUT_reg[4]  ( .D(1'b0), .CK(CLK), .RN(n385), .SN(n386), .Q(
        DATA_OUT[4]) );
  DFFRS_X1 \DATA_OUT_reg[3]  ( .D(1'b0), .CK(CLK), .RN(n381), .SN(n382), .Q(
        DATA_OUT[3]) );
  DFFRS_X1 \DATA_OUT_reg[2]  ( .D(1'b0), .CK(CLK), .RN(n377), .SN(n378), .Q(
        DATA_OUT[2]) );
  DFFRS_X1 \DATA_OUT_reg[1]  ( .D(1'b0), .CK(CLK), .RN(n373), .SN(n374), .Q(
        DATA_OUT[1]) );
  DFFRS_X1 \DATA_OUT_reg[0]  ( .D(1'b0), .CK(CLK), .RN(n369), .SN(n370), .Q(
        DATA_OUT[0]) );
  AND2_X1 U4 ( .A1(n300), .A2(n281), .ZN(n1) );
  INV_X1 U5 ( .A(n245), .ZN(n235) );
  INV_X1 U6 ( .A(n245), .ZN(n236) );
  BUF_X1 U7 ( .A(n1), .Z(n245) );
  INV_X1 U8 ( .A(n265), .ZN(n256) );
  BUF_X1 U10 ( .A(n1), .Z(n244) );
  BUF_X1 U11 ( .A(n1), .Z(n243) );
  BUF_X1 U12 ( .A(n1), .Z(n242) );
  BUF_X1 U13 ( .A(n1), .Z(n241) );
  BUF_X1 U14 ( .A(n1), .Z(n240) );
  BUF_X1 U16 ( .A(n1), .Z(n239) );
  BUF_X1 U17 ( .A(n1), .Z(n238) );
  BUF_X1 U18 ( .A(n1), .Z(n237) );
  INV_X1 U19 ( .A(n255), .ZN(n246) );
  INV_X1 U20 ( .A(n275), .ZN(n266) );
  BUF_X1 U22 ( .A(n202), .Z(n265) );
  BUF_X1 U23 ( .A(n205), .Z(n255) );
  BUF_X1 U24 ( .A(n11), .Z(n275) );
  BUF_X1 U25 ( .A(n202), .Z(n264) );
  BUF_X1 U26 ( .A(n202), .Z(n263) );
  BUF_X1 U28 ( .A(n202), .Z(n262) );
  BUF_X1 U29 ( .A(n202), .Z(n261) );
  BUF_X1 U30 ( .A(n202), .Z(n260) );
  BUF_X1 U31 ( .A(n202), .Z(n259) );
  BUF_X1 U32 ( .A(n202), .Z(n258) );
  BUF_X1 U34 ( .A(n202), .Z(n257) );
  BUF_X1 U35 ( .A(n205), .Z(n254) );
  BUF_X1 U36 ( .A(n205), .Z(n253) );
  BUF_X1 U37 ( .A(n205), .Z(n252) );
  BUF_X1 U38 ( .A(n205), .Z(n251) );
  BUF_X1 U40 ( .A(n205), .Z(n250) );
  BUF_X1 U41 ( .A(n205), .Z(n249) );
  BUF_X1 U42 ( .A(n205), .Z(n248) );
  BUF_X1 U43 ( .A(n205), .Z(n247) );
  BUF_X1 U44 ( .A(n11), .Z(n274) );
  BUF_X1 U46 ( .A(n11), .Z(n273) );
  BUF_X1 U47 ( .A(n11), .Z(n272) );
  BUF_X1 U48 ( .A(n11), .Z(n271) );
  BUF_X1 U49 ( .A(n11), .Z(n270) );
  BUF_X1 U50 ( .A(n11), .Z(n269) );
  BUF_X1 U52 ( .A(n11), .Z(n268) );
  BUF_X1 U53 ( .A(n11), .Z(n267) );
  NOR2_X1 U54 ( .A1(n288), .A2(n287), .ZN(n202) );
  NOR2_X1 U55 ( .A1(n288), .A2(n282), .ZN(n205) );
  BUF_X1 U56 ( .A(n9), .Z(n281) );
  INV_X1 U58 ( .A(n289), .ZN(n288) );
  NAND2_X1 U59 ( .A1(n300), .A2(n278), .ZN(n11) );
  BUF_X1 U60 ( .A(n9), .Z(n279) );
  BUF_X1 U61 ( .A(n9), .Z(n280) );
  NOR2_X1 U62 ( .A1(n203), .A2(n206), .ZN(n9) );
  BUF_X1 U64 ( .A(n4), .Z(n287) );
  BUF_X1 U65 ( .A(n6), .Z(n282) );
  BUF_X1 U66 ( .A(n10), .Z(n278) );
  BUF_X1 U67 ( .A(n4), .Z(n285) );
  BUF_X1 U68 ( .A(n4), .Z(n286) );
  BUF_X1 U70 ( .A(n10), .Z(n276) );
  BUF_X1 U71 ( .A(n10), .Z(n277) );
  BUF_X1 U72 ( .A(n6), .Z(n284) );
  BUF_X1 U73 ( .A(n6), .Z(n283) );
  OAI22_X1 U74 ( .A1(n12), .A2(n256), .B1(n264), .B2(n17), .ZN(n497) );
  OAI22_X1 U76 ( .A1(n19), .A2(n256), .B1(n264), .B2(n20), .ZN(n498) );
  OAI22_X1 U77 ( .A1(n25), .A2(n256), .B1(n264), .B2(n22), .ZN(n499) );
  OAI22_X1 U78 ( .A1(n31), .A2(n256), .B1(n264), .B2(n23), .ZN(n500) );
  OAI22_X1 U79 ( .A1(n37), .A2(n256), .B1(n263), .B2(n26), .ZN(n501) );
  OAI22_X1 U80 ( .A1(n43), .A2(n256), .B1(n263), .B2(n28), .ZN(n502) );
  OAI22_X1 U82 ( .A1(n49), .A2(n256), .B1(n263), .B2(n29), .ZN(n503) );
  OAI22_X1 U83 ( .A1(n55), .A2(n256), .B1(n263), .B2(n32), .ZN(n504) );
  OAI22_X1 U84 ( .A1(n61), .A2(n256), .B1(n262), .B2(n34), .ZN(n505) );
  OAI22_X1 U85 ( .A1(n67), .A2(n256), .B1(n262), .B2(n35), .ZN(n506) );
  OAI22_X1 U86 ( .A1(n73), .A2(n256), .B1(n262), .B2(n38), .ZN(n507) );
  OAI22_X1 U88 ( .A1(n79), .A2(n256), .B1(n262), .B2(n40), .ZN(n508) );
  OAI22_X1 U89 ( .A1(n85), .A2(n256), .B1(n261), .B2(n41), .ZN(n509) );
  OAI22_X1 U90 ( .A1(n91), .A2(n256), .B1(n261), .B2(n44), .ZN(n510) );
  OAI22_X1 U91 ( .A1(n97), .A2(n256), .B1(n261), .B2(n46), .ZN(n511) );
  OAI22_X1 U92 ( .A1(n103), .A2(n256), .B1(n261), .B2(n47), .ZN(n512) );
  OAI22_X1 U94 ( .A1(n109), .A2(n256), .B1(n260), .B2(n50), .ZN(n513) );
  OAI22_X1 U95 ( .A1(n115), .A2(n256), .B1(n260), .B2(n52), .ZN(n514) );
  OAI22_X1 U96 ( .A1(n121), .A2(n256), .B1(n260), .B2(n53), .ZN(n515) );
  OAI22_X1 U97 ( .A1(n127), .A2(n256), .B1(n260), .B2(n56), .ZN(n516) );
  OAI22_X1 U98 ( .A1(n133), .A2(n256), .B1(n259), .B2(n58), .ZN(n517) );
  OAI22_X1 U100 ( .A1(n139), .A2(n256), .B1(n259), .B2(n59), .ZN(n518) );
  OAI22_X1 U101 ( .A1(n145), .A2(n256), .B1(n259), .B2(n62), .ZN(n519) );
  OAI22_X1 U102 ( .A1(n151), .A2(n256), .B1(n259), .B2(n64), .ZN(n520) );
  OAI22_X1 U103 ( .A1(n157), .A2(n256), .B1(n258), .B2(n65), .ZN(n521) );
  OAI22_X1 U104 ( .A1(n163), .A2(n256), .B1(n258), .B2(n68), .ZN(n522) );
  OAI22_X1 U106 ( .A1(n169), .A2(n256), .B1(n258), .B2(n2), .ZN(n523) );
  OAI22_X1 U107 ( .A1(n175), .A2(n256), .B1(n258), .B2(n5), .ZN(n524) );
  OAI22_X1 U108 ( .A1(n181), .A2(n256), .B1(n257), .B2(n7), .ZN(n525) );
  OAI22_X1 U109 ( .A1(n187), .A2(n256), .B1(n257), .B2(n13), .ZN(n526) );
  OAI22_X1 U110 ( .A1(n193), .A2(n256), .B1(n257), .B2(n14), .ZN(n527) );
  OAI22_X1 U112 ( .A1(n199), .A2(n256), .B1(n257), .B2(n16), .ZN(n528) );
  OAI22_X1 U113 ( .A1(n12), .A2(n246), .B1(n254), .B2(n82), .ZN(n529) );
  OAI22_X1 U114 ( .A1(n19), .A2(n246), .B1(n254), .B2(n83), .ZN(n530) );
  OAI22_X1 U115 ( .A1(n25), .A2(n246), .B1(n254), .B2(n86), .ZN(n531) );
  OAI22_X1 U116 ( .A1(n31), .A2(n246), .B1(n254), .B2(n88), .ZN(n532) );
  OAI22_X1 U118 ( .A1(n37), .A2(n246), .B1(n253), .B2(n89), .ZN(n533) );
  OAI22_X1 U119 ( .A1(n43), .A2(n246), .B1(n253), .B2(n92), .ZN(n534) );
  OAI22_X1 U120 ( .A1(n49), .A2(n246), .B1(n253), .B2(n94), .ZN(n535) );
  OAI22_X1 U121 ( .A1(n55), .A2(n246), .B1(n253), .B2(n95), .ZN(n536) );
  OAI22_X1 U122 ( .A1(n61), .A2(n246), .B1(n252), .B2(n98), .ZN(n537) );
  OAI22_X1 U124 ( .A1(n67), .A2(n246), .B1(n252), .B2(n100), .ZN(n538) );
  OAI22_X1 U125 ( .A1(n73), .A2(n246), .B1(n252), .B2(n101), .ZN(n539) );
  OAI22_X1 U126 ( .A1(n79), .A2(n246), .B1(n252), .B2(n104), .ZN(n540) );
  OAI22_X1 U127 ( .A1(n85), .A2(n246), .B1(n251), .B2(n106), .ZN(n541) );
  OAI22_X1 U128 ( .A1(n91), .A2(n246), .B1(n251), .B2(n107), .ZN(n542) );
  OAI22_X1 U130 ( .A1(n97), .A2(n246), .B1(n251), .B2(n110), .ZN(n543) );
  OAI22_X1 U131 ( .A1(n103), .A2(n246), .B1(n251), .B2(n112), .ZN(n544) );
  OAI22_X1 U132 ( .A1(n109), .A2(n246), .B1(n250), .B2(n113), .ZN(n545) );
  OAI22_X1 U133 ( .A1(n115), .A2(n246), .B1(n250), .B2(n116), .ZN(n546) );
  OAI22_X1 U134 ( .A1(n121), .A2(n246), .B1(n250), .B2(n118), .ZN(n547) );
  OAI22_X1 U136 ( .A1(n127), .A2(n246), .B1(n250), .B2(n119), .ZN(n548) );
  OAI22_X1 U137 ( .A1(n133), .A2(n246), .B1(n249), .B2(n122), .ZN(n549) );
  OAI22_X1 U138 ( .A1(n139), .A2(n246), .B1(n249), .B2(n124), .ZN(n550) );
  OAI22_X1 U139 ( .A1(n145), .A2(n246), .B1(n249), .B2(n125), .ZN(n551) );
  OAI22_X1 U140 ( .A1(n151), .A2(n246), .B1(n249), .B2(n128), .ZN(n552) );
  OAI22_X1 U142 ( .A1(n157), .A2(n246), .B1(n248), .B2(n130), .ZN(n553) );
  OAI22_X1 U143 ( .A1(n163), .A2(n246), .B1(n248), .B2(n131), .ZN(n554) );
  OAI22_X1 U144 ( .A1(n169), .A2(n246), .B1(n248), .B2(n70), .ZN(n555) );
  OAI22_X1 U145 ( .A1(n175), .A2(n246), .B1(n248), .B2(n71), .ZN(n556) );
  OAI22_X1 U146 ( .A1(n181), .A2(n246), .B1(n247), .B2(n74), .ZN(n557) );
  OAI22_X1 U148 ( .A1(n187), .A2(n246), .B1(n247), .B2(n76), .ZN(n558) );
  OAI22_X1 U149 ( .A1(n193), .A2(n246), .B1(n247), .B2(n77), .ZN(n559) );
  OAI22_X1 U150 ( .A1(n199), .A2(n246), .B1(n247), .B2(n80), .ZN(n560) );
  INV_X1 U151 ( .A(ADDR[0]), .ZN(n206) );
  INV_X1 U152 ( .A(DATA_IN[0]), .ZN(n12) );
  INV_X1 U154 ( .A(DATA_IN[1]), .ZN(n19) );
  INV_X1 U155 ( .A(DATA_IN[2]), .ZN(n25) );
  INV_X1 U156 ( .A(DATA_IN[3]), .ZN(n31) );
  INV_X1 U157 ( .A(DATA_IN[4]), .ZN(n37) );
  INV_X1 U158 ( .A(DATA_IN[5]), .ZN(n43) );
  INV_X1 U160 ( .A(DATA_IN[6]), .ZN(n49) );
  INV_X1 U161 ( .A(DATA_IN[7]), .ZN(n55) );
  INV_X1 U162 ( .A(DATA_IN[8]), .ZN(n61) );
  INV_X1 U163 ( .A(DATA_IN[9]), .ZN(n67) );
  INV_X1 U164 ( .A(DATA_IN[10]), .ZN(n73) );
  INV_X1 U166 ( .A(DATA_IN[11]), .ZN(n79) );
  INV_X1 U167 ( .A(DATA_IN[12]), .ZN(n85) );
  INV_X1 U168 ( .A(DATA_IN[13]), .ZN(n91) );
  INV_X1 U169 ( .A(DATA_IN[14]), .ZN(n97) );
  INV_X1 U170 ( .A(DATA_IN[15]), .ZN(n103) );
  INV_X1 U172 ( .A(DATA_IN[16]), .ZN(n109) );
  INV_X1 U173 ( .A(DATA_IN[17]), .ZN(n115) );
  INV_X1 U174 ( .A(DATA_IN[18]), .ZN(n121) );
  INV_X1 U175 ( .A(DATA_IN[19]), .ZN(n127) );
  INV_X1 U176 ( .A(DATA_IN[20]), .ZN(n133) );
  INV_X1 U178 ( .A(DATA_IN[21]), .ZN(n139) );
  INV_X1 U179 ( .A(DATA_IN[22]), .ZN(n145) );
  INV_X1 U180 ( .A(DATA_IN[23]), .ZN(n151) );
  INV_X1 U181 ( .A(DATA_IN[24]), .ZN(n157) );
  INV_X1 U182 ( .A(DATA_IN[25]), .ZN(n163) );
  INV_X1 U184 ( .A(DATA_IN[26]), .ZN(n169) );
  INV_X1 U185 ( .A(DATA_IN[27]), .ZN(n175) );
  INV_X1 U186 ( .A(DATA_IN[28]), .ZN(n181) );
  INV_X1 U187 ( .A(DATA_IN[29]), .ZN(n187) );
  INV_X1 U188 ( .A(DATA_IN[30]), .ZN(n193) );
  INV_X1 U190 ( .A(DATA_IN[31]), .ZN(n199) );
  INV_X1 U191 ( .A(ADDR[1]), .ZN(n203) );
  NOR2_X1 U192 ( .A1(ADDR[0]), .A2(ADDR[1]), .ZN(n10) );
  OR2_X1 U193 ( .A1(n3), .A2(n289), .ZN(n369) );
  OR2_X1 U194 ( .A1(n195), .A2(n300), .ZN(n493) );
  OR2_X1 U195 ( .A1(n165), .A2(n298), .ZN(n473) );
  OR2_X1 U196 ( .A1(n171), .A2(n298), .ZN(n477) );
  OR2_X1 U197 ( .A1(n177), .A2(n299), .ZN(n481) );
  OR2_X1 U198 ( .A1(n183), .A2(n299), .ZN(n485) );
  OR2_X1 U199 ( .A1(n189), .A2(n299), .ZN(n489) );
  OR2_X1 U200 ( .A1(n15), .A2(n290), .ZN(n373) );
  OR2_X1 U201 ( .A1(n21), .A2(n290), .ZN(n377) );
  OR2_X1 U202 ( .A1(n27), .A2(n290), .ZN(n381) );
  OR2_X1 U203 ( .A1(n33), .A2(n291), .ZN(n385) );
  OR2_X1 U204 ( .A1(n39), .A2(n291), .ZN(n389) );
  OR2_X1 U205 ( .A1(n45), .A2(n291), .ZN(n393) );
  OR2_X1 U206 ( .A1(n51), .A2(n292), .ZN(n397) );
  OR2_X1 U207 ( .A1(n57), .A2(n292), .ZN(n401) );
  OR2_X1 U208 ( .A1(n63), .A2(n292), .ZN(n405) );
  OR2_X1 U209 ( .A1(n69), .A2(n293), .ZN(n409) );
  OR2_X1 U210 ( .A1(n75), .A2(n293), .ZN(n413) );
  OR2_X1 U211 ( .A1(n81), .A2(n293), .ZN(n417) );
  OR2_X1 U212 ( .A1(n87), .A2(n294), .ZN(n421) );
  OR2_X1 U213 ( .A1(n93), .A2(n294), .ZN(n425) );
  OR2_X1 U214 ( .A1(n99), .A2(n294), .ZN(n429) );
  OR2_X1 U215 ( .A1(n105), .A2(n295), .ZN(n433) );
  OR2_X1 U216 ( .A1(n111), .A2(n295), .ZN(n437) );
  OR2_X1 U217 ( .A1(n117), .A2(n295), .ZN(n441) );
  OR2_X1 U218 ( .A1(n123), .A2(n296), .ZN(n445) );
  OR2_X1 U219 ( .A1(n129), .A2(n296), .ZN(n449) );
  OR2_X1 U220 ( .A1(n135), .A2(n296), .ZN(n453) );
  OR2_X1 U221 ( .A1(n141), .A2(n297), .ZN(n457) );
  OR2_X1 U222 ( .A1(n147), .A2(n297), .ZN(n461) );
  OR2_X1 U223 ( .A1(n153), .A2(n297), .ZN(n465) );
  OR2_X1 U224 ( .A1(n159), .A2(n298), .ZN(n469) );
  OAI22_X1 U225 ( .A1(n268), .A2(n169), .B1(n266), .B2(n197), .ZN(n476) );
  OAI22_X1 U226 ( .A1(n268), .A2(n175), .B1(n266), .B2(n200), .ZN(n480) );
  OAI22_X1 U227 ( .A1(n267), .A2(n181), .B1(n266), .B2(n201), .ZN(n484) );
  OAI22_X1 U228 ( .A1(n267), .A2(n187), .B1(n266), .B2(n204), .ZN(n488) );
  OAI22_X1 U229 ( .A1(n267), .A2(n193), .B1(n266), .B2(n207), .ZN(n492) );
  OAI22_X1 U230 ( .A1(n267), .A2(n199), .B1(n266), .B2(n208), .ZN(n496) );
  OAI22_X1 U231 ( .A1(n274), .A2(n12), .B1(n266), .B2(n209), .ZN(n372) );
  OAI22_X1 U232 ( .A1(n274), .A2(n19), .B1(n266), .B2(n210), .ZN(n376) );
  OAI22_X1 U233 ( .A1(n274), .A2(n25), .B1(n266), .B2(n211), .ZN(n380) );
  OAI22_X1 U234 ( .A1(n274), .A2(n31), .B1(n266), .B2(n212), .ZN(n384) );
  OAI22_X1 U235 ( .A1(n273), .A2(n37), .B1(n266), .B2(n213), .ZN(n388) );
  OAI22_X1 U236 ( .A1(n273), .A2(n43), .B1(n266), .B2(n214), .ZN(n392) );
  OAI22_X1 U237 ( .A1(n273), .A2(n49), .B1(n266), .B2(n215), .ZN(n396) );
  OAI22_X1 U238 ( .A1(n273), .A2(n55), .B1(n266), .B2(n216), .ZN(n400) );
  OAI22_X1 U239 ( .A1(n272), .A2(n61), .B1(n266), .B2(n217), .ZN(n404) );
  OAI22_X1 U240 ( .A1(n272), .A2(n67), .B1(n266), .B2(n218), .ZN(n408) );
  OAI22_X1 U241 ( .A1(n272), .A2(n73), .B1(n266), .B2(n219), .ZN(n412) );
  OAI22_X1 U242 ( .A1(n272), .A2(n79), .B1(n266), .B2(n220), .ZN(n416) );
  OAI22_X1 U243 ( .A1(n271), .A2(n85), .B1(n266), .B2(n221), .ZN(n420) );
  OAI22_X1 U244 ( .A1(n271), .A2(n91), .B1(n266), .B2(n222), .ZN(n424) );
  OAI22_X1 U245 ( .A1(n271), .A2(n97), .B1(n266), .B2(n223), .ZN(n428) );
  OAI22_X1 U246 ( .A1(n271), .A2(n103), .B1(n266), .B2(n224), .ZN(n432) );
  OAI22_X1 U247 ( .A1(n270), .A2(n109), .B1(n266), .B2(n225), .ZN(n436) );
  OAI22_X1 U248 ( .A1(n270), .A2(n115), .B1(n266), .B2(n226), .ZN(n440) );
  OAI22_X1 U249 ( .A1(n270), .A2(n121), .B1(n266), .B2(n227), .ZN(n444) );
  OAI22_X1 U250 ( .A1(n270), .A2(n127), .B1(n266), .B2(n228), .ZN(n448) );
  OAI22_X1 U251 ( .A1(n269), .A2(n133), .B1(n266), .B2(n229), .ZN(n452) );
  OAI22_X1 U252 ( .A1(n269), .A2(n139), .B1(n266), .B2(n230), .ZN(n456) );
  OAI22_X1 U253 ( .A1(n269), .A2(n145), .B1(n266), .B2(n231), .ZN(n460) );
  OAI22_X1 U254 ( .A1(n269), .A2(n151), .B1(n266), .B2(n232), .ZN(n464) );
  OAI22_X1 U255 ( .A1(n268), .A2(n157), .B1(n266), .B2(n233), .ZN(n468) );
  OAI22_X1 U256 ( .A1(n268), .A2(n163), .B1(n266), .B2(n234), .ZN(n472) );
  OAI22_X1 U257 ( .A1(n12), .A2(n235), .B1(n244), .B2(n134), .ZN(n561) );
  OAI22_X1 U258 ( .A1(n19), .A2(n235), .B1(n244), .B2(n136), .ZN(n562) );
  OAI22_X1 U259 ( .A1(n25), .A2(n235), .B1(n244), .B2(n137), .ZN(n563) );
  OAI22_X1 U260 ( .A1(n31), .A2(n235), .B1(n244), .B2(n140), .ZN(n564) );
  OAI22_X1 U261 ( .A1(n37), .A2(n235), .B1(n243), .B2(n142), .ZN(n565) );
  OAI22_X1 U262 ( .A1(n43), .A2(n235), .B1(n243), .B2(n143), .ZN(n566) );
  OAI22_X1 U263 ( .A1(n49), .A2(n235), .B1(n243), .B2(n146), .ZN(n567) );
  OAI22_X1 U265 ( .A1(n55), .A2(n235), .B1(n243), .B2(n148), .ZN(n568) );
  OAI22_X1 U266 ( .A1(n61), .A2(n235), .B1(n242), .B2(n149), .ZN(n569) );
  OAI22_X1 U267 ( .A1(n67), .A2(n235), .B1(n242), .B2(n152), .ZN(n570) );
  OAI22_X1 U268 ( .A1(n73), .A2(n235), .B1(n242), .B2(n154), .ZN(n571) );
  OAI22_X1 U269 ( .A1(n79), .A2(n235), .B1(n242), .B2(n155), .ZN(n572) );
  OAI22_X1 U270 ( .A1(n85), .A2(n235), .B1(n241), .B2(n158), .ZN(n573) );
  OAI22_X1 U271 ( .A1(n91), .A2(n236), .B1(n241), .B2(n160), .ZN(n574) );
  OAI22_X1 U272 ( .A1(n97), .A2(n236), .B1(n241), .B2(n161), .ZN(n575) );
  OAI22_X1 U273 ( .A1(n103), .A2(n236), .B1(n241), .B2(n164), .ZN(n576) );
  OAI22_X1 U274 ( .A1(n109), .A2(n236), .B1(n240), .B2(n166), .ZN(n577) );
  OAI22_X1 U275 ( .A1(n115), .A2(n236), .B1(n240), .B2(n167), .ZN(n578) );
  OAI22_X1 U276 ( .A1(n121), .A2(n236), .B1(n240), .B2(n170), .ZN(n579) );
  OAI22_X1 U277 ( .A1(n127), .A2(n236), .B1(n240), .B2(n172), .ZN(n580) );
  OAI22_X1 U278 ( .A1(n133), .A2(n236), .B1(n239), .B2(n173), .ZN(n581) );
  OAI22_X1 U279 ( .A1(n139), .A2(n236), .B1(n239), .B2(n176), .ZN(n582) );
  OAI22_X1 U280 ( .A1(n145), .A2(n236), .B1(n239), .B2(n178), .ZN(n583) );
  OAI22_X1 U281 ( .A1(n151), .A2(n236), .B1(n239), .B2(n179), .ZN(n584) );
  OAI22_X1 U282 ( .A1(n157), .A2(n236), .B1(n238), .B2(n182), .ZN(n585) );
  OAI22_X1 U283 ( .A1(n163), .A2(n236), .B1(n238), .B2(n184), .ZN(n586) );
  OAI22_X1 U284 ( .A1(n169), .A2(n235), .B1(n238), .B2(n185), .ZN(n587) );
  OAI22_X1 U285 ( .A1(n175), .A2(n236), .B1(n238), .B2(n188), .ZN(n588) );
  OAI22_X1 U286 ( .A1(n181), .A2(n235), .B1(n237), .B2(n190), .ZN(n589) );
  OAI22_X1 U287 ( .A1(n187), .A2(n236), .B1(n237), .B2(n191), .ZN(n590) );
  OAI22_X1 U288 ( .A1(n193), .A2(n235), .B1(n237), .B2(n194), .ZN(n591) );
  OAI22_X1 U289 ( .A1(n199), .A2(n236), .B1(n237), .B2(n196), .ZN(n592) );
  OAI221_X1 U290 ( .B1(n287), .B2(n2), .C1(n282), .C2(n70), .A(n168), .ZN(n165) );
  AOI22_X1 U291 ( .A1(\CACHE_MEM[3][26] ), .A2(n281), .B1(\CACHE_MEM[0][26] ), 
        .B2(n278), .ZN(n168) );
  OAI221_X1 U292 ( .B1(n287), .B2(n5), .C1(n282), .C2(n71), .A(n174), .ZN(n171) );
  AOI22_X1 U293 ( .A1(\CACHE_MEM[3][27] ), .A2(n281), .B1(\CACHE_MEM[0][27] ), 
        .B2(n278), .ZN(n174) );
  OAI221_X1 U294 ( .B1(n287), .B2(n7), .C1(n282), .C2(n74), .A(n180), .ZN(n177) );
  AOI22_X1 U295 ( .A1(\CACHE_MEM[3][28] ), .A2(n281), .B1(\CACHE_MEM[0][28] ), 
        .B2(n278), .ZN(n180) );
  OAI221_X1 U296 ( .B1(n287), .B2(n13), .C1(n282), .C2(n76), .A(n186), .ZN(
        n183) );
  AOI22_X1 U297 ( .A1(\CACHE_MEM[3][29] ), .A2(n281), .B1(\CACHE_MEM[0][29] ), 
        .B2(n278), .ZN(n186) );
  OAI221_X1 U298 ( .B1(n287), .B2(n14), .C1(n282), .C2(n77), .A(n192), .ZN(
        n189) );
  AOI22_X1 U299 ( .A1(\CACHE_MEM[3][30] ), .A2(n281), .B1(\CACHE_MEM[0][30] ), 
        .B2(n278), .ZN(n192) );
  OAI221_X1 U300 ( .B1(n287), .B2(n16), .C1(n282), .C2(n80), .A(n198), .ZN(
        n195) );
  AOI22_X1 U301 ( .A1(\CACHE_MEM[3][31] ), .A2(n281), .B1(\CACHE_MEM[0][31] ), 
        .B2(n278), .ZN(n198) );
  OAI221_X1 U302 ( .B1(n285), .B2(n17), .C1(n284), .C2(n82), .A(n8), .ZN(n3)
         );
  AOI22_X1 U303 ( .A1(\CACHE_MEM[3][0] ), .A2(n279), .B1(\CACHE_MEM[0][0] ), 
        .B2(n276), .ZN(n8) );
  OAI221_X1 U304 ( .B1(n285), .B2(n20), .C1(n284), .C2(n83), .A(n18), .ZN(n15)
         );
  AOI22_X1 U305 ( .A1(\CACHE_MEM[3][1] ), .A2(n279), .B1(\CACHE_MEM[0][1] ), 
        .B2(n276), .ZN(n18) );
  OAI221_X1 U306 ( .B1(n285), .B2(n22), .C1(n284), .C2(n86), .A(n24), .ZN(n21)
         );
  AOI22_X1 U307 ( .A1(\CACHE_MEM[3][2] ), .A2(n279), .B1(\CACHE_MEM[0][2] ), 
        .B2(n276), .ZN(n24) );
  OAI221_X1 U308 ( .B1(n285), .B2(n23), .C1(n284), .C2(n88), .A(n30), .ZN(n27)
         );
  AOI22_X1 U309 ( .A1(\CACHE_MEM[3][3] ), .A2(n279), .B1(\CACHE_MEM[0][3] ), 
        .B2(n276), .ZN(n30) );
  OAI221_X1 U310 ( .B1(n285), .B2(n26), .C1(n284), .C2(n89), .A(n36), .ZN(n33)
         );
  AOI22_X1 U311 ( .A1(\CACHE_MEM[3][4] ), .A2(n279), .B1(\CACHE_MEM[0][4] ), 
        .B2(n276), .ZN(n36) );
  OAI221_X1 U312 ( .B1(n285), .B2(n28), .C1(n283), .C2(n92), .A(n42), .ZN(n39)
         );
  AOI22_X1 U313 ( .A1(\CACHE_MEM[3][5] ), .A2(n279), .B1(\CACHE_MEM[0][5] ), 
        .B2(n276), .ZN(n42) );
  OAI221_X1 U314 ( .B1(n285), .B2(n29), .C1(n283), .C2(n94), .A(n48), .ZN(n45)
         );
  AOI22_X1 U315 ( .A1(\CACHE_MEM[3][6] ), .A2(n279), .B1(\CACHE_MEM[0][6] ), 
        .B2(n276), .ZN(n48) );
  OAI221_X1 U316 ( .B1(n285), .B2(n32), .C1(n283), .C2(n95), .A(n54), .ZN(n51)
         );
  AOI22_X1 U317 ( .A1(\CACHE_MEM[3][7] ), .A2(n279), .B1(\CACHE_MEM[0][7] ), 
        .B2(n276), .ZN(n54) );
  OAI221_X1 U318 ( .B1(n285), .B2(n34), .C1(n283), .C2(n98), .A(n60), .ZN(n57)
         );
  AOI22_X1 U319 ( .A1(\CACHE_MEM[3][8] ), .A2(n279), .B1(\CACHE_MEM[0][8] ), 
        .B2(n276), .ZN(n60) );
  OAI221_X1 U320 ( .B1(n285), .B2(n35), .C1(n283), .C2(n100), .A(n66), .ZN(n63) );
  AOI22_X1 U321 ( .A1(\CACHE_MEM[3][9] ), .A2(n279), .B1(\CACHE_MEM[0][9] ), 
        .B2(n276), .ZN(n66) );
  OAI221_X1 U322 ( .B1(n285), .B2(n38), .C1(n283), .C2(n101), .A(n72), .ZN(n69) );
  AOI22_X1 U323 ( .A1(\CACHE_MEM[3][10] ), .A2(n279), .B1(\CACHE_MEM[0][10] ), 
        .B2(n276), .ZN(n72) );
  OAI221_X1 U324 ( .B1(n285), .B2(n40), .C1(n283), .C2(n104), .A(n78), .ZN(n75) );
  AOI22_X1 U325 ( .A1(\CACHE_MEM[3][11] ), .A2(n279), .B1(\CACHE_MEM[0][11] ), 
        .B2(n276), .ZN(n78) );
  OAI221_X1 U326 ( .B1(n285), .B2(n41), .C1(n283), .C2(n106), .A(n84), .ZN(n81) );
  AOI22_X1 U327 ( .A1(\CACHE_MEM[3][12] ), .A2(n279), .B1(\CACHE_MEM[0][12] ), 
        .B2(n276), .ZN(n84) );
  OAI221_X1 U328 ( .B1(n286), .B2(n44), .C1(n283), .C2(n107), .A(n90), .ZN(n87) );
  AOI22_X1 U329 ( .A1(\CACHE_MEM[3][13] ), .A2(n280), .B1(\CACHE_MEM[0][13] ), 
        .B2(n277), .ZN(n90) );
  OAI221_X1 U330 ( .B1(n286), .B2(n46), .C1(n283), .C2(n110), .A(n96), .ZN(n93) );
  AOI22_X1 U332 ( .A1(\CACHE_MEM[3][14] ), .A2(n280), .B1(\CACHE_MEM[0][14] ), 
        .B2(n277), .ZN(n96) );
  OAI221_X1 U333 ( .B1(n286), .B2(n47), .C1(n283), .C2(n112), .A(n102), .ZN(
        n99) );
  AOI22_X1 U334 ( .A1(\CACHE_MEM[3][15] ), .A2(n280), .B1(\CACHE_MEM[0][15] ), 
        .B2(n277), .ZN(n102) );
  OAI221_X1 U335 ( .B1(n286), .B2(n50), .C1(n283), .C2(n113), .A(n108), .ZN(
        n105) );
  AOI22_X1 U336 ( .A1(\CACHE_MEM[3][16] ), .A2(n280), .B1(\CACHE_MEM[0][16] ), 
        .B2(n277), .ZN(n108) );
  OAI221_X1 U337 ( .B1(n286), .B2(n52), .C1(n283), .C2(n116), .A(n114), .ZN(
        n111) );
  AOI22_X1 U338 ( .A1(\CACHE_MEM[3][17] ), .A2(n280), .B1(\CACHE_MEM[0][17] ), 
        .B2(n277), .ZN(n114) );
  OAI221_X1 U339 ( .B1(n286), .B2(n53), .C1(n283), .C2(n118), .A(n120), .ZN(
        n117) );
  AOI22_X1 U340 ( .A1(\CACHE_MEM[3][18] ), .A2(n280), .B1(\CACHE_MEM[0][18] ), 
        .B2(n277), .ZN(n120) );
  OAI221_X1 U341 ( .B1(n286), .B2(n56), .C1(n282), .C2(n119), .A(n126), .ZN(
        n123) );
  AOI22_X1 U342 ( .A1(\CACHE_MEM[3][19] ), .A2(n280), .B1(\CACHE_MEM[0][19] ), 
        .B2(n277), .ZN(n126) );
  OAI221_X1 U343 ( .B1(n286), .B2(n58), .C1(n282), .C2(n122), .A(n132), .ZN(
        n129) );
  AOI22_X1 U344 ( .A1(\CACHE_MEM[3][20] ), .A2(n280), .B1(\CACHE_MEM[0][20] ), 
        .B2(n277), .ZN(n132) );
  OAI221_X1 U345 ( .B1(n286), .B2(n59), .C1(n282), .C2(n124), .A(n138), .ZN(
        n135) );
  AOI22_X1 U346 ( .A1(\CACHE_MEM[3][21] ), .A2(n280), .B1(\CACHE_MEM[0][21] ), 
        .B2(n277), .ZN(n138) );
  OAI221_X1 U347 ( .B1(n286), .B2(n62), .C1(n282), .C2(n125), .A(n144), .ZN(
        n141) );
  AOI22_X1 U348 ( .A1(\CACHE_MEM[3][22] ), .A2(n280), .B1(\CACHE_MEM[0][22] ), 
        .B2(n277), .ZN(n144) );
  OAI221_X1 U349 ( .B1(n286), .B2(n64), .C1(n282), .C2(n128), .A(n150), .ZN(
        n147) );
  AOI22_X1 U350 ( .A1(\CACHE_MEM[3][23] ), .A2(n280), .B1(\CACHE_MEM[0][23] ), 
        .B2(n277), .ZN(n150) );
  OAI221_X1 U351 ( .B1(n286), .B2(n65), .C1(n282), .C2(n130), .A(n156), .ZN(
        n153) );
  AOI22_X1 U352 ( .A1(\CACHE_MEM[3][24] ), .A2(n280), .B1(\CACHE_MEM[0][24] ), 
        .B2(n277), .ZN(n156) );
  OAI221_X1 U353 ( .B1(n286), .B2(n68), .C1(n282), .C2(n131), .A(n162), .ZN(
        n159) );
  AOI22_X1 U354 ( .A1(\CACHE_MEM[3][25] ), .A2(n280), .B1(\CACHE_MEM[0][25] ), 
        .B2(n277), .ZN(n162) );
  CLKBUF_X1 U355 ( .A(WE), .Z(n289) );
  CLKBUF_X1 U356 ( .A(WE), .Z(n290) );
  CLKBUF_X1 U357 ( .A(WE), .Z(n291) );
  CLKBUF_X1 U358 ( .A(WE), .Z(n292) );
  CLKBUF_X1 U359 ( .A(WE), .Z(n293) );
  CLKBUF_X1 U360 ( .A(WE), .Z(n294) );
  CLKBUF_X1 U361 ( .A(WE), .Z(n295) );
  CLKBUF_X1 U362 ( .A(WE), .Z(n296) );
  CLKBUF_X1 U363 ( .A(WE), .Z(n297) );
  CLKBUF_X1 U364 ( .A(WE), .Z(n298) );
  CLKBUF_X1 U365 ( .A(WE), .Z(n299) );
  CLKBUF_X1 U366 ( .A(WE), .Z(n300) );
endmodule


module MUX21_GEN_N2 ( A, B, SEL, Y );
  input [1:0] A;
  input [1:0] B;
  output [1:0] Y;
  input SEL;
  wire   SB;
  wire   [1:0] Y1;
  wire   [1:0] Y2;

  INV_1_120 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_1023 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_1022 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_1021 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_1020 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_1019 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_1018 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
endmodule


module SYNC_COUNTER_2BIT ( EN, RST, CLK, COUNT );
  output [1:0] COUNT;
  input EN, RST, CLK;


  FFT_2 FFT_1 ( .T(1'b1), .CLK(CLK), .EN(EN), .RST(RST), .Q(COUNT[0]) );
  FFT_1 FFT_2 ( .T(COUNT[0]), .CLK(CLK), .EN(EN), .RST(RST), .Q(COUNT[1]) );
endmodule


module BPU_ENCODER ( A, Y );
  input [3:0] A;
  output [1:0] Y;


  OR_GATE_309 OR_1 ( .A(A[1]), .B(A[3]), .Y(Y[0]) );
  OR_GATE_308 OR_2 ( .A(A[2]), .B(A[3]), .Y(Y[1]) );
endmodule


module N_OR_N4 ( A, Y );
  input [3:0] A;
  output Y;


  OR4_X1 U1 ( .A1(A[1]), .A2(A[0]), .A3(A[3]), .A4(A[2]), .ZN(Y) );
endmodule


module EQU_COMPARATOR_N32_0 ( A, B, Y );
  input [31:0] A;
  input [31:0] B;
  output Y;

  wire   [31:0] L;

  XNOR_GATE_160 XNORING_0 ( .A(A[0]), .B(B[0]), .Y(L[0]) );
  XNOR_GATE_159 XNORING_1 ( .A(A[1]), .B(B[1]), .Y(L[1]) );
  XNOR_GATE_158 XNORING_2 ( .A(A[2]), .B(B[2]), .Y(L[2]) );
  XNOR_GATE_157 XNORING_3 ( .A(A[3]), .B(B[3]), .Y(L[3]) );
  XNOR_GATE_156 XNORING_4 ( .A(A[4]), .B(B[4]), .Y(L[4]) );
  XNOR_GATE_155 XNORING_5 ( .A(A[5]), .B(B[5]), .Y(L[5]) );
  XNOR_GATE_154 XNORING_6 ( .A(A[6]), .B(B[6]), .Y(L[6]) );
  XNOR_GATE_153 XNORING_7 ( .A(A[7]), .B(B[7]), .Y(L[7]) );
  XNOR_GATE_152 XNORING_8 ( .A(A[8]), .B(B[8]), .Y(L[8]) );
  XNOR_GATE_151 XNORING_9 ( .A(A[9]), .B(B[9]), .Y(L[9]) );
  XNOR_GATE_150 XNORING_10 ( .A(A[10]), .B(B[10]), .Y(L[10]) );
  XNOR_GATE_149 XNORING_11 ( .A(A[11]), .B(B[11]), .Y(L[11]) );
  XNOR_GATE_148 XNORING_12 ( .A(A[12]), .B(B[12]), .Y(L[12]) );
  XNOR_GATE_147 XNORING_13 ( .A(A[13]), .B(B[13]), .Y(L[13]) );
  XNOR_GATE_146 XNORING_14 ( .A(A[14]), .B(B[14]), .Y(L[14]) );
  XNOR_GATE_145 XNORING_15 ( .A(A[15]), .B(B[15]), .Y(L[15]) );
  XNOR_GATE_144 XNORING_16 ( .A(A[16]), .B(B[16]), .Y(L[16]) );
  XNOR_GATE_143 XNORING_17 ( .A(A[17]), .B(B[17]), .Y(L[17]) );
  XNOR_GATE_142 XNORING_18 ( .A(A[18]), .B(B[18]), .Y(L[18]) );
  XNOR_GATE_141 XNORING_19 ( .A(A[19]), .B(B[19]), .Y(L[19]) );
  XNOR_GATE_140 XNORING_20 ( .A(A[20]), .B(B[20]), .Y(L[20]) );
  XNOR_GATE_139 XNORING_21 ( .A(A[21]), .B(B[21]), .Y(L[21]) );
  XNOR_GATE_138 XNORING_22 ( .A(A[22]), .B(B[22]), .Y(L[22]) );
  XNOR_GATE_137 XNORING_23 ( .A(A[23]), .B(B[23]), .Y(L[23]) );
  XNOR_GATE_136 XNORING_24 ( .A(A[24]), .B(B[24]), .Y(L[24]) );
  XNOR_GATE_135 XNORING_25 ( .A(A[25]), .B(B[25]), .Y(L[25]) );
  XNOR_GATE_134 XNORING_26 ( .A(A[26]), .B(B[26]), .Y(L[26]) );
  XNOR_GATE_133 XNORING_27 ( .A(A[27]), .B(B[27]), .Y(L[27]) );
  XNOR_GATE_132 XNORING_28 ( .A(A[28]), .B(B[28]), .Y(L[28]) );
  XNOR_GATE_131 XNORING_29 ( .A(A[29]), .B(B[29]), .Y(L[29]) );
  XNOR_GATE_130 XNORING_30 ( .A(A[30]), .B(B[30]), .Y(L[30]) );
  XNOR_GATE_129 XNORING_31 ( .A(A[31]), .B(B[31]), .Y(L[31]) );
  N_AND_N32_0 ANDING ( .A(L), .Y(Y) );
endmodule


module CAM_BPU_N32_SET_BIT2 ( ADDR, RST, WE, DATA_IN, ADDR_OUT_1, ADDR_OUT_2, 
        ADDR_OUT_3, ADDR_OUT_4, VALID_1, VALID_2, VALID_3, VALID_4 );
  input [1:0] ADDR;
  input [31:0] DATA_IN;
  output [31:0] ADDR_OUT_1;
  output [31:0] ADDR_OUT_2;
  output [31:0] ADDR_OUT_3;
  output [31:0] ADDR_OUT_4;
  input RST, WE;
  output VALID_1, VALID_2, VALID_3, VALID_4;
  wire   \CAM_MEM[3][31] , \CAM_MEM[3][30] , \CAM_MEM[3][29] ,
         \CAM_MEM[3][28] , \CAM_MEM[3][27] , \CAM_MEM[3][26] ,
         \CAM_MEM[3][25] , \CAM_MEM[3][24] , \CAM_MEM[3][23] ,
         \CAM_MEM[3][22] , \CAM_MEM[3][21] , \CAM_MEM[3][20] ,
         \CAM_MEM[3][19] , \CAM_MEM[3][18] , \CAM_MEM[3][17] ,
         \CAM_MEM[3][16] , \CAM_MEM[3][15] , \CAM_MEM[3][14] ,
         \CAM_MEM[3][13] , \CAM_MEM[3][12] , \CAM_MEM[3][11] ,
         \CAM_MEM[3][10] , \CAM_MEM[3][9] , \CAM_MEM[3][8] , \CAM_MEM[3][7] ,
         \CAM_MEM[3][6] , \CAM_MEM[3][5] , \CAM_MEM[3][4] , \CAM_MEM[3][3] ,
         \CAM_MEM[3][2] , \CAM_MEM[3][1] , \CAM_MEM[3][0] , \CAM_MEM[2][31] ,
         \CAM_MEM[2][30] , \CAM_MEM[2][29] , \CAM_MEM[2][28] ,
         \CAM_MEM[2][27] , \CAM_MEM[2][26] , \CAM_MEM[2][25] ,
         \CAM_MEM[2][24] , \CAM_MEM[2][23] , \CAM_MEM[2][22] ,
         \CAM_MEM[2][21] , \CAM_MEM[2][20] , \CAM_MEM[2][19] ,
         \CAM_MEM[2][18] , \CAM_MEM[2][17] , \CAM_MEM[2][16] ,
         \CAM_MEM[2][15] , \CAM_MEM[2][14] , \CAM_MEM[2][13] ,
         \CAM_MEM[2][12] , \CAM_MEM[2][11] , \CAM_MEM[2][10] , \CAM_MEM[2][9] ,
         \CAM_MEM[2][8] , \CAM_MEM[2][7] , \CAM_MEM[2][6] , \CAM_MEM[2][5] ,
         \CAM_MEM[2][4] , \CAM_MEM[2][3] , \CAM_MEM[2][2] , \CAM_MEM[2][1] ,
         \CAM_MEM[2][0] , \CAM_MEM[1][31] , \CAM_MEM[1][30] , \CAM_MEM[1][29] ,
         \CAM_MEM[1][28] , \CAM_MEM[1][27] , \CAM_MEM[1][26] ,
         \CAM_MEM[1][25] , \CAM_MEM[1][24] , \CAM_MEM[1][23] ,
         \CAM_MEM[1][22] , \CAM_MEM[1][21] , \CAM_MEM[1][20] ,
         \CAM_MEM[1][19] , \CAM_MEM[1][18] , \CAM_MEM[1][17] ,
         \CAM_MEM[1][16] , \CAM_MEM[1][15] , \CAM_MEM[1][14] ,
         \CAM_MEM[1][13] , \CAM_MEM[1][12] , \CAM_MEM[1][11] ,
         \CAM_MEM[1][10] , \CAM_MEM[1][9] , \CAM_MEM[1][8] , \CAM_MEM[1][7] ,
         \CAM_MEM[1][6] , \CAM_MEM[1][5] , \CAM_MEM[1][4] , \CAM_MEM[1][3] ,
         \CAM_MEM[1][2] , \CAM_MEM[1][1] , \CAM_MEM[1][0] , \CAM_MEM[0][31] ,
         \CAM_MEM[0][30] , \CAM_MEM[0][29] , \CAM_MEM[0][28] ,
         \CAM_MEM[0][27] , \CAM_MEM[0][26] , \CAM_MEM[0][25] ,
         \CAM_MEM[0][24] , \CAM_MEM[0][23] , \CAM_MEM[0][22] ,
         \CAM_MEM[0][21] , \CAM_MEM[0][20] , \CAM_MEM[0][19] ,
         \CAM_MEM[0][18] , \CAM_MEM[0][17] , \CAM_MEM[0][16] ,
         \CAM_MEM[0][15] , \CAM_MEM[0][14] , \CAM_MEM[0][13] ,
         \CAM_MEM[0][12] , \CAM_MEM[0][11] , \CAM_MEM[0][10] , \CAM_MEM[0][9] ,
         \CAM_MEM[0][8] , \CAM_MEM[0][7] , \CAM_MEM[0][6] , \CAM_MEM[0][5] ,
         \CAM_MEM[0][4] , \CAM_MEM[0][3] , \CAM_MEM[0][2] , \CAM_MEM[0][1] ,
         \CAM_MEM[0][0] , N190, N222, N254, N286, N417, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n1, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23;
  wire   [3:0] VALID_BIT;

  DLL_X1 \VALID_BIT_reg[3]  ( .D(n23), .GN(n7), .Q(VALID_BIT[3]) );
  DLL_X1 \VALID_BIT_reg[2]  ( .D(n23), .GN(n10), .Q(VALID_BIT[2]) );
  DLH_X1 VALID_3_reg ( .G(n22), .D(VALID_BIT[2]), .Q(VALID_3) );
  DLL_X1 \VALID_BIT_reg[1]  ( .D(n23), .GN(n11), .Q(VALID_BIT[1]) );
  DLL_X1 \VALID_BIT_reg[0]  ( .D(n23), .GN(n12), .Q(VALID_BIT[0]) );
  DLH_X1 VALID_4_reg ( .G(n22), .D(VALID_BIT[3]), .Q(VALID_4) );
  DLH_X1 \CAM_MEM_reg[3][31]  ( .G(N286), .D(DATA_IN[31]), .Q(\CAM_MEM[3][31] ) );
  DLH_X1 \CAM_MEM_reg[3][30]  ( .G(N286), .D(DATA_IN[30]), .Q(\CAM_MEM[3][30] ) );
  DLH_X1 \CAM_MEM_reg[3][29]  ( .G(N286), .D(DATA_IN[29]), .Q(\CAM_MEM[3][29] ) );
  DLH_X1 \CAM_MEM_reg[3][28]  ( .G(N286), .D(DATA_IN[28]), .Q(\CAM_MEM[3][28] ) );
  DLH_X1 \CAM_MEM_reg[3][27]  ( .G(N286), .D(DATA_IN[27]), .Q(\CAM_MEM[3][27] ) );
  DLH_X1 \CAM_MEM_reg[3][26]  ( .G(N286), .D(DATA_IN[26]), .Q(\CAM_MEM[3][26] ) );
  DLH_X1 \CAM_MEM_reg[3][25]  ( .G(N286), .D(DATA_IN[25]), .Q(\CAM_MEM[3][25] ) );
  DLH_X1 \CAM_MEM_reg[3][24]  ( .G(N286), .D(DATA_IN[24]), .Q(\CAM_MEM[3][24] ) );
  DLH_X1 \CAM_MEM_reg[3][23]  ( .G(N286), .D(DATA_IN[23]), .Q(\CAM_MEM[3][23] ) );
  DLH_X1 \CAM_MEM_reg[3][22]  ( .G(N286), .D(DATA_IN[22]), .Q(\CAM_MEM[3][22] ) );
  DLH_X1 \CAM_MEM_reg[3][21]  ( .G(N286), .D(DATA_IN[21]), .Q(\CAM_MEM[3][21] ) );
  DLH_X1 \CAM_MEM_reg[3][20]  ( .G(N286), .D(DATA_IN[20]), .Q(\CAM_MEM[3][20] ) );
  DLH_X1 \CAM_MEM_reg[3][19]  ( .G(N286), .D(DATA_IN[19]), .Q(\CAM_MEM[3][19] ) );
  DLH_X1 \CAM_MEM_reg[3][18]  ( .G(N286), .D(DATA_IN[18]), .Q(\CAM_MEM[3][18] ) );
  DLH_X1 \CAM_MEM_reg[3][17]  ( .G(N286), .D(DATA_IN[17]), .Q(\CAM_MEM[3][17] ) );
  DLH_X1 \CAM_MEM_reg[3][16]  ( .G(N286), .D(DATA_IN[16]), .Q(\CAM_MEM[3][16] ) );
  DLH_X1 \CAM_MEM_reg[3][15]  ( .G(N286), .D(DATA_IN[15]), .Q(\CAM_MEM[3][15] ) );
  DLH_X1 \CAM_MEM_reg[3][14]  ( .G(N286), .D(DATA_IN[14]), .Q(\CAM_MEM[3][14] ) );
  DLH_X1 \CAM_MEM_reg[3][13]  ( .G(N286), .D(DATA_IN[13]), .Q(\CAM_MEM[3][13] ) );
  DLH_X1 \CAM_MEM_reg[3][12]  ( .G(N286), .D(DATA_IN[12]), .Q(\CAM_MEM[3][12] ) );
  DLH_X1 \CAM_MEM_reg[3][11]  ( .G(N286), .D(DATA_IN[11]), .Q(\CAM_MEM[3][11] ) );
  DLH_X1 \CAM_MEM_reg[3][10]  ( .G(N286), .D(DATA_IN[10]), .Q(\CAM_MEM[3][10] ) );
  DLH_X1 \CAM_MEM_reg[3][9]  ( .G(N286), .D(DATA_IN[9]), .Q(\CAM_MEM[3][9] )
         );
  DLH_X1 \CAM_MEM_reg[3][8]  ( .G(N286), .D(DATA_IN[8]), .Q(\CAM_MEM[3][8] )
         );
  DLH_X1 \CAM_MEM_reg[3][7]  ( .G(N286), .D(DATA_IN[7]), .Q(\CAM_MEM[3][7] )
         );
  DLH_X1 \CAM_MEM_reg[3][6]  ( .G(N286), .D(DATA_IN[6]), .Q(\CAM_MEM[3][6] )
         );
  DLH_X1 \CAM_MEM_reg[3][5]  ( .G(N286), .D(DATA_IN[5]), .Q(\CAM_MEM[3][5] )
         );
  DLH_X1 \CAM_MEM_reg[3][4]  ( .G(N286), .D(DATA_IN[4]), .Q(\CAM_MEM[3][4] )
         );
  DLH_X1 \CAM_MEM_reg[3][3]  ( .G(N286), .D(DATA_IN[3]), .Q(\CAM_MEM[3][3] )
         );
  DLH_X1 \CAM_MEM_reg[3][2]  ( .G(N286), .D(DATA_IN[2]), .Q(\CAM_MEM[3][2] )
         );
  DLH_X1 \CAM_MEM_reg[3][1]  ( .G(N286), .D(DATA_IN[1]), .Q(\CAM_MEM[3][1] )
         );
  DLH_X1 \CAM_MEM_reg[3][0]  ( .G(N286), .D(DATA_IN[0]), .Q(\CAM_MEM[3][0] )
         );
  DLH_X1 \CAM_MEM_reg[2][31]  ( .G(N254), .D(DATA_IN[31]), .Q(\CAM_MEM[2][31] ) );
  DLH_X1 \CAM_MEM_reg[2][30]  ( .G(N254), .D(DATA_IN[30]), .Q(\CAM_MEM[2][30] ) );
  DLH_X1 \CAM_MEM_reg[2][29]  ( .G(N254), .D(DATA_IN[29]), .Q(\CAM_MEM[2][29] ) );
  DLH_X1 \CAM_MEM_reg[2][28]  ( .G(N254), .D(DATA_IN[28]), .Q(\CAM_MEM[2][28] ) );
  DLH_X1 \CAM_MEM_reg[2][27]  ( .G(N254), .D(DATA_IN[27]), .Q(\CAM_MEM[2][27] ) );
  DLH_X1 \CAM_MEM_reg[2][26]  ( .G(N254), .D(DATA_IN[26]), .Q(\CAM_MEM[2][26] ) );
  DLH_X1 \CAM_MEM_reg[2][25]  ( .G(N254), .D(DATA_IN[25]), .Q(\CAM_MEM[2][25] ) );
  DLH_X1 \CAM_MEM_reg[2][24]  ( .G(N254), .D(DATA_IN[24]), .Q(\CAM_MEM[2][24] ) );
  DLH_X1 \CAM_MEM_reg[2][23]  ( .G(N254), .D(DATA_IN[23]), .Q(\CAM_MEM[2][23] ) );
  DLH_X1 \CAM_MEM_reg[2][22]  ( .G(N254), .D(DATA_IN[22]), .Q(\CAM_MEM[2][22] ) );
  DLH_X1 \CAM_MEM_reg[2][21]  ( .G(N254), .D(DATA_IN[21]), .Q(\CAM_MEM[2][21] ) );
  DLH_X1 \CAM_MEM_reg[2][20]  ( .G(N254), .D(DATA_IN[20]), .Q(\CAM_MEM[2][20] ) );
  DLH_X1 \CAM_MEM_reg[2][19]  ( .G(N254), .D(DATA_IN[19]), .Q(\CAM_MEM[2][19] ) );
  DLH_X1 \CAM_MEM_reg[2][18]  ( .G(N254), .D(DATA_IN[18]), .Q(\CAM_MEM[2][18] ) );
  DLH_X1 \CAM_MEM_reg[2][17]  ( .G(N254), .D(DATA_IN[17]), .Q(\CAM_MEM[2][17] ) );
  DLH_X1 \CAM_MEM_reg[2][16]  ( .G(N254), .D(DATA_IN[16]), .Q(\CAM_MEM[2][16] ) );
  DLH_X1 \CAM_MEM_reg[2][15]  ( .G(N254), .D(DATA_IN[15]), .Q(\CAM_MEM[2][15] ) );
  DLH_X1 \CAM_MEM_reg[2][14]  ( .G(N254), .D(DATA_IN[14]), .Q(\CAM_MEM[2][14] ) );
  DLH_X1 \CAM_MEM_reg[2][13]  ( .G(N254), .D(DATA_IN[13]), .Q(\CAM_MEM[2][13] ) );
  DLH_X1 \CAM_MEM_reg[2][12]  ( .G(N254), .D(DATA_IN[12]), .Q(\CAM_MEM[2][12] ) );
  DLH_X1 \CAM_MEM_reg[2][11]  ( .G(N254), .D(DATA_IN[11]), .Q(\CAM_MEM[2][11] ) );
  DLH_X1 \CAM_MEM_reg[2][10]  ( .G(N254), .D(DATA_IN[10]), .Q(\CAM_MEM[2][10] ) );
  DLH_X1 \CAM_MEM_reg[2][9]  ( .G(N254), .D(DATA_IN[9]), .Q(\CAM_MEM[2][9] )
         );
  DLH_X1 \CAM_MEM_reg[2][8]  ( .G(N254), .D(DATA_IN[8]), .Q(\CAM_MEM[2][8] )
         );
  DLH_X1 \CAM_MEM_reg[2][7]  ( .G(N254), .D(DATA_IN[7]), .Q(\CAM_MEM[2][7] )
         );
  DLH_X1 \CAM_MEM_reg[2][6]  ( .G(N254), .D(DATA_IN[6]), .Q(\CAM_MEM[2][6] )
         );
  DLH_X1 \CAM_MEM_reg[2][5]  ( .G(N254), .D(DATA_IN[5]), .Q(\CAM_MEM[2][5] )
         );
  DLH_X1 \CAM_MEM_reg[2][4]  ( .G(N254), .D(DATA_IN[4]), .Q(\CAM_MEM[2][4] )
         );
  DLH_X1 \CAM_MEM_reg[2][3]  ( .G(N254), .D(DATA_IN[3]), .Q(\CAM_MEM[2][3] )
         );
  DLH_X1 \CAM_MEM_reg[2][2]  ( .G(N254), .D(DATA_IN[2]), .Q(\CAM_MEM[2][2] )
         );
  DLH_X1 \CAM_MEM_reg[2][1]  ( .G(N254), .D(DATA_IN[1]), .Q(\CAM_MEM[2][1] )
         );
  DLH_X1 \CAM_MEM_reg[2][0]  ( .G(N254), .D(DATA_IN[0]), .Q(\CAM_MEM[2][0] )
         );
  DLH_X1 \CAM_MEM_reg[1][31]  ( .G(N222), .D(DATA_IN[31]), .Q(\CAM_MEM[1][31] ) );
  DLH_X1 \CAM_MEM_reg[1][30]  ( .G(N222), .D(DATA_IN[30]), .Q(\CAM_MEM[1][30] ) );
  DLH_X1 \CAM_MEM_reg[1][29]  ( .G(N222), .D(DATA_IN[29]), .Q(\CAM_MEM[1][29] ) );
  DLH_X1 \CAM_MEM_reg[1][28]  ( .G(N222), .D(DATA_IN[28]), .Q(\CAM_MEM[1][28] ) );
  DLH_X1 \CAM_MEM_reg[1][27]  ( .G(N222), .D(DATA_IN[27]), .Q(\CAM_MEM[1][27] ) );
  DLH_X1 \CAM_MEM_reg[1][26]  ( .G(N222), .D(DATA_IN[26]), .Q(\CAM_MEM[1][26] ) );
  DLH_X1 \CAM_MEM_reg[1][25]  ( .G(N222), .D(DATA_IN[25]), .Q(\CAM_MEM[1][25] ) );
  DLH_X1 \CAM_MEM_reg[1][24]  ( .G(N222), .D(DATA_IN[24]), .Q(\CAM_MEM[1][24] ) );
  DLH_X1 \CAM_MEM_reg[1][23]  ( .G(N222), .D(DATA_IN[23]), .Q(\CAM_MEM[1][23] ) );
  DLH_X1 \CAM_MEM_reg[1][22]  ( .G(N222), .D(DATA_IN[22]), .Q(\CAM_MEM[1][22] ) );
  DLH_X1 \CAM_MEM_reg[1][21]  ( .G(N222), .D(DATA_IN[21]), .Q(\CAM_MEM[1][21] ) );
  DLH_X1 \CAM_MEM_reg[1][20]  ( .G(N222), .D(DATA_IN[20]), .Q(\CAM_MEM[1][20] ) );
  DLH_X1 \CAM_MEM_reg[1][19]  ( .G(N222), .D(DATA_IN[19]), .Q(\CAM_MEM[1][19] ) );
  DLH_X1 \CAM_MEM_reg[1][18]  ( .G(N222), .D(DATA_IN[18]), .Q(\CAM_MEM[1][18] ) );
  DLH_X1 \CAM_MEM_reg[1][17]  ( .G(N222), .D(DATA_IN[17]), .Q(\CAM_MEM[1][17] ) );
  DLH_X1 \CAM_MEM_reg[1][16]  ( .G(N222), .D(DATA_IN[16]), .Q(\CAM_MEM[1][16] ) );
  DLH_X1 \CAM_MEM_reg[1][15]  ( .G(N222), .D(DATA_IN[15]), .Q(\CAM_MEM[1][15] ) );
  DLH_X1 \CAM_MEM_reg[1][14]  ( .G(N222), .D(DATA_IN[14]), .Q(\CAM_MEM[1][14] ) );
  DLH_X1 \CAM_MEM_reg[1][13]  ( .G(N222), .D(DATA_IN[13]), .Q(\CAM_MEM[1][13] ) );
  DLH_X1 \CAM_MEM_reg[1][12]  ( .G(N222), .D(DATA_IN[12]), .Q(\CAM_MEM[1][12] ) );
  DLH_X1 \CAM_MEM_reg[1][11]  ( .G(N222), .D(DATA_IN[11]), .Q(\CAM_MEM[1][11] ) );
  DLH_X1 \CAM_MEM_reg[1][10]  ( .G(N222), .D(DATA_IN[10]), .Q(\CAM_MEM[1][10] ) );
  DLH_X1 \CAM_MEM_reg[1][9]  ( .G(N222), .D(DATA_IN[9]), .Q(\CAM_MEM[1][9] )
         );
  DLH_X1 \CAM_MEM_reg[1][8]  ( .G(N222), .D(DATA_IN[8]), .Q(\CAM_MEM[1][8] )
         );
  DLH_X1 \CAM_MEM_reg[1][7]  ( .G(N222), .D(DATA_IN[7]), .Q(\CAM_MEM[1][7] )
         );
  DLH_X1 \CAM_MEM_reg[1][6]  ( .G(N222), .D(DATA_IN[6]), .Q(\CAM_MEM[1][6] )
         );
  DLH_X1 \CAM_MEM_reg[1][5]  ( .G(N222), .D(DATA_IN[5]), .Q(\CAM_MEM[1][5] )
         );
  DLH_X1 \CAM_MEM_reg[1][4]  ( .G(N222), .D(DATA_IN[4]), .Q(\CAM_MEM[1][4] )
         );
  DLH_X1 \CAM_MEM_reg[1][3]  ( .G(N222), .D(DATA_IN[3]), .Q(\CAM_MEM[1][3] )
         );
  DLH_X1 \CAM_MEM_reg[1][2]  ( .G(N222), .D(DATA_IN[2]), .Q(\CAM_MEM[1][2] )
         );
  DLH_X1 \CAM_MEM_reg[1][1]  ( .G(N222), .D(DATA_IN[1]), .Q(\CAM_MEM[1][1] )
         );
  DLH_X1 \CAM_MEM_reg[1][0]  ( .G(N222), .D(DATA_IN[0]), .Q(\CAM_MEM[1][0] )
         );
  DLH_X1 \CAM_MEM_reg[0][31]  ( .G(N190), .D(DATA_IN[31]), .Q(\CAM_MEM[0][31] ) );
  DLH_X1 \CAM_MEM_reg[0][30]  ( .G(N190), .D(DATA_IN[30]), .Q(\CAM_MEM[0][30] ) );
  DLH_X1 \CAM_MEM_reg[0][29]  ( .G(N190), .D(DATA_IN[29]), .Q(\CAM_MEM[0][29] ) );
  DLH_X1 \CAM_MEM_reg[0][28]  ( .G(N190), .D(DATA_IN[28]), .Q(\CAM_MEM[0][28] ) );
  DLH_X1 \CAM_MEM_reg[0][27]  ( .G(N190), .D(DATA_IN[27]), .Q(\CAM_MEM[0][27] ) );
  DLH_X1 \CAM_MEM_reg[0][26]  ( .G(N190), .D(DATA_IN[26]), .Q(\CAM_MEM[0][26] ) );
  DLH_X1 \CAM_MEM_reg[0][25]  ( .G(N190), .D(DATA_IN[25]), .Q(\CAM_MEM[0][25] ) );
  DLH_X1 \CAM_MEM_reg[0][24]  ( .G(N190), .D(DATA_IN[24]), .Q(\CAM_MEM[0][24] ) );
  DLH_X1 \CAM_MEM_reg[0][23]  ( .G(N190), .D(DATA_IN[23]), .Q(\CAM_MEM[0][23] ) );
  DLH_X1 \CAM_MEM_reg[0][22]  ( .G(N190), .D(DATA_IN[22]), .Q(\CAM_MEM[0][22] ) );
  DLH_X1 \CAM_MEM_reg[0][21]  ( .G(N190), .D(DATA_IN[21]), .Q(\CAM_MEM[0][21] ) );
  DLH_X1 \CAM_MEM_reg[0][20]  ( .G(N190), .D(DATA_IN[20]), .Q(\CAM_MEM[0][20] ) );
  DLH_X1 \CAM_MEM_reg[0][19]  ( .G(N190), .D(DATA_IN[19]), .Q(\CAM_MEM[0][19] ) );
  DLH_X1 \CAM_MEM_reg[0][18]  ( .G(N190), .D(DATA_IN[18]), .Q(\CAM_MEM[0][18] ) );
  DLH_X1 \CAM_MEM_reg[0][17]  ( .G(N190), .D(DATA_IN[17]), .Q(\CAM_MEM[0][17] ) );
  DLH_X1 \CAM_MEM_reg[0][16]  ( .G(N190), .D(DATA_IN[16]), .Q(\CAM_MEM[0][16] ) );
  DLH_X1 \CAM_MEM_reg[0][15]  ( .G(N190), .D(DATA_IN[15]), .Q(\CAM_MEM[0][15] ) );
  DLH_X1 \CAM_MEM_reg[0][14]  ( .G(N190), .D(DATA_IN[14]), .Q(\CAM_MEM[0][14] ) );
  DLH_X1 \CAM_MEM_reg[0][13]  ( .G(N190), .D(DATA_IN[13]), .Q(\CAM_MEM[0][13] ) );
  DLH_X1 \CAM_MEM_reg[0][12]  ( .G(N190), .D(DATA_IN[12]), .Q(\CAM_MEM[0][12] ) );
  DLH_X1 \CAM_MEM_reg[0][11]  ( .G(N190), .D(DATA_IN[11]), .Q(\CAM_MEM[0][11] ) );
  DLH_X1 \CAM_MEM_reg[0][10]  ( .G(N190), .D(DATA_IN[10]), .Q(\CAM_MEM[0][10] ) );
  DLH_X1 \CAM_MEM_reg[0][9]  ( .G(N190), .D(DATA_IN[9]), .Q(\CAM_MEM[0][9] )
         );
  DLH_X1 \CAM_MEM_reg[0][8]  ( .G(N190), .D(DATA_IN[8]), .Q(\CAM_MEM[0][8] )
         );
  DLH_X1 \CAM_MEM_reg[0][7]  ( .G(N190), .D(DATA_IN[7]), .Q(\CAM_MEM[0][7] )
         );
  DLH_X1 \CAM_MEM_reg[0][6]  ( .G(N190), .D(DATA_IN[6]), .Q(\CAM_MEM[0][6] )
         );
  DLH_X1 \CAM_MEM_reg[0][5]  ( .G(N190), .D(DATA_IN[5]), .Q(\CAM_MEM[0][5] )
         );
  DLH_X1 \CAM_MEM_reg[0][4]  ( .G(N190), .D(DATA_IN[4]), .Q(\CAM_MEM[0][4] )
         );
  DLH_X1 \CAM_MEM_reg[0][3]  ( .G(N190), .D(DATA_IN[3]), .Q(\CAM_MEM[0][3] )
         );
  DLH_X1 \CAM_MEM_reg[0][2]  ( .G(N190), .D(DATA_IN[2]), .Q(\CAM_MEM[0][2] )
         );
  DLH_X1 \CAM_MEM_reg[0][1]  ( .G(N190), .D(DATA_IN[1]), .Q(\CAM_MEM[0][1] )
         );
  DLH_X1 \CAM_MEM_reg[0][0]  ( .G(N190), .D(DATA_IN[0]), .Q(\CAM_MEM[0][0] )
         );
  DLH_X1 \ADDR_OUT_1_reg[31]  ( .G(n21), .D(\CAM_MEM[0][31] ), .Q(
        ADDR_OUT_1[31]) );
  DLH_X1 \ADDR_OUT_1_reg[30]  ( .G(n21), .D(\CAM_MEM[0][30] ), .Q(
        ADDR_OUT_1[30]) );
  DLH_X1 \ADDR_OUT_1_reg[29]  ( .G(n21), .D(\CAM_MEM[0][29] ), .Q(
        ADDR_OUT_1[29]) );
  DLH_X1 \ADDR_OUT_1_reg[28]  ( .G(n21), .D(\CAM_MEM[0][28] ), .Q(
        ADDR_OUT_1[28]) );
  DLH_X1 \ADDR_OUT_1_reg[27]  ( .G(n21), .D(\CAM_MEM[0][27] ), .Q(
        ADDR_OUT_1[27]) );
  DLH_X1 \ADDR_OUT_1_reg[26]  ( .G(n21), .D(\CAM_MEM[0][26] ), .Q(
        ADDR_OUT_1[26]) );
  DLH_X1 \ADDR_OUT_1_reg[25]  ( .G(n21), .D(\CAM_MEM[0][25] ), .Q(
        ADDR_OUT_1[25]) );
  DLH_X1 \ADDR_OUT_1_reg[24]  ( .G(n21), .D(\CAM_MEM[0][24] ), .Q(
        ADDR_OUT_1[24]) );
  DLH_X1 \ADDR_OUT_1_reg[23]  ( .G(n21), .D(\CAM_MEM[0][23] ), .Q(
        ADDR_OUT_1[23]) );
  DLH_X1 \ADDR_OUT_1_reg[22]  ( .G(n21), .D(\CAM_MEM[0][22] ), .Q(
        ADDR_OUT_1[22]) );
  DLH_X1 \ADDR_OUT_1_reg[21]  ( .G(n21), .D(\CAM_MEM[0][21] ), .Q(
        ADDR_OUT_1[21]) );
  DLH_X1 \ADDR_OUT_1_reg[20]  ( .G(n21), .D(\CAM_MEM[0][20] ), .Q(
        ADDR_OUT_1[20]) );
  DLH_X1 \ADDR_OUT_1_reg[19]  ( .G(n21), .D(\CAM_MEM[0][19] ), .Q(
        ADDR_OUT_1[19]) );
  DLH_X1 \ADDR_OUT_1_reg[18]  ( .G(n20), .D(\CAM_MEM[0][18] ), .Q(
        ADDR_OUT_1[18]) );
  DLH_X1 \ADDR_OUT_1_reg[17]  ( .G(n20), .D(\CAM_MEM[0][17] ), .Q(
        ADDR_OUT_1[17]) );
  DLH_X1 \ADDR_OUT_1_reg[16]  ( .G(n20), .D(\CAM_MEM[0][16] ), .Q(
        ADDR_OUT_1[16]) );
  DLH_X1 \ADDR_OUT_1_reg[15]  ( .G(n20), .D(\CAM_MEM[0][15] ), .Q(
        ADDR_OUT_1[15]) );
  DLH_X1 \ADDR_OUT_1_reg[14]  ( .G(n20), .D(\CAM_MEM[0][14] ), .Q(
        ADDR_OUT_1[14]) );
  DLH_X1 \ADDR_OUT_1_reg[13]  ( .G(n20), .D(\CAM_MEM[0][13] ), .Q(
        ADDR_OUT_1[13]) );
  DLH_X1 \ADDR_OUT_1_reg[12]  ( .G(n20), .D(\CAM_MEM[0][12] ), .Q(
        ADDR_OUT_1[12]) );
  DLH_X1 \ADDR_OUT_1_reg[11]  ( .G(n20), .D(\CAM_MEM[0][11] ), .Q(
        ADDR_OUT_1[11]) );
  DLH_X1 \ADDR_OUT_1_reg[10]  ( .G(n20), .D(\CAM_MEM[0][10] ), .Q(
        ADDR_OUT_1[10]) );
  DLH_X1 \ADDR_OUT_1_reg[9]  ( .G(n20), .D(\CAM_MEM[0][9] ), .Q(ADDR_OUT_1[9])
         );
  DLH_X1 \ADDR_OUT_1_reg[8]  ( .G(n20), .D(\CAM_MEM[0][8] ), .Q(ADDR_OUT_1[8])
         );
  DLH_X1 \ADDR_OUT_1_reg[7]  ( .G(n20), .D(\CAM_MEM[0][7] ), .Q(ADDR_OUT_1[7])
         );
  DLH_X1 \ADDR_OUT_1_reg[6]  ( .G(n20), .D(\CAM_MEM[0][6] ), .Q(ADDR_OUT_1[6])
         );
  DLH_X1 \ADDR_OUT_1_reg[5]  ( .G(n19), .D(\CAM_MEM[0][5] ), .Q(ADDR_OUT_1[5])
         );
  DLH_X1 \ADDR_OUT_1_reg[4]  ( .G(n19), .D(\CAM_MEM[0][4] ), .Q(ADDR_OUT_1[4])
         );
  DLH_X1 \ADDR_OUT_1_reg[3]  ( .G(n19), .D(\CAM_MEM[0][3] ), .Q(ADDR_OUT_1[3])
         );
  DLH_X1 \ADDR_OUT_1_reg[2]  ( .G(n19), .D(\CAM_MEM[0][2] ), .Q(ADDR_OUT_1[2])
         );
  DLH_X1 \ADDR_OUT_1_reg[1]  ( .G(n19), .D(\CAM_MEM[0][1] ), .Q(ADDR_OUT_1[1])
         );
  DLH_X1 \ADDR_OUT_1_reg[0]  ( .G(n19), .D(\CAM_MEM[0][0] ), .Q(ADDR_OUT_1[0])
         );
  DLH_X1 \ADDR_OUT_2_reg[31]  ( .G(n19), .D(\CAM_MEM[1][31] ), .Q(
        ADDR_OUT_2[31]) );
  DLH_X1 \ADDR_OUT_2_reg[30]  ( .G(n19), .D(\CAM_MEM[1][30] ), .Q(
        ADDR_OUT_2[30]) );
  DLH_X1 \ADDR_OUT_2_reg[29]  ( .G(n19), .D(\CAM_MEM[1][29] ), .Q(
        ADDR_OUT_2[29]) );
  DLH_X1 \ADDR_OUT_2_reg[28]  ( .G(n19), .D(\CAM_MEM[1][28] ), .Q(
        ADDR_OUT_2[28]) );
  DLH_X1 \ADDR_OUT_2_reg[27]  ( .G(n19), .D(\CAM_MEM[1][27] ), .Q(
        ADDR_OUT_2[27]) );
  DLH_X1 \ADDR_OUT_2_reg[26]  ( .G(n19), .D(\CAM_MEM[1][26] ), .Q(
        ADDR_OUT_2[26]) );
  DLH_X1 \ADDR_OUT_2_reg[25]  ( .G(n19), .D(\CAM_MEM[1][25] ), .Q(
        ADDR_OUT_2[25]) );
  DLH_X1 \ADDR_OUT_2_reg[24]  ( .G(n18), .D(\CAM_MEM[1][24] ), .Q(
        ADDR_OUT_2[24]) );
  DLH_X1 \ADDR_OUT_2_reg[23]  ( .G(n18), .D(\CAM_MEM[1][23] ), .Q(
        ADDR_OUT_2[23]) );
  DLH_X1 \ADDR_OUT_2_reg[22]  ( .G(n18), .D(\CAM_MEM[1][22] ), .Q(
        ADDR_OUT_2[22]) );
  DLH_X1 \ADDR_OUT_2_reg[21]  ( .G(n18), .D(\CAM_MEM[1][21] ), .Q(
        ADDR_OUT_2[21]) );
  DLH_X1 \ADDR_OUT_2_reg[20]  ( .G(n18), .D(\CAM_MEM[1][20] ), .Q(
        ADDR_OUT_2[20]) );
  DLH_X1 \ADDR_OUT_2_reg[19]  ( .G(n18), .D(\CAM_MEM[1][19] ), .Q(
        ADDR_OUT_2[19]) );
  DLH_X1 \ADDR_OUT_2_reg[18]  ( .G(n18), .D(\CAM_MEM[1][18] ), .Q(
        ADDR_OUT_2[18]) );
  DLH_X1 \ADDR_OUT_2_reg[17]  ( .G(n18), .D(\CAM_MEM[1][17] ), .Q(
        ADDR_OUT_2[17]) );
  DLH_X1 \ADDR_OUT_2_reg[16]  ( .G(n18), .D(\CAM_MEM[1][16] ), .Q(
        ADDR_OUT_2[16]) );
  DLH_X1 \ADDR_OUT_2_reg[15]  ( .G(n18), .D(\CAM_MEM[1][15] ), .Q(
        ADDR_OUT_2[15]) );
  DLH_X1 \ADDR_OUT_2_reg[14]  ( .G(n18), .D(\CAM_MEM[1][14] ), .Q(
        ADDR_OUT_2[14]) );
  DLH_X1 \ADDR_OUT_2_reg[13]  ( .G(n18), .D(\CAM_MEM[1][13] ), .Q(
        ADDR_OUT_2[13]) );
  DLH_X1 \ADDR_OUT_2_reg[12]  ( .G(n18), .D(\CAM_MEM[1][12] ), .Q(
        ADDR_OUT_2[12]) );
  DLH_X1 \ADDR_OUT_2_reg[11]  ( .G(n17), .D(\CAM_MEM[1][11] ), .Q(
        ADDR_OUT_2[11]) );
  DLH_X1 \ADDR_OUT_2_reg[10]  ( .G(n17), .D(\CAM_MEM[1][10] ), .Q(
        ADDR_OUT_2[10]) );
  DLH_X1 \ADDR_OUT_2_reg[9]  ( .G(n17), .D(\CAM_MEM[1][9] ), .Q(ADDR_OUT_2[9])
         );
  DLH_X1 \ADDR_OUT_2_reg[8]  ( .G(n17), .D(\CAM_MEM[1][8] ), .Q(ADDR_OUT_2[8])
         );
  DLH_X1 \ADDR_OUT_2_reg[7]  ( .G(n17), .D(\CAM_MEM[1][7] ), .Q(ADDR_OUT_2[7])
         );
  DLH_X1 \ADDR_OUT_2_reg[6]  ( .G(n17), .D(\CAM_MEM[1][6] ), .Q(ADDR_OUT_2[6])
         );
  DLH_X1 \ADDR_OUT_2_reg[5]  ( .G(n17), .D(\CAM_MEM[1][5] ), .Q(ADDR_OUT_2[5])
         );
  DLH_X1 \ADDR_OUT_2_reg[4]  ( .G(n17), .D(\CAM_MEM[1][4] ), .Q(ADDR_OUT_2[4])
         );
  DLH_X1 \ADDR_OUT_2_reg[3]  ( .G(n17), .D(\CAM_MEM[1][3] ), .Q(ADDR_OUT_2[3])
         );
  DLH_X1 \ADDR_OUT_2_reg[2]  ( .G(n17), .D(\CAM_MEM[1][2] ), .Q(ADDR_OUT_2[2])
         );
  DLH_X1 \ADDR_OUT_2_reg[1]  ( .G(n17), .D(\CAM_MEM[1][1] ), .Q(ADDR_OUT_2[1])
         );
  DLH_X1 \ADDR_OUT_2_reg[0]  ( .G(n17), .D(\CAM_MEM[1][0] ), .Q(ADDR_OUT_2[0])
         );
  DLH_X1 \ADDR_OUT_3_reg[31]  ( .G(n17), .D(\CAM_MEM[2][31] ), .Q(
        ADDR_OUT_3[31]) );
  DLH_X1 \ADDR_OUT_3_reg[30]  ( .G(n16), .D(\CAM_MEM[2][30] ), .Q(
        ADDR_OUT_3[30]) );
  DLH_X1 \ADDR_OUT_3_reg[29]  ( .G(n16), .D(\CAM_MEM[2][29] ), .Q(
        ADDR_OUT_3[29]) );
  DLH_X1 \ADDR_OUT_3_reg[28]  ( .G(n16), .D(\CAM_MEM[2][28] ), .Q(
        ADDR_OUT_3[28]) );
  DLH_X1 \ADDR_OUT_3_reg[27]  ( .G(n16), .D(\CAM_MEM[2][27] ), .Q(
        ADDR_OUT_3[27]) );
  DLH_X1 \ADDR_OUT_3_reg[26]  ( .G(n16), .D(\CAM_MEM[2][26] ), .Q(
        ADDR_OUT_3[26]) );
  DLH_X1 \ADDR_OUT_3_reg[25]  ( .G(n16), .D(\CAM_MEM[2][25] ), .Q(
        ADDR_OUT_3[25]) );
  DLH_X1 \ADDR_OUT_3_reg[24]  ( .G(n16), .D(\CAM_MEM[2][24] ), .Q(
        ADDR_OUT_3[24]) );
  DLH_X1 \ADDR_OUT_3_reg[23]  ( .G(n16), .D(\CAM_MEM[2][23] ), .Q(
        ADDR_OUT_3[23]) );
  DLH_X1 \ADDR_OUT_3_reg[22]  ( .G(n16), .D(\CAM_MEM[2][22] ), .Q(
        ADDR_OUT_3[22]) );
  DLH_X1 \ADDR_OUT_3_reg[21]  ( .G(n16), .D(\CAM_MEM[2][21] ), .Q(
        ADDR_OUT_3[21]) );
  DLH_X1 \ADDR_OUT_3_reg[20]  ( .G(n16), .D(\CAM_MEM[2][20] ), .Q(
        ADDR_OUT_3[20]) );
  DLH_X1 \ADDR_OUT_3_reg[19]  ( .G(n16), .D(\CAM_MEM[2][19] ), .Q(
        ADDR_OUT_3[19]) );
  DLH_X1 \ADDR_OUT_3_reg[18]  ( .G(n16), .D(\CAM_MEM[2][18] ), .Q(
        ADDR_OUT_3[18]) );
  DLH_X1 \ADDR_OUT_3_reg[17]  ( .G(n15), .D(\CAM_MEM[2][17] ), .Q(
        ADDR_OUT_3[17]) );
  DLH_X1 \ADDR_OUT_3_reg[16]  ( .G(n15), .D(\CAM_MEM[2][16] ), .Q(
        ADDR_OUT_3[16]) );
  DLH_X1 \ADDR_OUT_3_reg[15]  ( .G(n15), .D(\CAM_MEM[2][15] ), .Q(
        ADDR_OUT_3[15]) );
  DLH_X1 \ADDR_OUT_3_reg[14]  ( .G(n15), .D(\CAM_MEM[2][14] ), .Q(
        ADDR_OUT_3[14]) );
  DLH_X1 \ADDR_OUT_3_reg[13]  ( .G(n15), .D(\CAM_MEM[2][13] ), .Q(
        ADDR_OUT_3[13]) );
  DLH_X1 \ADDR_OUT_3_reg[12]  ( .G(n15), .D(\CAM_MEM[2][12] ), .Q(
        ADDR_OUT_3[12]) );
  DLH_X1 \ADDR_OUT_3_reg[11]  ( .G(n15), .D(\CAM_MEM[2][11] ), .Q(
        ADDR_OUT_3[11]) );
  DLH_X1 \ADDR_OUT_3_reg[10]  ( .G(n15), .D(\CAM_MEM[2][10] ), .Q(
        ADDR_OUT_3[10]) );
  DLH_X1 \ADDR_OUT_3_reg[9]  ( .G(n15), .D(\CAM_MEM[2][9] ), .Q(ADDR_OUT_3[9])
         );
  DLH_X1 \ADDR_OUT_3_reg[8]  ( .G(n15), .D(\CAM_MEM[2][8] ), .Q(ADDR_OUT_3[8])
         );
  DLH_X1 \ADDR_OUT_3_reg[7]  ( .G(n15), .D(\CAM_MEM[2][7] ), .Q(ADDR_OUT_3[7])
         );
  DLH_X1 \ADDR_OUT_3_reg[6]  ( .G(n15), .D(\CAM_MEM[2][6] ), .Q(ADDR_OUT_3[6])
         );
  DLH_X1 \ADDR_OUT_3_reg[5]  ( .G(n15), .D(\CAM_MEM[2][5] ), .Q(ADDR_OUT_3[5])
         );
  DLH_X1 \ADDR_OUT_3_reg[4]  ( .G(n14), .D(\CAM_MEM[2][4] ), .Q(ADDR_OUT_3[4])
         );
  DLH_X1 \ADDR_OUT_3_reg[3]  ( .G(n14), .D(\CAM_MEM[2][3] ), .Q(ADDR_OUT_3[3])
         );
  DLH_X1 \ADDR_OUT_3_reg[2]  ( .G(n14), .D(\CAM_MEM[2][2] ), .Q(ADDR_OUT_3[2])
         );
  DLH_X1 \ADDR_OUT_3_reg[1]  ( .G(n14), .D(\CAM_MEM[2][1] ), .Q(ADDR_OUT_3[1])
         );
  DLH_X1 \ADDR_OUT_3_reg[0]  ( .G(n14), .D(\CAM_MEM[2][0] ), .Q(ADDR_OUT_3[0])
         );
  DLH_X1 \ADDR_OUT_4_reg[31]  ( .G(n14), .D(\CAM_MEM[3][31] ), .Q(
        ADDR_OUT_4[31]) );
  DLH_X1 \ADDR_OUT_4_reg[30]  ( .G(n14), .D(\CAM_MEM[3][30] ), .Q(
        ADDR_OUT_4[30]) );
  DLH_X1 \ADDR_OUT_4_reg[29]  ( .G(n14), .D(\CAM_MEM[3][29] ), .Q(
        ADDR_OUT_4[29]) );
  DLH_X1 \ADDR_OUT_4_reg[28]  ( .G(n14), .D(\CAM_MEM[3][28] ), .Q(
        ADDR_OUT_4[28]) );
  DLH_X1 \ADDR_OUT_4_reg[27]  ( .G(n14), .D(\CAM_MEM[3][27] ), .Q(
        ADDR_OUT_4[27]) );
  DLH_X1 \ADDR_OUT_4_reg[26]  ( .G(n14), .D(\CAM_MEM[3][26] ), .Q(
        ADDR_OUT_4[26]) );
  DLH_X1 \ADDR_OUT_4_reg[25]  ( .G(n14), .D(\CAM_MEM[3][25] ), .Q(
        ADDR_OUT_4[25]) );
  DLH_X1 \ADDR_OUT_4_reg[24]  ( .G(n14), .D(\CAM_MEM[3][24] ), .Q(
        ADDR_OUT_4[24]) );
  DLH_X1 \ADDR_OUT_4_reg[23]  ( .G(n13), .D(\CAM_MEM[3][23] ), .Q(
        ADDR_OUT_4[23]) );
  DLH_X1 \ADDR_OUT_4_reg[22]  ( .G(n13), .D(\CAM_MEM[3][22] ), .Q(
        ADDR_OUT_4[22]) );
  DLH_X1 \ADDR_OUT_4_reg[21]  ( .G(n13), .D(\CAM_MEM[3][21] ), .Q(
        ADDR_OUT_4[21]) );
  DLH_X1 \ADDR_OUT_4_reg[20]  ( .G(n13), .D(\CAM_MEM[3][20] ), .Q(
        ADDR_OUT_4[20]) );
  DLH_X1 \ADDR_OUT_4_reg[19]  ( .G(n13), .D(\CAM_MEM[3][19] ), .Q(
        ADDR_OUT_4[19]) );
  DLH_X1 \ADDR_OUT_4_reg[18]  ( .G(n13), .D(\CAM_MEM[3][18] ), .Q(
        ADDR_OUT_4[18]) );
  DLH_X1 \ADDR_OUT_4_reg[17]  ( .G(n13), .D(\CAM_MEM[3][17] ), .Q(
        ADDR_OUT_4[17]) );
  DLH_X1 \ADDR_OUT_4_reg[16]  ( .G(n13), .D(\CAM_MEM[3][16] ), .Q(
        ADDR_OUT_4[16]) );
  DLH_X1 \ADDR_OUT_4_reg[15]  ( .G(n13), .D(\CAM_MEM[3][15] ), .Q(
        ADDR_OUT_4[15]) );
  DLH_X1 \ADDR_OUT_4_reg[14]  ( .G(n13), .D(\CAM_MEM[3][14] ), .Q(
        ADDR_OUT_4[14]) );
  DLH_X1 \ADDR_OUT_4_reg[13]  ( .G(n13), .D(\CAM_MEM[3][13] ), .Q(
        ADDR_OUT_4[13]) );
  DLH_X1 \ADDR_OUT_4_reg[12]  ( .G(n13), .D(\CAM_MEM[3][12] ), .Q(
        ADDR_OUT_4[12]) );
  DLH_X1 \ADDR_OUT_4_reg[11]  ( .G(n13), .D(\CAM_MEM[3][11] ), .Q(
        ADDR_OUT_4[11]) );
  DLH_X1 \ADDR_OUT_4_reg[10]  ( .G(n1), .D(\CAM_MEM[3][10] ), .Q(
        ADDR_OUT_4[10]) );
  DLH_X1 \ADDR_OUT_4_reg[9]  ( .G(n1), .D(\CAM_MEM[3][9] ), .Q(ADDR_OUT_4[9])
         );
  DLH_X1 \ADDR_OUT_4_reg[8]  ( .G(n1), .D(\CAM_MEM[3][8] ), .Q(ADDR_OUT_4[8])
         );
  DLH_X1 \ADDR_OUT_4_reg[7]  ( .G(n1), .D(\CAM_MEM[3][7] ), .Q(ADDR_OUT_4[7])
         );
  DLH_X1 \ADDR_OUT_4_reg[6]  ( .G(n1), .D(\CAM_MEM[3][6] ), .Q(ADDR_OUT_4[6])
         );
  DLH_X1 \ADDR_OUT_4_reg[5]  ( .G(n1), .D(\CAM_MEM[3][5] ), .Q(ADDR_OUT_4[5])
         );
  DLH_X1 \ADDR_OUT_4_reg[4]  ( .G(n1), .D(\CAM_MEM[3][4] ), .Q(ADDR_OUT_4[4])
         );
  DLH_X1 \ADDR_OUT_4_reg[3]  ( .G(n1), .D(\CAM_MEM[3][3] ), .Q(ADDR_OUT_4[3])
         );
  DLH_X1 \ADDR_OUT_4_reg[2]  ( .G(n1), .D(\CAM_MEM[3][2] ), .Q(ADDR_OUT_4[2])
         );
  DLH_X1 \ADDR_OUT_4_reg[1]  ( .G(n1), .D(\CAM_MEM[3][1] ), .Q(ADDR_OUT_4[1])
         );
  DLH_X1 \ADDR_OUT_4_reg[0]  ( .G(n1), .D(\CAM_MEM[3][0] ), .Q(ADDR_OUT_4[0])
         );
  DLH_X1 VALID_1_reg ( .G(n1), .D(VALID_BIT[0]), .Q(VALID_1) );
  DLH_X1 VALID_2_reg ( .G(n1), .D(VALID_BIT[1]), .Q(VALID_2) );
  AND2_X1 U3 ( .A1(n2), .A2(n3), .ZN(N286) );
  NOR2_X1 U4 ( .A1(RST), .A2(WE), .ZN(N417) );
  AOI21_X1 U5 ( .B1(WE), .B2(n2), .A(RST), .ZN(n7) );
  AND2_X1 U6 ( .A1(WE), .A2(n23), .ZN(n3) );
  AND2_X1 U7 ( .A1(n6), .A2(n3), .ZN(N190) );
  AND2_X1 U8 ( .A1(n5), .A2(n3), .ZN(N222) );
  AND2_X1 U9 ( .A1(n4), .A2(n3), .ZN(N254) );
  INV_X1 U10 ( .A(RST), .ZN(n23) );
  NOR2_X1 U11 ( .A1(n8), .A2(n9), .ZN(n2) );
  AOI21_X1 U12 ( .B1(WE), .B2(n6), .A(RST), .ZN(n12) );
  AOI21_X1 U13 ( .B1(WE), .B2(n5), .A(RST), .ZN(n11) );
  AOI21_X1 U14 ( .B1(WE), .B2(n4), .A(RST), .ZN(n10) );
  NOR2_X1 U15 ( .A1(ADDR[0]), .A2(ADDR[1]), .ZN(n6) );
  NOR2_X1 U16 ( .A1(n8), .A2(ADDR[0]), .ZN(n4) );
  NOR2_X1 U17 ( .A1(n9), .A2(ADDR[1]), .ZN(n5) );
  INV_X1 U18 ( .A(ADDR[0]), .ZN(n9) );
  INV_X1 U19 ( .A(ADDR[1]), .ZN(n8) );
  CLKBUF_X1 U20 ( .A(N417), .Z(n1) );
  CLKBUF_X1 U21 ( .A(N417), .Z(n13) );
  CLKBUF_X1 U22 ( .A(N417), .Z(n14) );
  CLKBUF_X1 U23 ( .A(N417), .Z(n15) );
  CLKBUF_X1 U24 ( .A(N417), .Z(n16) );
  CLKBUF_X1 U25 ( .A(N417), .Z(n17) );
  CLKBUF_X1 U26 ( .A(N417), .Z(n18) );
  CLKBUF_X1 U27 ( .A(N417), .Z(n19) );
  CLKBUF_X1 U28 ( .A(N417), .Z(n20) );
  CLKBUF_X1 U29 ( .A(N417), .Z(n21) );
  CLKBUF_X1 U30 ( .A(N417), .Z(n22) );
endmodule


module NAND_GATE_0 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module INV_1_0 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module FA_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   OUT_XOR, n1;
  wire   [1:0] OUT_AND;

  XOR_GATE_1_637 XOR_GATE_1 ( .A(A), .B(B), .Y(OUT_XOR) );
  XOR_GATE_1_636 XOR_GATE_2 ( .A(n1), .B(Ci), .Y(S) );
  AND_GATE_1_702 AND_GATE_1 ( .A(A), .B(B), .Y(OUT_AND[0]) );
  AND_GATE_1_701 AND_GATE_2 ( .A(OUT_XOR), .B(Ci), .Y(OUT_AND[1]) );
  OR_GATE_338 OR_GATE_1 ( .A(OUT_AND[0]), .B(OUT_AND[1]), .Y(Co) );
  CLKBUF_X1 U1 ( .A(OUT_XOR), .Z(n1) );
endmodule


module HA_0 ( A, B, S, Co );
  input A, B;
  output S, Co;


  XOR_GATE_1_638 XOR_GATE_INST ( .A(A), .B(B), .Y(S) );
  AND_GATE_1_703 AND_GATE_INST ( .A(A), .B(B), .Y(Co) );
endmodule


module SYNC_COUNTER_5BIT ( EN, RST, CLK, COUNT );
  output [4:0] COUNT;
  input EN, RST, CLK;

  wire   [2:0] AND_SIG;

  FFT_0 FFT_1 ( .T(1'b1), .CLK(CLK), .EN(EN), .RST(RST), .Q(COUNT[0]) );
  FFT_6 FFT_2 ( .T(COUNT[0]), .CLK(CLK), .EN(EN), .RST(RST), .Q(COUNT[1]) );
  AND_GATE_1_706 AND_1 ( .A(COUNT[0]), .B(COUNT[1]), .Y(AND_SIG[0]) );
  FFT_5 FFT_3 ( .T(AND_SIG[0]), .CLK(CLK), .EN(EN), .RST(RST), .Q(COUNT[2]) );
  AND_GATE_1_705 AND_2 ( .A(AND_SIG[0]), .B(COUNT[2]), .Y(AND_SIG[1]) );
  FFT_4 FFT_4 ( .T(AND_SIG[1]), .CLK(CLK), .EN(EN), .RST(RST), .Q(COUNT[3]) );
  AND_GATE_1_704 AND_3 ( .A(AND_SIG[1]), .B(COUNT[3]), .Y(AND_SIG[2]) );
  FFT_3 FFT_5 ( .T(AND_SIG[2]), .CLK(CLK), .EN(EN), .RST(RST), .Q(COUNT[4]) );
endmodule


module EQU_COMPARATOR_N23 ( A, B, Y );
  input [22:0] A;
  input [22:0] B;
  output Y;

  wire   [22:0] L;

  XNOR_GATE_183 XNORING_0 ( .A(A[0]), .B(B[0]), .Y(L[0]) );
  XNOR_GATE_182 XNORING_1 ( .A(A[1]), .B(B[1]), .Y(L[1]) );
  XNOR_GATE_181 XNORING_2 ( .A(A[2]), .B(B[2]), .Y(L[2]) );
  XNOR_GATE_180 XNORING_3 ( .A(A[3]), .B(B[3]), .Y(L[3]) );
  XNOR_GATE_179 XNORING_4 ( .A(A[4]), .B(B[4]), .Y(L[4]) );
  XNOR_GATE_178 XNORING_5 ( .A(A[5]), .B(B[5]), .Y(L[5]) );
  XNOR_GATE_177 XNORING_6 ( .A(A[6]), .B(B[6]), .Y(L[6]) );
  XNOR_GATE_176 XNORING_7 ( .A(A[7]), .B(B[7]), .Y(L[7]) );
  XNOR_GATE_175 XNORING_8 ( .A(A[8]), .B(B[8]), .Y(L[8]) );
  XNOR_GATE_174 XNORING_9 ( .A(A[9]), .B(B[9]), .Y(L[9]) );
  XNOR_GATE_173 XNORING_10 ( .A(A[10]), .B(B[10]), .Y(L[10]) );
  XNOR_GATE_172 XNORING_11 ( .A(A[11]), .B(B[11]), .Y(L[11]) );
  XNOR_GATE_171 XNORING_12 ( .A(A[12]), .B(B[12]), .Y(L[12]) );
  XNOR_GATE_170 XNORING_13 ( .A(A[13]), .B(B[13]), .Y(L[13]) );
  XNOR_GATE_169 XNORING_14 ( .A(A[14]), .B(B[14]), .Y(L[14]) );
  XNOR_GATE_168 XNORING_15 ( .A(A[15]), .B(B[15]), .Y(L[15]) );
  XNOR_GATE_167 XNORING_16 ( .A(A[16]), .B(B[16]), .Y(L[16]) );
  XNOR_GATE_166 XNORING_17 ( .A(A[17]), .B(B[17]), .Y(L[17]) );
  XNOR_GATE_165 XNORING_18 ( .A(A[18]), .B(B[18]), .Y(L[18]) );
  XNOR_GATE_164 XNORING_19 ( .A(A[19]), .B(B[19]), .Y(L[19]) );
  XNOR_GATE_163 XNORING_20 ( .A(A[20]), .B(B[20]), .Y(L[20]) );
  XNOR_GATE_162 XNORING_21 ( .A(A[21]), .B(B[21]), .Y(L[21]) );
  XNOR_GATE_161 XNORING_22 ( .A(A[22]), .B(B[22]), .Y(L[22]) );
  N_AND_N23 ANDING ( .A(L), .Y(Y) );
endmodule


module CACHE_DATA_N32_N_DATA5_SET_BIT4 ( DATA_IN, DATA_OUT, ADDR, OFFSET, CLK, 
        WE );
  input [7:0] DATA_IN;
  output [31:0] DATA_OUT;
  input [3:0] ADDR;
  input [4:0] OFFSET;
  input CLK, WE;
  wire   N28803, N147559, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n77, n78, n79, n81, n82, n84, n85, n87, n88, n90, n91, n93, n94, n96,
         n97, n99, n100, n102, n103, n105, n106, n108, n109, n111, n112, n114,
         n115, n117, n118, n120, n121, n123, n124, n126, n127, n129, n130,
         n132, n133, n135, n136, n138, n139, n141, n142, n144, n145, n147,
         n148, n150, n151, n153, n154, n156, n157, n159, n160, n162, n163,
         n165, n166, n168, n169, n171, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1183, n1186, n1187, n1188,
         n1189, n1192, n1195, n1196, n1197, n1198, n1201, n1204, n1205, n1206,
         n1207, n1210, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1223, n1226, n1227, n1228, n1229, n1232, n1235, n1236, n1237, n1238,
         n1241, n1244, n1245, n1246, n1247, n1250, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1263, n1266, n1267, n1268, n1269, n1272,
         n1275, n1276, n1277, n1278, n1281, n1284, n1285, n1286, n1287, n1290,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1303, n1306,
         n1307, n1308, n1309, n1312, n1315, n1316, n1317, n1318, n1321, n1324,
         n1325, n1326, n1327, n1330, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1347, n1350, n1351, n1352,
         n1355, n1358, n1359, n1360, n1363, n1366, n1367, n1368, n1371, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1383, n1386, n1387, n1388,
         n1391, n1394, n1395, n1396, n1399, n1402, n1403, n1404, n1407, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1419, n1422, n1423, n1424,
         n1427, n1430, n1431, n1432, n1435, n1438, n1439, n1440, n1443, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1455, n1458, n1459, n1460,
         n1463, n1466, n1467, n1468, n1471, n1474, n1475, n1476, n1479, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1496, n1499, n1500, n1501, n1504, n1507, n1508, n1509, n1512,
         n1515, n1516, n1517, n1520, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1532, n1535, n1536, n1537, n1540, n1543, n1544, n1545, n1548,
         n1551, n1552, n1553, n1556, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1568, n1571, n1572, n1573, n1576, n1579, n1580, n1581, n1584,
         n1587, n1588, n1589, n1592, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1604, n1607, n1608, n1609, n1612, n1615, n1616, n1617, n1620,
         n1623, n1624, n1625, n1628, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1645, n1648, n1649, n1650,
         n1653, n1656, n1657, n1658, n1661, n1664, n1665, n1666, n1669, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1681, n1684, n1685, n1686,
         n1689, n1692, n1693, n1694, n1697, n1700, n1701, n1702, n1705, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1717, n1720, n1721, n1722,
         n1725, n1728, n1729, n1730, n1733, n1736, n1737, n1738, n1741, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1753, n1756, n1757, n1758,
         n1761, n1764, n1765, n1766, n1769, n1772, n1773, n1774, n1777, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1794, n1797, n1798, n1799, n1802, n1805, n1806, n1807, n1810,
         n1813, n1814, n1815, n1818, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1830, n1833, n1834, n1835, n1838, n1841, n1842, n1843, n1846,
         n1849, n1850, n1851, n1854, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1866, n1869, n1870, n1871, n1874, n1877, n1878, n1879, n1882,
         n1885, n1886, n1887, n1890, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1902, n1905, n1906, n1907, n1910, n1913, n1914, n1915, n1918,
         n1921, n1922, n1923, n1926, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1943, n1946, n1947, n1948,
         n1951, n1954, n1955, n1956, n1959, n1962, n1963, n1964, n1967, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1979, n1982, n1983, n1984,
         n1987, n1990, n1991, n1992, n1995, n1998, n1999, n2000, n2003, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2015, n2018, n2019, n2020,
         n2023, n2026, n2027, n2028, n2031, n2034, n2035, n2036, n2039, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2051, n2054, n2055, n2056,
         n2059, n2062, n2063, n2064, n2067, n2070, n2071, n2072, n2075, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2092, n2095, n2096, n2097, n2100, n2103, n2104, n2105, n2108,
         n2111, n2112, n2113, n2116, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2128, n2131, n2132, n2133, n2136, n2139, n2140, n2141, n2144,
         n2147, n2148, n2149, n2152, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2164, n2167, n2168, n2169, n2172, n2175, n2176, n2177, n2180,
         n2183, n2184, n2185, n2188, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2200, n2203, n2204, n2205, n2208, n2211, n2212, n2213, n2216,
         n2219, n2220, n2221, n2224, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2241, n2244, n2245, n2246,
         n2249, n2252, n2253, n2254, n2257, n2260, n2261, n2262, n2265, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2277, n2280, n2281, n2282,
         n2285, n2288, n2289, n2290, n2293, n2296, n2297, n2298, n2301, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2313, n2316, n2317, n2318,
         n2321, n2324, n2325, n2326, n2329, n2332, n2333, n2334, n2337, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2349, n2352, n2353, n2354,
         n2357, n2360, n2361, n2362, n2365, n2368, n2369, n2370, n2373, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2390, n2393, n2394, n2395, n2398, n2401, n2402, n2403, n2406,
         n2409, n2410, n2411, n2414, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2426, n2429, n2430, n2431, n2434, n2437, n2438, n2439, n2442,
         n2445, n2446, n2447, n2450, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2462, n2465, n2466, n2467, n2470, n2473, n2474, n2475, n2478,
         n2481, n2482, n2483, n2486, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2498, n2501, n2502, n2503, n2506, n2509, n2510, n2511, n2514,
         n2517, n2518, n2519, n2522, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2539, n2542, n2543, n2544,
         n2547, n2550, n2551, n2552, n2555, n2558, n2559, n2560, n2563, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2575, n2578, n2579, n2580,
         n2583, n2586, n2587, n2588, n2591, n2594, n2595, n2596, n2599, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2611, n2614, n2615, n2616,
         n2619, n2622, n2623, n2624, n2627, n2630, n2631, n2632, n2635, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2647, n2650, n2651, n2652,
         n2655, n2658, n2659, n2660, n2663, n2666, n2667, n2668, n2671, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2688, n2691, n2692, n2693, n2696, n2699, n2700, n2701, n2704,
         n2707, n2708, n2709, n2712, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2724, n2727, n2728, n2729, n2732, n2735, n2736, n2737, n2740,
         n2743, n2744, n2745, n2748, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2760, n2763, n2764, n2765, n2768, n2771, n2772, n2773, n2776,
         n2779, n2780, n2781, n2784, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2796, n2799, n2800, n2801, n2804, n2807, n2808, n2809, n2812,
         n2815, n2816, n2817, n2820, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2837, n2840, n2841, n2842,
         n2845, n2848, n2849, n2850, n2853, n2856, n2857, n2858, n2861, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2873, n2876, n2877, n2878,
         n2881, n2884, n2885, n2886, n2889, n2892, n2893, n2894, n2897, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2909, n2912, n2913, n2914,
         n2917, n2920, n2921, n2922, n2925, n2928, n2929, n2930, n2933, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2945, n2948, n2949, n2950,
         n2953, n2956, n2957, n2958, n2961, n2964, n2965, n2966, n2969, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2986, n2989, n2990, n2991, n2994, n2997, n2998, n2999, n3002,
         n3005, n3006, n3007, n3010, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3022, n3025, n3026, n3027, n3030, n3033, n3034, n3035, n3038,
         n3041, n3042, n3043, n3046, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3058, n3061, n3062, n3063, n3066, n3069, n3070, n3071, n3074,
         n3077, n3078, n3079, n3082, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3094, n3097, n3098, n3099, n3102, n3105, n3106, n3107, n3110,
         n3113, n3114, n3115, n3118, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3135, n3138, n3139, n3140,
         n3143, n3146, n3147, n3148, n3151, n3154, n3155, n3156, n3159, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3171, n3174, n3175, n3176,
         n3179, n3182, n3183, n3184, n3187, n3190, n3191, n3192, n3195, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3207, n3210, n3211, n3212,
         n3215, n3218, n3219, n3220, n3223, n3226, n3227, n3228, n3231, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3243, n3246, n3247, n3248,
         n3251, n3254, n3255, n3256, n3259, n3262, n3263, n3264, n3267, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3284, n3287, n3288, n3289, n3292, n3295, n3296, n3297, n3300,
         n3303, n3304, n3305, n3308, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3320, n3323, n3324, n3325, n3328, n3331, n3332, n3333, n3336,
         n3339, n3340, n3341, n3344, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3356, n3359, n3360, n3361, n3364, n3367, n3368, n3369, n3372,
         n3375, n3376, n3377, n3380, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3392, n3395, n3396, n3397, n3400, n3403, n3404, n3405, n3408,
         n3411, n3412, n3413, n3416, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3433, n3436, n3437, n3438,
         n3441, n3444, n3445, n3446, n3449, n3452, n3453, n3454, n3457, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3469, n3472, n3473, n3474,
         n3477, n3480, n3481, n3482, n3485, n3488, n3489, n3490, n3493, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3505, n3508, n3509, n3510,
         n3513, n3516, n3517, n3518, n3521, n3524, n3525, n3526, n3529, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3541, n3544, n3545, n3546,
         n3549, n3552, n3553, n3554, n3557, n3560, n3561, n3562, n3565, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3582, n3585, n3586, n3587, n3590, n3593, n3594, n3595, n3598,
         n3601, n3602, n3603, n3606, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3618, n3621, n3622, n3623, n3626, n3629, n3630, n3631, n3634,
         n3637, n3638, n3639, n3642, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3654, n3657, n3658, n3659, n3662, n3665, n3666, n3667, n3670,
         n3673, n3674, n3675, n3678, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3690, n3693, n3694, n3695, n3698, n3701, n3702, n3703, n3706,
         n3709, n3710, n3711, n3714, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3731, n3734, n3735, n3736,
         n3739, n3742, n3743, n3744, n3747, n3750, n3751, n3752, n3755, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3767, n3770, n3771, n3772,
         n3775, n3778, n3779, n3780, n3783, n3786, n3787, n3788, n3791, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3803, n3806, n3807, n3808,
         n3811, n3814, n3815, n3816, n3819, n3822, n3823, n3824, n3827, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3839, n3842, n3843, n3844,
         n3847, n3850, n3851, n3852, n3855, n3858, n3859, n3860, n3863, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3880, n3883, n3884, n3885, n3888, n3891, n3892, n3893, n3896,
         n3899, n3900, n3901, n3904, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3916, n3919, n3920, n3921, n3924, n3927, n3928, n3929, n3932,
         n3935, n3936, n3937, n3940, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3952, n3955, n3956, n3957, n3960, n3963, n3964, n3965, n3968,
         n3971, n3972, n3973, n3976, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3988, n3991, n3992, n3993, n3996, n3999, n4000, n4001, n4004,
         n4007, n4008, n4009, n4012, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4029, n4032, n4033, n4034,
         n4037, n4040, n4041, n4042, n4045, n4048, n4049, n4050, n4053, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4065, n4068, n4069, n4070,
         n4073, n4076, n4077, n4078, n4081, n4084, n4085, n4086, n4089, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4101, n4104, n4105, n4106,
         n4109, n4112, n4113, n4114, n4117, n4120, n4121, n4122, n4125, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4137, n4140, n4141, n4142,
         n4145, n4148, n4149, n4150, n4153, n4156, n4157, n4158, n4161, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4178, n4181, n4182, n4183, n4186, n4189, n4190, n4191, n4194,
         n4197, n4198, n4199, n4202, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4214, n4217, n4218, n4219, n4222, n4225, n4226, n4227, n4230,
         n4233, n4234, n4235, n4238, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4250, n4253, n4254, n4255, n4258, n4261, n4262, n4263, n4266,
         n4269, n4270, n4271, n4274, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4286, n4289, n4290, n4291, n4294, n4297, n4298, n4299, n4302,
         n4305, n4306, n4307, n4310, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4327, n4330, n4331, n4332,
         n4335, n4338, n4339, n4340, n4343, n4346, n4347, n4348, n4351, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4363, n4366, n4367, n4368,
         n4371, n4374, n4375, n4376, n4379, n4382, n4383, n4384, n4387, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4399, n4402, n4403, n4404,
         n4407, n4410, n4411, n4412, n4415, n4418, n4419, n4420, n4423, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4435, n4438, n4439, n4440,
         n4443, n4446, n4447, n4448, n4451, n4454, n4455, n4456, n4459, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4476, n4479, n4480, n4481, n4484, n4487, n4488, n4489, n4492,
         n4495, n4496, n4497, n4500, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4512, n4515, n4516, n4517, n4520, n4523, n4524, n4525, n4528,
         n4531, n4532, n4533, n4536, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4548, n4551, n4552, n4553, n4556, n4559, n4560, n4561, n4564,
         n4567, n4568, n4569, n4572, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4584, n4587, n4588, n4589, n4592, n4595, n4596, n4597, n4600,
         n4603, n4604, n4605, n4608, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4625, n4628, n4629, n4630,
         n4633, n4636, n4637, n4638, n4641, n4644, n4645, n4646, n4649, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4661, n4664, n4665, n4666,
         n4669, n4672, n4673, n4674, n4677, n4680, n4681, n4682, n4685, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4697, n4700, n4701, n4702,
         n4705, n4708, n4709, n4710, n4713, n4716, n4717, n4718, n4721, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4733, n4736, n4737, n4738,
         n4741, n4744, n4745, n4746, n4749, n4752, n4753, n4754, n4757, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4774, n4777, n4778, n4779, n4782, n4785, n4786, n4787, n4790,
         n4793, n4794, n4795, n4798, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4810, n4813, n4814, n4815, n4818, n4821, n4822, n4823, n4826,
         n4829, n4830, n4831, n4834, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4846, n4849, n4850, n4851, n4854, n4857, n4858, n4859, n4862,
         n4865, n4866, n4867, n4870, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4882, n4885, n4886, n4887, n4890, n4893, n4894, n4895, n4898,
         n4901, n4902, n4903, n4906, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4923, n4926, n4927, n4928,
         n4931, n4934, n4935, n4936, n4939, n4942, n4943, n4944, n4947, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4959, n4962, n4963, n4964,
         n4967, n4970, n4971, n4972, n4975, n4978, n4979, n4980, n4983, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4995, n4998, n4999, n5000,
         n5003, n5006, n5007, n5008, n5011, n5014, n5015, n5016, n5019, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5031, n5034, n5035, n5036,
         n5039, n5042, n5043, n5044, n5047, n5050, n5051, n5052, n5055, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5072, n5075, n5076, n5077, n5080, n5083, n5084, n5085, n5088,
         n5091, n5092, n5093, n5096, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5108, n5111, n5112, n5113, n5116, n5119, n5120, n5121, n5124,
         n5127, n5128, n5129, n5132, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5144, n5147, n5148, n5149, n5152, n5155, n5156, n5157, n5160,
         n5163, n5164, n5165, n5168, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5180, n5183, n5184, n5185, n5188, n5191, n5192, n5193, n5196,
         n5199, n5200, n5201, n5204, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5221, n5224, n5225, n5226,
         n5229, n5232, n5233, n5234, n5237, n5240, n5241, n5242, n5245, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5257, n5260, n5261, n5262,
         n5265, n5268, n5269, n5270, n5273, n5276, n5277, n5278, n5281, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5293, n5296, n5297, n5298,
         n5301, n5304, n5305, n5306, n5309, n5312, n5313, n5314, n5317, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5329, n5332, n5333, n5334,
         n5337, n5340, n5341, n5342, n5345, n5348, n5349, n5350, n5353, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5370, n5373, n5374, n5375, n5378, n5381, n5382, n5383, n5386,
         n5389, n5390, n5391, n5394, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5406, n5409, n5410, n5411, n5414, n5417, n5418, n5419, n5422,
         n5425, n5426, n5427, n5430, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5442, n5445, n5446, n5447, n5450, n5453, n5454, n5455, n5458,
         n5461, n5462, n5463, n5466, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5478, n5481, n5482, n5483, n5486, n5489, n5490, n5491, n5494,
         n5497, n5498, n5499, n5502, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5519, n5522, n5523, n5524,
         n5527, n5530, n5531, n5532, n5535, n5538, n5539, n5540, n5543, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5555, n5558, n5559, n5560,
         n5563, n5566, n5567, n5568, n5571, n5574, n5575, n5576, n5579, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5591, n5594, n5595, n5596,
         n5599, n5602, n5603, n5604, n5607, n5610, n5611, n5612, n5615, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5627, n5630, n5631, n5632,
         n5635, n5638, n5639, n5640, n5643, n5646, n5647, n5648, n5651, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5668, n5671, n5672, n5673, n5676, n5679, n5680, n5681, n5684,
         n5687, n5688, n5689, n5692, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5704, n5707, n5708, n5709, n5712, n5715, n5716, n5717, n5720,
         n5723, n5724, n5725, n5728, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5740, n5743, n5744, n5745, n5748, n5751, n5752, n5753, n5756,
         n5759, n5760, n5761, n5764, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5776, n5779, n5780, n5781, n5784, n5787, n5788, n5789, n5792,
         n5795, n5796, n5797, n5800, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5817, n5820, n5821, n5822,
         n5825, n5828, n5829, n5830, n5833, n5836, n5837, n5838, n5841, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5853, n5856, n5857, n5858,
         n5861, n5864, n5865, n5866, n5869, n5872, n5873, n5874, n5877, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5891, n5894,
         n5895, n5896, n5899, n5902, n5903, n5904, n5907, n5910, n5911, n5912,
         n5915, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5927, n5930,
         n5931, n5932, n5935, n5938, n5939, n5940, n5943, n5946, n5947, n5948,
         n5951, n5952, n5953, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n76, n80, n83, n86, n89, n92, n95, n98, n101, n104, n107, n110, n113,
         n116, n119, n122, n125, n128, n131, n134, n137, n140, n143, n146,
         n149, n152, n155, n158, n161, n164, n167, n170, n172, n238, n1181,
         n1182, n1184, n1185, n1190, n1191, n1193, n1194, n1199, n1200, n1202,
         n1203, n1208, n1209, n1211, n1212, n1221, n1222, n1224, n1225, n1230,
         n1231, n1233, n1234, n1239, n1240, n1242, n1243, n1248, n1249, n1251,
         n1252, n1261, n1262, n1264, n1265, n1270, n1271, n1273, n1274, n1279,
         n1280, n1282, n1283, n1288, n1289, n1291, n1292, n1301, n1302, n1304,
         n1305, n1310, n1311, n1313, n1314, n1319, n1320, n1322, n1323, n1328,
         n1329, n1331, n1332, n1345, n1346, n1348, n1349, n1353, n1354, n1356,
         n1357, n1361, n1362, n1364, n1365, n1369, n1370, n1372, n1373, n1381,
         n1382, n1384, n1385, n1389, n1390, n1392, n1393, n1397, n1398, n1400,
         n1401, n1405, n1406, n1408, n1409, n1417, n1418, n1420, n1421, n1425,
         n1426, n1428, n1429, n1433, n1434, n1436, n1437, n1441, n1442, n1444,
         n1445, n1453, n1454, n1456, n1457, n1461, n1462, n1464, n1465, n1469,
         n1470, n1472, n1473, n1477, n1478, n1480, n1481, n1494, n1495, n1497,
         n1498, n1502, n1503, n1505, n1506, n1510, n1511, n1513, n1514, n1518,
         n1519, n1521, n1522, n1530, n1531, n1533, n1534, n1538, n1539, n1541,
         n1542, n1546, n1547, n1549, n1550, n1554, n1555, n1557, n1558, n1566,
         n1567, n1569, n1570, n1574, n1575, n1577, n1578, n1582, n1583, n1585,
         n1586, n1590, n1591, n1593, n1594, n1602, n1603, n1605, n1606, n1610,
         n1611, n1613, n1614, n1618, n1619, n1621, n1622, n1626, n1627, n1629,
         n1630, n1643, n1644, n1646, n1647, n1651, n1652, n1654, n1655, n1659,
         n1660, n1662, n1663, n1667, n1668, n1670, n1671, n1679, n1680, n1682,
         n1683, n1687, n1688, n1690, n1691, n1695, n1696, n1698, n1699, n1703,
         n1704, n1706, n1707, n1715, n1716, n1718, n1719, n1723, n1724, n1726,
         n1727, n1731, n1732, n1734, n1735, n1739, n1740, n1742, n1743, n1751,
         n1752, n1754, n1755, n1759, n1760, n1762, n1763, n1767, n1768, n1770,
         n1771, n1775, n1776, n1778, n1779, n1792, n1793, n1795, n1796, n1800,
         n1801, n1803, n1804, n1808, n1809, n1811, n1812, n1816, n1817, n1819,
         n1820, n1828, n1829, n1831, n1832, n1836, n1837, n1839, n1840, n1844,
         n1845, n1847, n1848, n1852, n1853, n1855, n1856, n1864, n1865, n1867,
         n1868, n1872, n1873, n1875, n1876, n1880, n1881, n1883, n1884, n1888,
         n1889, n1891, n1892, n1900, n1901, n1903, n1904, n1908, n1909, n1911,
         n1912, n1916, n1917, n1919, n1920, n1924, n1925, n1927, n1928, n1941,
         n1942, n1944, n1945, n1949, n1950, n1952, n1953, n1957, n1958, n1960,
         n1961, n1965, n1966, n1968, n1969, n1977, n1978, n1980, n1981, n1985,
         n1986, n1988, n1989, n1993, n1994, n1996, n1997, n2001, n2002, n2004,
         n2005, n2013, n2014, n2016, n2017, n2021, n2022, n2024, n2025, n2029,
         n2030, n2032, n2033, n2037, n2038, n2040, n2041, n2049, n2050, n2052,
         n2053, n2057, n2058, n2060, n2061, n2065, n2066, n2068, n2069, n2073,
         n2074, n2076, n2077, n2090, n2091, n2093, n2094, n2098, n2099, n2101,
         n2102, n2106, n2107, n2109, n2110, n2114, n2115, n2117, n2118, n2126,
         n2127, n2129, n2130, n2134, n2135, n2137, n2138, n2142, n2143, n2145,
         n2146, n2150, n2151, n2153, n2154, n2162, n2163, n2165, n2166, n2170,
         n2171, n2173, n2174, n2178, n2179, n2181, n2182, n2186, n2187, n2189,
         n2190, n2198, n2199, n2201, n2202, n2206, n2207, n2209, n2210, n2214,
         n2215, n2217, n2218, n2222, n2223, n2225, n2226, n2239, n2240, n2242,
         n2243, n2247, n2248, n2250, n2251, n2255, n2256, n2258, n2259, n2263,
         n2264, n2266, n2267, n2275, n2276, n2278, n2279, n2283, n2284, n2286,
         n2287, n2291, n2292, n2294, n2295, n2299, n2300, n2302, n2303, n2311,
         n2312, n2314, n2315, n2319, n2320, n2322, n2323, n2327, n2328, n2330,
         n2331, n2335, n2336, n2338, n2339, n2347, n2348, n2350, n2351, n2355,
         n2356, n2358, n2359, n2363, n2364, n2366, n2367, n2371, n2372, n2374,
         n2375, n2388, n2389, n2391, n2392, n2396, n2397, n2399, n2400, n2404,
         n2405, n2407, n2408, n2412, n2413, n2415, n2416, n2424, n2425, n2427,
         n2428, n2432, n2433, n2435, n2436, n2440, n2441, n2443, n2444, n2448,
         n2449, n2451, n2452, n2460, n2461, n2463, n2464, n2468, n2469, n2471,
         n2472, n2476, n2477, n2479, n2480, n2484, n2485, n2487, n2488, n2496,
         n2497, n2499, n2500, n2504, n2505, n2507, n2508, n2512, n2513, n2515,
         n2516, n2520, n2521, n2523, n2524, n2537, n2538, n2540, n2541, n2545,
         n2546, n2548, n2549, n2553, n2554, n2556, n2557, n2561, n2562, n2564,
         n2565, n2573, n2574, n2576, n2577, n2581, n2582, n2584, n2585, n2589,
         n2590, n2592, n2593, n2597, n2598, n2600, n2601, n2609, n2610, n2612,
         n2613, n2617, n2618, n2620, n2621, n2625, n2626, n2628, n2629, n2633,
         n2634, n2636, n2637, n2645, n2646, n2648, n2649, n2653, n2654, n2656,
         n2657, n2661, n2662, n2664, n2665, n2669, n2670, n2672, n2673, n2686,
         n2687, n2689, n2690, n2694, n2695, n2697, n2698, n2702, n2703, n2705,
         n2706, n2710, n2711, n2713, n2714, n2722, n2723, n2725, n2726, n2730,
         n2731, n2733, n2734, n2738, n2739, n2741, n2742, n2746, n2747, n2749,
         n2750, n2758, n2759, n2761, n2762, n2766, n2767, n2769, n2770, n2774,
         n2775, n2777, n2778, n2782, n2783, n2785, n2786, n2794, n2795, n2797,
         n2798, n2802, n2803, n2805, n2806, n2810, n2811, n2813, n2814, n2818,
         n2819, n2821, n2822, n2835, n2836, n2838, n2839, n2843, n2844, n2846,
         n2847, n2851, n2852, n2854, n2855, n2859, n2860, n2862, n2863, n2871,
         n2872, n2874, n2875, n2879, n2880, n2882, n2883, n2887, n2888, n2890,
         n2891, n2895, n2896, n2898, n2899, n2907, n2908, n2910, n2911, n2915,
         n2916, n2918, n2919, n2923, n2924, n2926, n2927, n2931, n2932, n2934,
         n2935, n2943, n2944, n2946, n2947, n2951, n2952, n2954, n2955, n2959,
         n2960, n2962, n2963, n2967, n2968, n2970, n2971, n2984, n2985, n2987,
         n2988, n2992, n2993, n2995, n2996, n3000, n3001, n3003, n3004, n3008,
         n3009, n3011, n3012, n3020, n3021, n3023, n3024, n3028, n3029, n3031,
         n3032, n3036, n3037, n3039, n3040, n3044, n3045, n3047, n3048, n3056,
         n3057, n3059, n3060, n3064, n3065, n3067, n3068, n3072, n3073, n3075,
         n3076, n3080, n3081, n3083, n3084, n3092, n3093, n3095, n3096, n3100,
         n3101, n3103, n3104, n3108, n3109, n3111, n3112, n3116, n3117, n3119,
         n3120, n3133, n3134, n3136, n3137, n3141, n3142, n3144, n3145, n3149,
         n3150, n3152, n3153, n3157, n3158, n3160, n3161, n3169, n3170, n3172,
         n3173, n3177, n3178, n3180, n3181, n3185, n3186, n3188, n3189, n3193,
         n3194, n3196, n3197, n3205, n3206, n3208, n3209, n3213, n3214, n3216,
         n3217, n3221, n3222, n3224, n3225, n3229, n3230, n3232, n3233, n3241,
         n3242, n3244, n3245, n3249, n3250, n3252, n3253, n3257, n3258, n3260,
         n3261, n3265, n3266, n3268, n3269, n3282, n3283, n3285, n3286, n3290,
         n3291, n3293, n3294, n3298, n3299, n3301, n3302, n3306, n3307, n3309,
         n3310, n3318, n3319, n3321, n3322, n3326, n3327, n3329, n3330, n3334,
         n3335, n3337, n3338, n3342, n3343, n3345, n3346, n3354, n3355, n3357,
         n3358, n3362, n3363, n3365, n3366, n3370, n3371, n3373, n3374, n3378,
         n3379, n3381, n3382, n3390, n3391, n3393, n3394, n3398, n3399, n3401,
         n3402, n3406, n3407, n3409, n3410, n3414, n3415, n3417, n3418, n3431,
         n3432, n3434, n3435, n3439, n3440, n3442, n3443, n3447, n3448, n3450,
         n3451, n3455, n3456, n3458, n3459, n3467, n3468, n3470, n3471, n3475,
         n3476, n3478, n3479, n3483, n3484, n3486, n3487, n3491, n3492, n3494,
         n3495, n3503, n3504, n3506, n3507, n3511, n3512, n3514, n3515, n3519,
         n3520, n3522, n3523, n3527, n3528, n3530, n3531, n3539, n3540, n3542,
         n3543, n3547, n3548, n3550, n3551, n3555, n3556, n3558, n3559, n3563,
         n3564, n3566, n3567, n3580, n3581, n3583, n3584, n3588, n3589, n3591,
         n3592, n3596, n3597, n3599, n3600, n3604, n3605, n3607, n3608, n3616,
         n3617, n3619, n3620, n3624, n3625, n3627, n3628, n3632, n3633, n3635,
         n3636, n3640, n3641, n3643, n3644, n3652, n3653, n3655, n3656, n3660,
         n3661, n3663, n3664, n3668, n3669, n3671, n3672, n3676, n3677, n3679,
         n3680, n3688, n3689, n3691, n3692, n3696, n3697, n3699, n3700, n3704,
         n3705, n3707, n3708, n3712, n3713, n3715, n3716, n3729, n3730, n3732,
         n3733, n3737, n3738, n3740, n3741, n3745, n3746, n3748, n3749, n3753,
         n3754, n3756, n3757, n3765, n3766, n3768, n3769, n3773, n3774, n3776,
         n3777, n3781, n3782, n3784, n3785, n3789, n3790, n3792, n3793, n3801,
         n3802, n3804, n3805, n3809, n3810, n3812, n3813, n3817, n3818, n3820,
         n3821, n3825, n3826, n3828, n3829, n3837, n3838, n3840, n3841, n3845,
         n3846, n3848, n3849, n3853, n3854, n3856, n3857, n3861, n3862, n3864,
         n3865, n3878, n3879, n3881, n3882, n3886, n3887, n3889, n3890, n3894,
         n3895, n3897, n3898, n3902, n3903, n3905, n3906, n3914, n3915, n3917,
         n3918, n3922, n3923, n3925, n3926, n3930, n3931, n3933, n3934, n3938,
         n3939, n3941, n3942, n3950, n3951, n3953, n3954, n3958, n3959, n3961,
         n3962, n3966, n3967, n3969, n3970, n3974, n3975, n3977, n3978, n3986,
         n3987, n3989, n3990, n3994, n3995, n3997, n3998, n4002, n4003, n4005,
         n4006, n4010, n4011, n4013, n4014, n4027, n4028, n4030, n4031, n4035,
         n4036, n4038, n4039, n4043, n4044, n4046, n4047, n4051, n4052, n4054,
         n4055, n4063, n4064, n4066, n4067, n4071, n4072, n4074, n4075, n4079,
         n4080, n4082, n4083, n4087, n4088, n4090, n4091, n4099, n4100, n4102,
         n4103, n4107, n4108, n4110, n4111, n4115, n4116, n4118, n4119, n4123,
         n4124, n4126, n4127, n4135, n4136, n4138, n4139, n4143, n4144, n4146,
         n4147, n4151, n4152, n4154, n4155, n4159, n4160, n4162, n4163, n4176,
         n4177, n4179, n4180, n4184, n4185, n4187, n4188, n4192, n4193, n4195,
         n4196, n4200, n4201, n4203, n4204, n4212, n4213, n4215, n4216, n4220,
         n4221, n4223, n4224, n4228, n4229, n4231, n4232, n4236, n4237, n4239,
         n4240, n4248, n4249, n4251, n4252, n4256, n4257, n4259, n4260, n4264,
         n4265, n4267, n4268, n4272, n4273, n4275, n4276, n4284, n4285, n4287,
         n4288, n4292, n4293, n4295, n4296, n4300, n4301, n4303, n4304, n4308,
         n4309, n4311, n4312, n4325, n4326, n4328, n4329, n4333, n4334, n4336,
         n4337, n4341, n4342, n4344, n4345, n4349, n4350, n4352, n4353, n4361,
         n4362, n4364, n4365, n4369, n4370, n4372, n4373, n4377, n4378, n4380,
         n4381, n4385, n4386, n4388, n4389, n4397, n4398, n4400, n4401, n4405,
         n4406, n4408, n4409, n4413, n4414, n4416, n4417, n4421, n4422, n4424,
         n4425, n4433, n4434, n4436, n4437, n4441, n4442, n4444, n4445, n4449,
         n4450, n4452, n4453, n4457, n4458, n4460, n4461, n4474, n4475, n4477,
         n4478, n4482, n4483, n4485, n4486, n4490, n4491, n4493, n4494, n4498,
         n4499, n4501, n4502, n4510, n4511, n4513, n4514, n4518, n4519, n4521,
         n4522, n4526, n4527, n4529, n4530, n4534, n4535, n4537, n4538, n4546,
         n4547, n4549, n4550, n4554, n4555, n4557, n4558, n4562, n4563, n4565,
         n4566, n4570, n4571, n4573, n4574, n4582, n4583, n4585, n4586, n4590,
         n4591, n4593, n4594, n4598, n4599, n4601, n4602, n4606, n4607, n4609,
         n4610, n4623, n4624, n4626, n4627, n4631, n4632, n4634, n4635, n4639,
         n4640, n4642, n4643, n4647, n4648, n4650, n4651, n4659, n4660, n4662,
         n4663, n4667, n4668, n4670, n4671, n4675, n4676, n4678, n4679, n4683,
         n4684, n4686, n4687, n4695, n4696, n4698, n4699, n4703, n4704, n4706,
         n4707, n4711, n4712, n4714, n4715, n4719, n4720, n4722, n4723, n4731,
         n4732, n4734, n4735, n4739, n4740, n4742, n4743, n4747, n4748, n4750,
         n4751, n4755, n4756, n4758, n4759, n4772, n4773, n4775, n4776, n4780,
         n4781, n4783, n4784, n4788, n4789, n4791, n4792, n4796, n4797, n4799,
         n4800, n4808, n4809, n4811, n4812, n4816, n4817, n4819, n4820, n4824,
         n4825, n4827, n4828, n4832, n4833, n4835, n4836, n4844, n4845, n4847,
         n4848, n4852, n4853, n4855, n4856, n4860, n4861, n4863, n4864, n4868,
         n4869, n4871, n4872, n4880, n4881, n4883, n4884, n4888, n4889, n4891,
         n4892, n4896, n4897, n4899, n4900, n4904, n4905, n4907, n4908, n4921,
         n4922, n4924, n4925, n4929, n4930, n4932, n4933, n4937, n4938, n4940,
         n4941, n4945, n4946, n4948, n4949, n4957, n4958, n4960, n4961, n4965,
         n4966, n4968, n4969, n4973, n4974, n4976, n4977, n4981, n4982, n4984,
         n4985, n4993, n4994, n4996, n4997, n5001, n5002, n5004, n5005, n5009,
         n5010, n5012, n5013, n5017, n5018, n5020, n5021, n5029, n5030, n5032,
         n5033, n5037, n5038, n5040, n5041, n5045, n5046, n5048, n5049, n5053,
         n5054, n5056, n5057, n5070, n5071, n5073, n5074, n5078, n5079, n5081,
         n5082, n5086, n5087, n5089, n5090, n5094, n5095, n5097, n5098, n5106,
         n5107, n5109, n5110, n5114, n5115, n5117, n5118, n5122, n5123, n5125,
         n5126, n5130, n5131, n5133, n5134, n5142, n5143, n5145, n5146, n5150,
         n5151, n5153, n5154, n5158, n5159, n5161, n5162, n5166, n5167, n5169,
         n5170, n5178, n5179, n5181, n5182, n5186, n5187, n5189, n5190, n5194,
         n5195, n5197, n5198, n5202, n5203, n5205, n5206, n5219, n5220, n5222,
         n5223, n5227, n5228, n5230, n5231, n5235, n5236, n5238, n5239, n5243,
         n5244, n5246, n5247, n5255, n5256, n5258, n5259, n5263, n5264, n5266,
         n5267, n5271, n5272, n5274, n5275, n5279, n5280, n5282, n5283, n5291,
         n5292, n5294, n5295, n5299, n5300, n5302, n5303, n5307, n5308, n5310,
         n5311, n5315, n5316, n5318, n5319, n5327, n5328, n5330, n5331, n5335,
         n5336, n5338, n5339, n5343, n5344, n5346, n5347, n5351, n5352, n5354,
         n5355, n5368, n5369, n5371, n5372, n5376, n5377, n5379, n5380, n5384,
         n5385, n5387, n5388, n5392, n5393, n5395, n5396, n5404, n5405, n5407,
         n5408, n5412, n5413, n5415, n5416, n5420, n5421, n5423, n5424, n5428,
         n5429, n5431, n5432, n5440, n5441, n5443, n5444, n5448, n5449, n5451,
         n5452, n5456, n5457, n5459, n5460, n5464, n5465, n5467, n5468, n5476,
         n5477, n5479, n5480, n5484, n5485, n5487, n5488, n5492, n5493, n5495,
         n5496, n5500, n5501, n5503, n5504, n5517, n5518, n5520, n5521, n5525,
         n5526, n5528, n5529, n5533, n5534, n5536, n5537, n5541, n5542, n5544,
         n5545, n5553, n5554, n5556, n5557, n5561, n5562, n5564, n5565, n5569,
         n5570, n5572, n5573, n5577, n5578, n5580, n5581, n5589, n5590, n5592,
         n5593, n5597, n5598, n5600, n5601, n5605, n5606, n5608, n5609, n5613,
         n5614, n5616, n5617, n5625, n5626, n5628, n5629, n5633, n5634, n5636,
         n5637, n5641, n5642, n5644, n5645, n5649, n5650, n5652, n5653, n5666,
         n5667, n5669, n5670, n5674, n5675, n5677, n5678, n5682, n5683, n5685,
         n5686, n5690, n5691, n5693, n5694, n5702, n5703, n5705, n5706, n5710,
         n5711, n5713, n5714, n5718, n5719, n5721, n5722, n5726, n5727, n5729,
         n5730, n5738, n5739, n5741, n5742, n5746, n5747, n5749, n5750, n5754,
         n5755, n5757, n5758, n5762, n5763, n5765, n5766, n5774, n5775, n5777,
         n5778, n5782, n5783, n5785, n5786, n5790, n5791, n5793, n5794, n5798,
         n5799, n5801, n5802, n5815, n5816, n5818, n5819, n5823, n5824, n5826,
         n5827, n5831, n5832, n5834, n5835, n5839, n5840, n5842, n5843, n5851,
         n5852, n5854, n5855, n5859, n5860, n5862, n5863, n5867, n5868, n5870,
         n5871, n5875, n5876, n5878, n5879, n5889, n5890, n5892, n5893, n5897,
         n5898, n5900, n5901, n5905, n5906, n5908, n5909, n5913, n5914, n5916,
         n5917, n5925, n5926, n5928, n5929, n5933, n5934, n5936, n5937, n5941,
         n5942, n5944, n5945, n5949, n5950, n5954, n5955, n5956, n5957, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988;
  assign N147559 = DATA_IN[0];

  DFF_X1 \CACHE_MEM_reg[15][255]  ( .D(n14183), .CK(N28803), .Q(n5266), .QN(
        n6006) );
  DFF_X1 \CACHE_MEM_reg[15][254]  ( .D(n14182), .CK(N28803), .Q(n5255), .QN(
        n6022) );
  DFF_X1 \CACHE_MEM_reg[15][253]  ( .D(n14181), .CK(N28803), .Q(n5238), .QN(
        n6038) );
  DFF_X1 \CACHE_MEM_reg[15][252]  ( .D(n14180), .CK(N28803), .Q(n5227), .QN(
        n6054) );
  DFF_X1 \CACHE_MEM_reg[15][251]  ( .D(n14179), .CK(N28803), .Q(n5205), .QN(
        n6070) );
  DFF_X1 \CACHE_MEM_reg[15][250]  ( .D(n14178), .CK(N28803), .Q(n5194), .QN(
        n6086) );
  DFF_X1 \CACHE_MEM_reg[15][249]  ( .D(n14177), .CK(N28803), .Q(n5181), .QN(
        n6102) );
  DFF_X1 \CACHE_MEM_reg[15][248]  ( .D(n14176), .CK(N28803), .Q(n5166), .QN(
        n6118) );
  DFF_X1 \CACHE_MEM_reg[15][247]  ( .D(n14175), .CK(N28803), .Q(n5153), .QN(
        n6134) );
  DFF_X1 \CACHE_MEM_reg[15][246]  ( .D(n14174), .CK(N28803), .Q(n5142), .QN(
        n6150) );
  DFF_X1 \CACHE_MEM_reg[15][245]  ( .D(n14173), .CK(N28803), .Q(n5125), .QN(
        n6166) );
  DFF_X1 \CACHE_MEM_reg[15][244]  ( .D(n14172), .CK(N28803), .Q(n5114), .QN(
        n6182) );
  DFF_X1 \CACHE_MEM_reg[15][243]  ( .D(n14171), .CK(N28803), .Q(n5097), .QN(
        n6198) );
  DFF_X1 \CACHE_MEM_reg[15][242]  ( .D(n14170), .CK(N28803), .Q(n5086), .QN(
        n6214) );
  DFF_X1 \CACHE_MEM_reg[15][241]  ( .D(n14169), .CK(N28803), .Q(n5073), .QN(
        n6230) );
  DFF_X1 \CACHE_MEM_reg[15][240]  ( .D(n14168), .CK(N28803), .Q(n5721), .QN(
        n6246) );
  DFF_X1 \CACHE_MEM_reg[15][239]  ( .D(n14167), .CK(N28803), .Q(n5045), .QN(
        n6262) );
  DFF_X1 \CACHE_MEM_reg[15][238]  ( .D(n14166), .CK(N28803), .Q(n5032), .QN(
        n6278) );
  DFF_X1 \CACHE_MEM_reg[15][237]  ( .D(n14165), .CK(N28803), .Q(n5017), .QN(
        n6294) );
  DFF_X1 \CACHE_MEM_reg[15][236]  ( .D(n14164), .CK(N28803), .Q(n5004), .QN(
        n6310) );
  DFF_X1 \CACHE_MEM_reg[15][235]  ( .D(n14163), .CK(N28803), .Q(n4993), .QN(
        n6326) );
  DFF_X1 \CACHE_MEM_reg[15][234]  ( .D(n14162), .CK(N28803), .Q(n4976), .QN(
        n6342) );
  DFF_X1 \CACHE_MEM_reg[15][233]  ( .D(n14161), .CK(N28803), .Q(n4965), .QN(
        n6358) );
  DFF_X1 \CACHE_MEM_reg[15][232]  ( .D(n14160), .CK(N28803), .Q(n4948), .QN(
        n6374) );
  DFF_X1 \CACHE_MEM_reg[15][231]  ( .D(n14159), .CK(N28803), .Q(n4937), .QN(
        n6390) );
  DFF_X1 \CACHE_MEM_reg[15][230]  ( .D(n14158), .CK(N28803), .Q(n4924), .QN(
        n6406) );
  DFF_X1 \CACHE_MEM_reg[15][229]  ( .D(n14157), .CK(N28803), .Q(n4904), .QN(
        n6422) );
  DFF_X1 \CACHE_MEM_reg[15][228]  ( .D(n14156), .CK(N28803), .Q(n4891), .QN(
        n6438) );
  DFF_X1 \CACHE_MEM_reg[15][227]  ( .D(n14155), .CK(N28803), .Q(n4880), .QN(
        n6454) );
  DFF_X1 \CACHE_MEM_reg[15][226]  ( .D(n14154), .CK(N28803), .Q(n4863), .QN(
        n6470) );
  DFF_X1 \CACHE_MEM_reg[15][225]  ( .D(n14153), .CK(N28803), .Q(n4852), .QN(
        n6486) );
  DFF_X1 \CACHE_MEM_reg[15][224]  ( .D(n14152), .CK(N28803), .Q(n4835), .QN(
        n6502) );
  DFF_X1 \CACHE_MEM_reg[15][223]  ( .D(n14151), .CK(N28803), .Q(n5271), .QN(
        n6518) );
  DFF_X1 \CACHE_MEM_reg[15][222]  ( .D(n14150), .CK(N28803), .Q(n5258), .QN(
        n6534) );
  DFF_X1 \CACHE_MEM_reg[15][221]  ( .D(n14149), .CK(N28803), .Q(n5243), .QN(
        n6550) );
  DFF_X1 \CACHE_MEM_reg[15][220]  ( .D(n14148), .CK(N28803), .Q(n5230), .QN(
        n6566) );
  DFF_X1 \CACHE_MEM_reg[15][219]  ( .D(n14147), .CK(N28803), .Q(n5219), .QN(
        n6582) );
  DFF_X1 \CACHE_MEM_reg[15][218]  ( .D(n14146), .CK(N28803), .Q(n5197), .QN(
        n6598) );
  DFF_X1 \CACHE_MEM_reg[15][217]  ( .D(n14145), .CK(N28803), .Q(n5186), .QN(
        n6614) );
  DFF_X1 \CACHE_MEM_reg[15][216]  ( .D(n14144), .CK(N28803), .Q(n5169), .QN(
        n6630) );
  DFF_X1 \CACHE_MEM_reg[15][215]  ( .D(n14143), .CK(N28803), .Q(n5158), .QN(
        n6646) );
  DFF_X1 \CACHE_MEM_reg[15][214]  ( .D(n14142), .CK(N28803), .Q(n5145), .QN(
        n6662) );
  DFF_X1 \CACHE_MEM_reg[15][213]  ( .D(n14141), .CK(N28803), .Q(n5130), .QN(
        n6678) );
  DFF_X1 \CACHE_MEM_reg[15][212]  ( .D(n14140), .CK(N28803), .Q(n5117), .QN(
        n6694) );
  DFF_X1 \CACHE_MEM_reg[15][211]  ( .D(n14139), .CK(N28803), .Q(n5106), .QN(
        n6710) );
  DFF_X1 \CACHE_MEM_reg[15][210]  ( .D(n14138), .CK(N28803), .Q(n5089), .QN(
        n6726) );
  DFF_X1 \CACHE_MEM_reg[15][209]  ( .D(n14137), .CK(N28803), .Q(n5078), .QN(
        n6742) );
  DFF_X1 \CACHE_MEM_reg[15][208]  ( .D(n14136), .CK(N28803), .Q(n5056), .QN(
        n6758) );
  DFF_X1 \CACHE_MEM_reg[15][207]  ( .D(n14135), .CK(N28803), .Q(n5048), .QN(
        n6774) );
  DFF_X1 \CACHE_MEM_reg[15][206]  ( .D(n14134), .CK(N28803), .Q(n5037), .QN(
        n6790) );
  DFF_X1 \CACHE_MEM_reg[15][205]  ( .D(n14133), .CK(N28803), .Q(n5020), .QN(
        n6806) );
  DFF_X1 \CACHE_MEM_reg[15][204]  ( .D(n14132), .CK(N28803), .Q(n5009), .QN(
        n6822) );
  DFF_X1 \CACHE_MEM_reg[15][203]  ( .D(n14131), .CK(N28803), .Q(n4996), .QN(
        n6838) );
  DFF_X1 \CACHE_MEM_reg[15][202]  ( .D(n14130), .CK(N28803), .Q(n4981), .QN(
        n6854) );
  DFF_X1 \CACHE_MEM_reg[15][201]  ( .D(n14129), .CK(N28803), .Q(n4968), .QN(
        n6870) );
  DFF_X1 \CACHE_MEM_reg[15][200]  ( .D(n14128), .CK(N28803), .Q(n4957), .QN(
        n6886) );
  DFF_X1 \CACHE_MEM_reg[15][199]  ( .D(n14127), .CK(N28803), .Q(n4940), .QN(
        n6902) );
  DFF_X1 \CACHE_MEM_reg[15][198]  ( .D(n14126), .CK(N28803), .Q(n4929), .QN(
        n6918) );
  DFF_X1 \CACHE_MEM_reg[15][197]  ( .D(n14125), .CK(N28803), .Q(n4907), .QN(
        n6934) );
  DFF_X1 \CACHE_MEM_reg[15][196]  ( .D(n14124), .CK(N28803), .Q(n4896), .QN(
        n6950) );
  DFF_X1 \CACHE_MEM_reg[15][195]  ( .D(n14123), .CK(N28803), .Q(n4883), .QN(
        n6966) );
  DFF_X1 \CACHE_MEM_reg[15][194]  ( .D(n14122), .CK(N28803), .Q(n4868), .QN(
        n6982) );
  DFF_X1 \CACHE_MEM_reg[15][193]  ( .D(n14121), .CK(N28803), .Q(n4855), .QN(
        n6998) );
  DFF_X1 \CACHE_MEM_reg[15][192]  ( .D(n14120), .CK(N28803), .Q(n4844), .QN(
        n7014) );
  DFF_X1 \CACHE_MEM_reg[15][191]  ( .D(n14119), .CK(N28803), .Q(n5713), .QN(
        n7030) );
  DFF_X1 \CACHE_MEM_reg[15][190]  ( .D(n14118), .CK(N28803), .Q(n5702), .QN(
        n7046) );
  DFF_X1 \CACHE_MEM_reg[15][189]  ( .D(n14117), .CK(N28803), .Q(n5685), .QN(
        n7062) );
  DFF_X1 \CACHE_MEM_reg[15][188]  ( .D(n14116), .CK(N28803), .Q(n5674), .QN(
        n7078) );
  DFF_X1 \CACHE_MEM_reg[15][187]  ( .D(n14115), .CK(N28803), .Q(n5652), .QN(
        n7094) );
  DFF_X1 \CACHE_MEM_reg[15][186]  ( .D(n14114), .CK(N28803), .Q(n5641), .QN(
        n7110) );
  DFF_X1 \CACHE_MEM_reg[15][185]  ( .D(n14113), .CK(N28803), .Q(n5628), .QN(
        n7126) );
  DFF_X1 \CACHE_MEM_reg[15][184]  ( .D(n14112), .CK(N28803), .Q(n5613), .QN(
        n7142) );
  DFF_X1 \CACHE_MEM_reg[15][183]  ( .D(n14111), .CK(N28803), .Q(n5600), .QN(
        n7158) );
  DFF_X1 \CACHE_MEM_reg[15][182]  ( .D(n14110), .CK(N28803), .Q(n5589), .QN(
        n7174) );
  DFF_X1 \CACHE_MEM_reg[15][181]  ( .D(n14109), .CK(N28803), .Q(n5572), .QN(
        n7190) );
  DFF_X1 \CACHE_MEM_reg[15][180]  ( .D(n14108), .CK(N28803), .Q(n5561), .QN(
        n7206) );
  DFF_X1 \CACHE_MEM_reg[15][179]  ( .D(n14107), .CK(N28803), .Q(n5544), .QN(
        n7222) );
  DFF_X1 \CACHE_MEM_reg[15][178]  ( .D(n14106), .CK(N28803), .Q(n5533), .QN(
        n7238) );
  DFF_X1 \CACHE_MEM_reg[15][177]  ( .D(n14105), .CK(N28803), .Q(n5520), .QN(
        n7254) );
  DFF_X1 \CACHE_MEM_reg[15][176]  ( .D(n14104), .CK(N28803), .Q(n5500), .QN(
        n7270) );
  DFF_X1 \CACHE_MEM_reg[15][175]  ( .D(n14103), .CK(N28803), .Q(n5487), .QN(
        n7286) );
  DFF_X1 \CACHE_MEM_reg[15][174]  ( .D(n14102), .CK(N28803), .Q(n5476), .QN(
        n7302) );
  DFF_X1 \CACHE_MEM_reg[15][173]  ( .D(n14101), .CK(N28803), .Q(n5459), .QN(
        n7318) );
  DFF_X1 \CACHE_MEM_reg[15][172]  ( .D(n14100), .CK(N28803), .Q(n5448), .QN(
        n7334) );
  DFF_X1 \CACHE_MEM_reg[15][171]  ( .D(n14099), .CK(N28803), .Q(n5431), .QN(
        n7350) );
  DFF_X1 \CACHE_MEM_reg[15][170]  ( .D(n14098), .CK(N28803), .Q(n5420), .QN(
        n7366) );
  DFF_X1 \CACHE_MEM_reg[15][169]  ( .D(n14097), .CK(N28803), .Q(n5407), .QN(
        n7382) );
  DFF_X1 \CACHE_MEM_reg[15][168]  ( .D(n14096), .CK(N28803), .Q(n5392), .QN(
        n7398) );
  DFF_X1 \CACHE_MEM_reg[15][167]  ( .D(n14095), .CK(N28803), .Q(n5379), .QN(
        n7414) );
  DFF_X1 \CACHE_MEM_reg[15][166]  ( .D(n14094), .CK(N28803), .Q(n5368), .QN(
        n7430) );
  DFF_X1 \CACHE_MEM_reg[15][165]  ( .D(n14093), .CK(N28803), .Q(n5346), .QN(
        n7446) );
  DFF_X1 \CACHE_MEM_reg[15][164]  ( .D(n14092), .CK(N28803), .Q(n5335), .QN(
        n7462) );
  DFF_X1 \CACHE_MEM_reg[15][163]  ( .D(n14091), .CK(N28803), .Q(n5318), .QN(
        n7478) );
  DFF_X1 \CACHE_MEM_reg[15][162]  ( .D(n14090), .CK(N28803), .Q(n5307), .QN(
        n7494) );
  DFF_X1 \CACHE_MEM_reg[15][161]  ( .D(n14089), .CK(N28803), .Q(n5294), .QN(
        n7510) );
  DFF_X1 \CACHE_MEM_reg[15][160]  ( .D(n14088), .CK(N28803), .Q(n5279), .QN(
        n7526) );
  DFF_X1 \CACHE_MEM_reg[15][159]  ( .D(n14087), .CK(N28803), .Q(n5718), .QN(
        n7542) );
  DFF_X1 \CACHE_MEM_reg[15][158]  ( .D(n14086), .CK(N28803), .Q(n5726), .QN(
        n7558) );
  DFF_X1 \CACHE_MEM_reg[15][157]  ( .D(n14085), .CK(N28803), .Q(n5690), .QN(
        n7574) );
  DFF_X1 \CACHE_MEM_reg[15][156]  ( .D(n14084), .CK(N28803), .Q(n5677), .QN(
        n7590) );
  DFF_X1 \CACHE_MEM_reg[15][155]  ( .D(n14083), .CK(N28803), .Q(n5666), .QN(
        n7606) );
  DFF_X1 \CACHE_MEM_reg[15][154]  ( .D(n14082), .CK(N28803), .Q(n5644), .QN(
        n7622) );
  DFF_X1 \CACHE_MEM_reg[15][153]  ( .D(n14081), .CK(N28803), .Q(n5633), .QN(
        n7638) );
  DFF_X1 \CACHE_MEM_reg[15][152]  ( .D(n14080), .CK(N28803), .Q(n5616), .QN(
        n7654) );
  DFF_X1 \CACHE_MEM_reg[15][151]  ( .D(n14079), .CK(N28803), .Q(n5605), .QN(
        n7670) );
  DFF_X1 \CACHE_MEM_reg[15][150]  ( .D(n14078), .CK(N28803), .Q(n5592), .QN(
        n7686) );
  DFF_X1 \CACHE_MEM_reg[15][149]  ( .D(n14077), .CK(N28803), .Q(n5577), .QN(
        n7702) );
  DFF_X1 \CACHE_MEM_reg[15][148]  ( .D(n14076), .CK(N28803), .Q(n5564), .QN(
        n7718) );
  DFF_X1 \CACHE_MEM_reg[15][147]  ( .D(n14075), .CK(N28803), .Q(n5553), .QN(
        n7734) );
  DFF_X1 \CACHE_MEM_reg[15][146]  ( .D(n14074), .CK(N28803), .Q(n5536), .QN(
        n7750) );
  DFF_X1 \CACHE_MEM_reg[15][145]  ( .D(n14073), .CK(N28803), .Q(n5525), .QN(
        n7766) );
  DFF_X1 \CACHE_MEM_reg[15][144]  ( .D(n14072), .CK(N28803), .Q(n5503), .QN(
        n7782) );
  DFF_X1 \CACHE_MEM_reg[15][143]  ( .D(n14071), .CK(N28803), .Q(n5492), .QN(
        n7798) );
  DFF_X1 \CACHE_MEM_reg[15][142]  ( .D(n14070), .CK(N28803), .Q(n5479), .QN(
        n7814) );
  DFF_X1 \CACHE_MEM_reg[15][141]  ( .D(n14069), .CK(N28803), .Q(n5464), .QN(
        n7830) );
  DFF_X1 \CACHE_MEM_reg[15][140]  ( .D(n14068), .CK(N28803), .Q(n5451), .QN(
        n7846) );
  DFF_X1 \CACHE_MEM_reg[15][139]  ( .D(n14067), .CK(N28803), .Q(n5440), .QN(
        n7862) );
  DFF_X1 \CACHE_MEM_reg[15][138]  ( .D(n14066), .CK(N28803), .Q(n5423), .QN(
        n7878) );
  DFF_X1 \CACHE_MEM_reg[15][137]  ( .D(n14065), .CK(N28803), .Q(n5412), .QN(
        n7894) );
  DFF_X1 \CACHE_MEM_reg[15][136]  ( .D(n14064), .CK(N28803), .Q(n5395), .QN(
        n7910) );
  DFF_X1 \CACHE_MEM_reg[15][135]  ( .D(n14063), .CK(N28803), .Q(n5384), .QN(
        n7926) );
  DFF_X1 \CACHE_MEM_reg[15][134]  ( .D(n14062), .CK(N28803), .Q(n5371), .QN(
        n7942) );
  DFF_X1 \CACHE_MEM_reg[15][133]  ( .D(n14061), .CK(N28803), .Q(n5351), .QN(
        n7958) );
  DFF_X1 \CACHE_MEM_reg[15][132]  ( .D(n14060), .CK(N28803), .Q(n5338), .QN(
        n7974) );
  DFF_X1 \CACHE_MEM_reg[15][131]  ( .D(n14059), .CK(N28803), .Q(n5327), .QN(
        n7990) );
  DFF_X1 \CACHE_MEM_reg[15][130]  ( .D(n14058), .CK(N28803), .Q(n5310), .QN(
        n8006) );
  DFF_X1 \CACHE_MEM_reg[15][129]  ( .D(n14057), .CK(N28803), .Q(n5299), .QN(
        n8022) );
  DFF_X1 \CACHE_MEM_reg[15][128]  ( .D(n14056), .CK(N28803), .Q(n5282), .QN(
        n8038) );
  DFF_X1 \CACHE_MEM_reg[15][127]  ( .D(n14055), .CK(N28803), .Q(n4377), .QN(
        n8054) );
  DFF_X1 \CACHE_MEM_reg[15][126]  ( .D(n14054), .CK(N28803), .Q(n4364), .QN(
        n8070) );
  DFF_X1 \CACHE_MEM_reg[15][125]  ( .D(n14053), .CK(N28803), .Q(n4344), .QN(
        n8086) );
  DFF_X1 \CACHE_MEM_reg[15][124]  ( .D(n14052), .CK(N28803), .Q(n4328), .QN(
        n8102) );
  DFF_X1 \CACHE_MEM_reg[15][123]  ( .D(n14051), .CK(N28803), .Q(n4303), .QN(
        n8118) );
  DFF_X1 \CACHE_MEM_reg[15][122]  ( .D(n14050), .CK(N28803), .Q(n4287), .QN(
        n8134) );
  DFF_X1 \CACHE_MEM_reg[15][121]  ( .D(n14049), .CK(N28803), .Q(n4267), .QN(
        n8150) );
  DFF_X1 \CACHE_MEM_reg[15][120]  ( .D(n14048), .CK(N28803), .Q(n4251), .QN(
        n8166) );
  DFF_X1 \CACHE_MEM_reg[15][119]  ( .D(n14047), .CK(N28803), .Q(n4231), .QN(
        n8182) );
  DFF_X1 \CACHE_MEM_reg[15][118]  ( .D(n14046), .CK(N28803), .Q(n4215), .QN(
        n8198) );
  DFF_X1 \CACHE_MEM_reg[15][117]  ( .D(n14045), .CK(N28803), .Q(n4195), .QN(
        n8214) );
  DFF_X1 \CACHE_MEM_reg[15][116]  ( .D(n14044), .CK(N28803), .Q(n4179), .QN(
        n8230) );
  DFF_X1 \CACHE_MEM_reg[15][115]  ( .D(n14043), .CK(N28803), .Q(n4154), .QN(
        n8246) );
  DFF_X1 \CACHE_MEM_reg[15][114]  ( .D(n14042), .CK(N28803), .Q(n4138), .QN(
        n8262) );
  DFF_X1 \CACHE_MEM_reg[15][113]  ( .D(n14041), .CK(N28803), .Q(n4118), .QN(
        n8278) );
  DFF_X1 \CACHE_MEM_reg[15][112]  ( .D(n14040), .CK(N28803), .Q(n4102), .QN(
        n8294) );
  DFF_X1 \CACHE_MEM_reg[15][111]  ( .D(n14039), .CK(N28803), .Q(n4082), .QN(
        n8310) );
  DFF_X1 \CACHE_MEM_reg[15][110]  ( .D(n14038), .CK(N28803), .Q(n4066), .QN(
        n8326) );
  DFF_X1 \CACHE_MEM_reg[15][109]  ( .D(n14037), .CK(N28803), .Q(n4046), .QN(
        n8342) );
  DFF_X1 \CACHE_MEM_reg[15][108]  ( .D(n14036), .CK(N28803), .Q(n4030), .QN(
        n8358) );
  DFF_X1 \CACHE_MEM_reg[15][107]  ( .D(n14035), .CK(N28803), .Q(n4005), .QN(
        n8374) );
  DFF_X1 \CACHE_MEM_reg[15][106]  ( .D(n14034), .CK(N28803), .Q(n3989), .QN(
        n8390) );
  DFF_X1 \CACHE_MEM_reg[15][105]  ( .D(n14033), .CK(N28803), .Q(n3969), .QN(
        n8406) );
  DFF_X1 \CACHE_MEM_reg[15][104]  ( .D(n14032), .CK(N28803), .Q(n3953), .QN(
        n8422) );
  DFF_X1 \CACHE_MEM_reg[15][103]  ( .D(n14031), .CK(N28803), .Q(n3933), .QN(
        n8438) );
  DFF_X1 \CACHE_MEM_reg[15][102]  ( .D(n14030), .CK(N28803), .Q(n3917), .QN(
        n8454) );
  DFF_X1 \CACHE_MEM_reg[15][101]  ( .D(n14029), .CK(N28803), .Q(n3897), .QN(
        n8470) );
  DFF_X1 \CACHE_MEM_reg[15][100]  ( .D(n14028), .CK(N28803), .Q(n3881), .QN(
        n8486) );
  DFF_X1 \CACHE_MEM_reg[15][99]  ( .D(n14027), .CK(N28803), .Q(n3856), .QN(
        n8502) );
  DFF_X1 \CACHE_MEM_reg[15][98]  ( .D(n14026), .CK(N28803), .Q(n3840), .QN(
        n8518) );
  DFF_X1 \CACHE_MEM_reg[15][97]  ( .D(n14025), .CK(N28803), .Q(n3820), .QN(
        n8534) );
  DFF_X1 \CACHE_MEM_reg[15][96]  ( .D(n14024), .CK(N28803), .Q(n3804), .QN(
        n8550) );
  DFF_X1 \CACHE_MEM_reg[15][95]  ( .D(n14023), .CK(N28803), .Q(n4380), .QN(
        n8566) );
  DFF_X1 \CACHE_MEM_reg[15][94]  ( .D(n14022), .CK(N28803), .Q(n4369), .QN(
        n8582) );
  DFF_X1 \CACHE_MEM_reg[15][93]  ( .D(n14021), .CK(N28803), .Q(n4349), .QN(
        n8598) );
  DFF_X1 \CACHE_MEM_reg[15][92]  ( .D(n14020), .CK(N28803), .Q(n4333), .QN(
        n8614) );
  DFF_X1 \CACHE_MEM_reg[15][91]  ( .D(n14019), .CK(N28803), .Q(n4308), .QN(
        n8630) );
  DFF_X1 \CACHE_MEM_reg[15][90]  ( .D(n14018), .CK(N28803), .Q(n4292), .QN(
        n8646) );
  DFF_X1 \CACHE_MEM_reg[15][89]  ( .D(n14017), .CK(N28803), .Q(n4272), .QN(
        n8662) );
  DFF_X1 \CACHE_MEM_reg[15][88]  ( .D(n14016), .CK(N28803), .Q(n4256), .QN(
        n8678) );
  DFF_X1 \CACHE_MEM_reg[15][87]  ( .D(n14015), .CK(N28803), .Q(n4236), .QN(
        n8694) );
  DFF_X1 \CACHE_MEM_reg[15][86]  ( .D(n14014), .CK(N28803), .Q(n4220), .QN(
        n8710) );
  DFF_X1 \CACHE_MEM_reg[15][85]  ( .D(n14013), .CK(N28803), .Q(n4200), .QN(
        n8726) );
  DFF_X1 \CACHE_MEM_reg[15][84]  ( .D(n14012), .CK(N28803), .Q(n4184), .QN(
        n8742) );
  DFF_X1 \CACHE_MEM_reg[15][83]  ( .D(n14011), .CK(N28803), .Q(n4159), .QN(
        n8758) );
  DFF_X1 \CACHE_MEM_reg[15][82]  ( .D(n14010), .CK(N28803), .Q(n4143), .QN(
        n8774) );
  DFF_X1 \CACHE_MEM_reg[15][81]  ( .D(n14009), .CK(N28803), .Q(n4123), .QN(
        n8790) );
  DFF_X1 \CACHE_MEM_reg[15][80]  ( .D(n14008), .CK(N28803), .Q(n4107), .QN(
        n8806) );
  DFF_X1 \CACHE_MEM_reg[15][79]  ( .D(n14007), .CK(N28803), .Q(n4087), .QN(
        n8822) );
  DFF_X1 \CACHE_MEM_reg[15][78]  ( .D(n14006), .CK(N28803), .Q(n4071), .QN(
        n8838) );
  DFF_X1 \CACHE_MEM_reg[15][77]  ( .D(n14005), .CK(N28803), .Q(n4051), .QN(
        n8854) );
  DFF_X1 \CACHE_MEM_reg[15][76]  ( .D(n14004), .CK(N28803), .Q(n4035), .QN(
        n8870) );
  DFF_X1 \CACHE_MEM_reg[15][75]  ( .D(n14003), .CK(N28803), .Q(n4010), .QN(
        n8886) );
  DFF_X1 \CACHE_MEM_reg[15][74]  ( .D(n14002), .CK(N28803), .Q(n3994), .QN(
        n8902) );
  DFF_X1 \CACHE_MEM_reg[15][73]  ( .D(n14001), .CK(N28803), .Q(n3974), .QN(
        n8918) );
  DFF_X1 \CACHE_MEM_reg[15][72]  ( .D(n14000), .CK(N28803), .Q(n3958), .QN(
        n8934) );
  DFF_X1 \CACHE_MEM_reg[15][71]  ( .D(n13999), .CK(N28803), .Q(n3938), .QN(
        n8950) );
  DFF_X1 \CACHE_MEM_reg[15][70]  ( .D(n13998), .CK(N28803), .Q(n3922), .QN(
        n8966) );
  DFF_X1 \CACHE_MEM_reg[15][69]  ( .D(n13997), .CK(N28803), .Q(n3902), .QN(
        n8982) );
  DFF_X1 \CACHE_MEM_reg[15][68]  ( .D(n13996), .CK(N28803), .Q(n3886), .QN(
        n8998) );
  DFF_X1 \CACHE_MEM_reg[15][67]  ( .D(n13995), .CK(N28803), .Q(n3861), .QN(
        n9014) );
  DFF_X1 \CACHE_MEM_reg[15][66]  ( .D(n13994), .CK(N28803), .Q(n3845), .QN(
        n9030) );
  DFF_X1 \CACHE_MEM_reg[15][65]  ( .D(n13993), .CK(N28803), .Q(n3825), .QN(
        n9046) );
  DFF_X1 \CACHE_MEM_reg[15][64]  ( .D(n13992), .CK(N28803), .Q(n3809), .QN(
        n9062) );
  DFF_X1 \CACHE_MEM_reg[15][63]  ( .D(n13991), .CK(N28803), .Q(n4824), .QN(
        n9078) );
  DFF_X1 \CACHE_MEM_reg[15][62]  ( .D(n13990), .CK(N28803), .Q(n4811), .QN(
        n9094) );
  DFF_X1 \CACHE_MEM_reg[15][61]  ( .D(n13989), .CK(N28803), .Q(n4796), .QN(
        n9110) );
  DFF_X1 \CACHE_MEM_reg[15][60]  ( .D(n13988), .CK(N28803), .Q(n4783), .QN(
        n9126) );
  DFF_X1 \CACHE_MEM_reg[15][59]  ( .D(n13987), .CK(N28803), .Q(n4772), .QN(
        n9142) );
  DFF_X1 \CACHE_MEM_reg[15][58]  ( .D(n13986), .CK(N28803), .Q(n4750), .QN(
        n9158) );
  DFF_X1 \CACHE_MEM_reg[15][57]  ( .D(n13985), .CK(N28803), .Q(n4739), .QN(
        n9174) );
  DFF_X1 \CACHE_MEM_reg[15][56]  ( .D(n13984), .CK(N28803), .Q(n4722), .QN(
        n9190) );
  DFF_X1 \CACHE_MEM_reg[15][55]  ( .D(n13983), .CK(N28803), .Q(n4711), .QN(
        n9206) );
  DFF_X1 \CACHE_MEM_reg[15][54]  ( .D(n13982), .CK(N28803), .Q(n4698), .QN(
        n9222) );
  DFF_X1 \CACHE_MEM_reg[15][53]  ( .D(n13981), .CK(N28803), .Q(n4683), .QN(
        n9238) );
  DFF_X1 \CACHE_MEM_reg[15][52]  ( .D(n13980), .CK(N28803), .Q(n4670), .QN(
        n9254) );
  DFF_X1 \CACHE_MEM_reg[15][51]  ( .D(n13979), .CK(N28803), .Q(n4659), .QN(
        n9270) );
  DFF_X1 \CACHE_MEM_reg[15][50]  ( .D(n13978), .CK(N28803), .Q(n4642), .QN(
        n9286) );
  DFF_X1 \CACHE_MEM_reg[15][49]  ( .D(n13977), .CK(N28803), .Q(n4631), .QN(
        n9302) );
  DFF_X1 \CACHE_MEM_reg[15][48]  ( .D(n13976), .CK(N28803), .Q(n4609), .QN(
        n9318) );
  DFF_X1 \CACHE_MEM_reg[15][47]  ( .D(n13975), .CK(N28803), .Q(n4598), .QN(
        n9334) );
  DFF_X1 \CACHE_MEM_reg[15][46]  ( .D(n13974), .CK(N28803), .Q(n4585), .QN(
        n9350) );
  DFF_X1 \CACHE_MEM_reg[15][45]  ( .D(n13973), .CK(N28803), .Q(n4570), .QN(
        n9366) );
  DFF_X1 \CACHE_MEM_reg[15][44]  ( .D(n13972), .CK(N28803), .Q(n4557), .QN(
        n9382) );
  DFF_X1 \CACHE_MEM_reg[15][43]  ( .D(n13971), .CK(N28803), .Q(n4546), .QN(
        n9398) );
  DFF_X1 \CACHE_MEM_reg[15][42]  ( .D(n13970), .CK(N28803), .Q(n4529), .QN(
        n9414) );
  DFF_X1 \CACHE_MEM_reg[15][41]  ( .D(n13969), .CK(N28803), .Q(n4518), .QN(
        n9430) );
  DFF_X1 \CACHE_MEM_reg[15][40]  ( .D(n13968), .CK(N28803), .Q(n4501), .QN(
        n9446) );
  DFF_X1 \CACHE_MEM_reg[15][39]  ( .D(n13967), .CK(N28803), .Q(n4490), .QN(
        n9462) );
  DFF_X1 \CACHE_MEM_reg[15][38]  ( .D(n13966), .CK(N28803), .Q(n4477), .QN(
        n9478) );
  DFF_X1 \CACHE_MEM_reg[15][37]  ( .D(n13965), .CK(N28803), .Q(n4457), .QN(
        n9494) );
  DFF_X1 \CACHE_MEM_reg[15][36]  ( .D(n13964), .CK(N28803), .Q(n4444), .QN(
        n9510) );
  DFF_X1 \CACHE_MEM_reg[15][35]  ( .D(n13963), .CK(N28803), .Q(n4433), .QN(
        n9526) );
  DFF_X1 \CACHE_MEM_reg[15][34]  ( .D(n13962), .CK(N28803), .Q(n4416), .QN(
        n9542) );
  DFF_X1 \CACHE_MEM_reg[15][33]  ( .D(n13961), .CK(N28803), .Q(n4405), .QN(
        n9558) );
  DFF_X1 \CACHE_MEM_reg[15][32]  ( .D(n13960), .CK(N28803), .Q(n4388), .QN(
        n9574) );
  DFF_X1 \CACHE_MEM_reg[15][31]  ( .D(n13959), .CK(N28803), .Q(n4827), .QN(
        n9590) );
  DFF_X1 \CACHE_MEM_reg[15][30]  ( .D(n13958), .CK(N28803), .Q(n4816), .QN(
        n9606) );
  DFF_X1 \CACHE_MEM_reg[15][29]  ( .D(n13957), .CK(N28803), .Q(n4799), .QN(
        n9622) );
  DFF_X1 \CACHE_MEM_reg[15][28]  ( .D(n13956), .CK(N28803), .Q(n4788), .QN(
        n9638) );
  DFF_X1 \CACHE_MEM_reg[15][27]  ( .D(n13955), .CK(N28803), .Q(n4775), .QN(
        n9654) );
  DFF_X1 \CACHE_MEM_reg[15][26]  ( .D(n13954), .CK(N28803), .Q(n4755), .QN(
        n9670) );
  DFF_X1 \CACHE_MEM_reg[15][25]  ( .D(n13953), .CK(N28803), .Q(n4742), .QN(
        n9686) );
  DFF_X1 \CACHE_MEM_reg[15][24]  ( .D(n13952), .CK(N28803), .Q(n4731), .QN(
        n9702) );
  DFF_X1 \CACHE_MEM_reg[15][23]  ( .D(n13951), .CK(N28803), .Q(n4714), .QN(
        n9718) );
  DFF_X1 \CACHE_MEM_reg[15][22]  ( .D(n13950), .CK(N28803), .Q(n4703), .QN(
        n9734) );
  DFF_X1 \CACHE_MEM_reg[15][21]  ( .D(n13949), .CK(N28803), .Q(n4686), .QN(
        n9750) );
  DFF_X1 \CACHE_MEM_reg[15][20]  ( .D(n13948), .CK(N28803), .Q(n4675), .QN(
        n9766) );
  DFF_X1 \CACHE_MEM_reg[15][19]  ( .D(n13947), .CK(N28803), .Q(n4662), .QN(
        n9782) );
  DFF_X1 \CACHE_MEM_reg[15][18]  ( .D(n13946), .CK(N28803), .Q(n4647), .QN(
        n9798) );
  DFF_X1 \CACHE_MEM_reg[15][17]  ( .D(n13945), .CK(N28803), .Q(n4634), .QN(
        n9814) );
  DFF_X1 \CACHE_MEM_reg[15][16]  ( .D(n13944), .CK(N28803), .Q(n4623), .QN(
        n9830) );
  DFF_X1 \CACHE_MEM_reg[15][15]  ( .D(n13943), .CK(N28803), .Q(n4601), .QN(
        n9846) );
  DFF_X1 \CACHE_MEM_reg[15][14]  ( .D(n13942), .CK(N28803), .Q(n4590), .QN(
        n9862) );
  DFF_X1 \CACHE_MEM_reg[15][13]  ( .D(n13941), .CK(N28803), .Q(n4573), .QN(
        n9878) );
  DFF_X1 \CACHE_MEM_reg[15][12]  ( .D(n13940), .CK(N28803), .Q(n4562), .QN(
        n9894) );
  DFF_X1 \CACHE_MEM_reg[15][11]  ( .D(n13939), .CK(N28803), .Q(n4549), .QN(
        n9910) );
  DFF_X1 \CACHE_MEM_reg[15][10]  ( .D(n13938), .CK(N28803), .Q(n4534), .QN(
        n9926) );
  DFF_X1 \CACHE_MEM_reg[15][9]  ( .D(n13937), .CK(N28803), .Q(n4521), .QN(
        n9942) );
  DFF_X1 \CACHE_MEM_reg[15][8]  ( .D(n13936), .CK(N28803), .Q(n4510), .QN(
        n9958) );
  DFF_X1 \CACHE_MEM_reg[15][7]  ( .D(n13935), .CK(N28803), .Q(n4493), .QN(
        n9974) );
  DFF_X1 \CACHE_MEM_reg[15][6]  ( .D(n13934), .CK(N28803), .Q(n4482), .QN(
        n9990) );
  DFF_X1 \CACHE_MEM_reg[15][5]  ( .D(n13933), .CK(N28803), .Q(n4460), .QN(
        n10006) );
  DFF_X1 \CACHE_MEM_reg[15][4]  ( .D(n13932), .CK(N28803), .Q(n4449), .QN(
        n10022) );
  DFF_X1 \CACHE_MEM_reg[15][3]  ( .D(n13931), .CK(N28803), .Q(n4436), .QN(
        n10038) );
  DFF_X1 \CACHE_MEM_reg[15][2]  ( .D(n13930), .CK(N28803), .Q(n4421), .QN(
        n10054) );
  DFF_X1 \CACHE_MEM_reg[15][1]  ( .D(n13929), .CK(N28803), .Q(n4408), .QN(
        n10070) );
  DFF_X1 \CACHE_MEM_reg[15][0]  ( .D(n13928), .CK(N28803), .Q(n4397), .QN(
        n10086) );
  DFF_X1 \CACHE_MEM_reg[14][255]  ( .D(n13927), .CK(N28803), .QN(n6002) );
  DFF_X1 \CACHE_MEM_reg[14][254]  ( .D(n13926), .CK(N28803), .QN(n6018) );
  DFF_X1 \CACHE_MEM_reg[14][253]  ( .D(n13925), .CK(N28803), .QN(n6034) );
  DFF_X1 \CACHE_MEM_reg[14][252]  ( .D(n13924), .CK(N28803), .QN(n6050) );
  DFF_X1 \CACHE_MEM_reg[14][251]  ( .D(n13923), .CK(N28803), .QN(n6066) );
  DFF_X1 \CACHE_MEM_reg[14][250]  ( .D(n13922), .CK(N28803), .QN(n6082) );
  DFF_X1 \CACHE_MEM_reg[14][249]  ( .D(n13921), .CK(N28803), .QN(n6098) );
  DFF_X1 \CACHE_MEM_reg[14][248]  ( .D(n13920), .CK(N28803), .QN(n6114) );
  DFF_X1 \CACHE_MEM_reg[14][247]  ( .D(n13919), .CK(N28803), .QN(n6130) );
  DFF_X1 \CACHE_MEM_reg[14][246]  ( .D(n13918), .CK(N28803), .QN(n6146) );
  DFF_X1 \CACHE_MEM_reg[14][245]  ( .D(n13917), .CK(N28803), .QN(n6162) );
  DFF_X1 \CACHE_MEM_reg[14][244]  ( .D(n13916), .CK(N28803), .QN(n6178) );
  DFF_X1 \CACHE_MEM_reg[14][243]  ( .D(n13915), .CK(N28803), .QN(n6194) );
  DFF_X1 \CACHE_MEM_reg[14][242]  ( .D(n13914), .CK(N28803), .QN(n6210) );
  DFF_X1 \CACHE_MEM_reg[14][241]  ( .D(n13913), .CK(N28803), .QN(n6226) );
  DFF_X1 \CACHE_MEM_reg[14][240]  ( .D(n13912), .CK(N28803), .QN(n6242) );
  DFF_X1 \CACHE_MEM_reg[14][239]  ( .D(n13911), .CK(N28803), .QN(n6258) );
  DFF_X1 \CACHE_MEM_reg[14][238]  ( .D(n13910), .CK(N28803), .QN(n6274) );
  DFF_X1 \CACHE_MEM_reg[14][237]  ( .D(n13909), .CK(N28803), .QN(n6290) );
  DFF_X1 \CACHE_MEM_reg[14][236]  ( .D(n13908), .CK(N28803), .QN(n6306) );
  DFF_X1 \CACHE_MEM_reg[14][235]  ( .D(n13907), .CK(N28803), .QN(n6322) );
  DFF_X1 \CACHE_MEM_reg[14][234]  ( .D(n13906), .CK(N28803), .QN(n6338) );
  DFF_X1 \CACHE_MEM_reg[14][233]  ( .D(n13905), .CK(N28803), .QN(n6354) );
  DFF_X1 \CACHE_MEM_reg[14][232]  ( .D(n13904), .CK(N28803), .QN(n6370) );
  DFF_X1 \CACHE_MEM_reg[14][231]  ( .D(n13903), .CK(N28803), .QN(n6386) );
  DFF_X1 \CACHE_MEM_reg[14][230]  ( .D(n13902), .CK(N28803), .QN(n6402) );
  DFF_X1 \CACHE_MEM_reg[14][229]  ( .D(n13901), .CK(N28803), .QN(n6418) );
  DFF_X1 \CACHE_MEM_reg[14][228]  ( .D(n13900), .CK(N28803), .QN(n6434) );
  DFF_X1 \CACHE_MEM_reg[14][227]  ( .D(n13899), .CK(N28803), .QN(n6450) );
  DFF_X1 \CACHE_MEM_reg[14][226]  ( .D(n13898), .CK(N28803), .QN(n6466) );
  DFF_X1 \CACHE_MEM_reg[14][225]  ( .D(n13897), .CK(N28803), .QN(n6482) );
  DFF_X1 \CACHE_MEM_reg[14][224]  ( .D(n13896), .CK(N28803), .QN(n6498) );
  DFF_X1 \CACHE_MEM_reg[14][223]  ( .D(n13895), .CK(N28803), .QN(n6514) );
  DFF_X1 \CACHE_MEM_reg[14][222]  ( .D(n13894), .CK(N28803), .QN(n6530) );
  DFF_X1 \CACHE_MEM_reg[14][221]  ( .D(n13893), .CK(N28803), .QN(n6546) );
  DFF_X1 \CACHE_MEM_reg[14][220]  ( .D(n13892), .CK(N28803), .QN(n6562) );
  DFF_X1 \CACHE_MEM_reg[14][219]  ( .D(n13891), .CK(N28803), .QN(n6578) );
  DFF_X1 \CACHE_MEM_reg[14][218]  ( .D(n13890), .CK(N28803), .QN(n6594) );
  DFF_X1 \CACHE_MEM_reg[14][217]  ( .D(n13889), .CK(N28803), .QN(n6610) );
  DFF_X1 \CACHE_MEM_reg[14][216]  ( .D(n13888), .CK(N28803), .QN(n6626) );
  DFF_X1 \CACHE_MEM_reg[14][215]  ( .D(n13887), .CK(N28803), .QN(n6642) );
  DFF_X1 \CACHE_MEM_reg[14][214]  ( .D(n13886), .CK(N28803), .QN(n6658) );
  DFF_X1 \CACHE_MEM_reg[14][213]  ( .D(n13885), .CK(N28803), .QN(n6674) );
  DFF_X1 \CACHE_MEM_reg[14][212]  ( .D(n13884), .CK(N28803), .QN(n6690) );
  DFF_X1 \CACHE_MEM_reg[14][211]  ( .D(n13883), .CK(N28803), .QN(n6706) );
  DFF_X1 \CACHE_MEM_reg[14][210]  ( .D(n13882), .CK(N28803), .QN(n6722) );
  DFF_X1 \CACHE_MEM_reg[14][209]  ( .D(n13881), .CK(N28803), .QN(n6738) );
  DFF_X1 \CACHE_MEM_reg[14][208]  ( .D(n13880), .CK(N28803), .QN(n6754) );
  DFF_X1 \CACHE_MEM_reg[14][207]  ( .D(n13879), .CK(N28803), .QN(n6770) );
  DFF_X1 \CACHE_MEM_reg[14][206]  ( .D(n13878), .CK(N28803), .QN(n6786) );
  DFF_X1 \CACHE_MEM_reg[14][205]  ( .D(n13877), .CK(N28803), .QN(n6802) );
  DFF_X1 \CACHE_MEM_reg[14][204]  ( .D(n13876), .CK(N28803), .QN(n6818) );
  DFF_X1 \CACHE_MEM_reg[14][203]  ( .D(n13875), .CK(N28803), .QN(n6834) );
  DFF_X1 \CACHE_MEM_reg[14][202]  ( .D(n13874), .CK(N28803), .QN(n6850) );
  DFF_X1 \CACHE_MEM_reg[14][201]  ( .D(n13873), .CK(N28803), .QN(n6866) );
  DFF_X1 \CACHE_MEM_reg[14][200]  ( .D(n13872), .CK(N28803), .QN(n6882) );
  DFF_X1 \CACHE_MEM_reg[14][199]  ( .D(n13871), .CK(N28803), .QN(n6898) );
  DFF_X1 \CACHE_MEM_reg[14][198]  ( .D(n13870), .CK(N28803), .QN(n6914) );
  DFF_X1 \CACHE_MEM_reg[14][197]  ( .D(n13869), .CK(N28803), .QN(n6930) );
  DFF_X1 \CACHE_MEM_reg[14][196]  ( .D(n13868), .CK(N28803), .QN(n6946) );
  DFF_X1 \CACHE_MEM_reg[14][195]  ( .D(n13867), .CK(N28803), .QN(n6962) );
  DFF_X1 \CACHE_MEM_reg[14][194]  ( .D(n13866), .CK(N28803), .QN(n6978) );
  DFF_X1 \CACHE_MEM_reg[14][193]  ( .D(n13865), .CK(N28803), .QN(n6994) );
  DFF_X1 \CACHE_MEM_reg[14][192]  ( .D(n13864), .CK(N28803), .QN(n7010) );
  DFF_X1 \CACHE_MEM_reg[14][191]  ( .D(n13863), .CK(N28803), .QN(n7026) );
  DFF_X1 \CACHE_MEM_reg[14][190]  ( .D(n13862), .CK(N28803), .QN(n7042) );
  DFF_X1 \CACHE_MEM_reg[14][189]  ( .D(n13861), .CK(N28803), .QN(n7058) );
  DFF_X1 \CACHE_MEM_reg[14][188]  ( .D(n13860), .CK(N28803), .QN(n7074) );
  DFF_X1 \CACHE_MEM_reg[14][187]  ( .D(n13859), .CK(N28803), .QN(n7090) );
  DFF_X1 \CACHE_MEM_reg[14][186]  ( .D(n13858), .CK(N28803), .QN(n7106) );
  DFF_X1 \CACHE_MEM_reg[14][185]  ( .D(n13857), .CK(N28803), .QN(n7122) );
  DFF_X1 \CACHE_MEM_reg[14][184]  ( .D(n13856), .CK(N28803), .QN(n7138) );
  DFF_X1 \CACHE_MEM_reg[14][183]  ( .D(n13855), .CK(N28803), .QN(n7154) );
  DFF_X1 \CACHE_MEM_reg[14][182]  ( .D(n13854), .CK(N28803), .QN(n7170) );
  DFF_X1 \CACHE_MEM_reg[14][181]  ( .D(n13853), .CK(N28803), .QN(n7186) );
  DFF_X1 \CACHE_MEM_reg[14][180]  ( .D(n13852), .CK(N28803), .QN(n7202) );
  DFF_X1 \CACHE_MEM_reg[14][179]  ( .D(n13851), .CK(N28803), .QN(n7218) );
  DFF_X1 \CACHE_MEM_reg[14][178]  ( .D(n13850), .CK(N28803), .QN(n7234) );
  DFF_X1 \CACHE_MEM_reg[14][177]  ( .D(n13849), .CK(N28803), .QN(n7250) );
  DFF_X1 \CACHE_MEM_reg[14][176]  ( .D(n13848), .CK(N28803), .QN(n7266) );
  DFF_X1 \CACHE_MEM_reg[14][175]  ( .D(n13847), .CK(N28803), .QN(n7282) );
  DFF_X1 \CACHE_MEM_reg[14][174]  ( .D(n13846), .CK(N28803), .QN(n7298) );
  DFF_X1 \CACHE_MEM_reg[14][173]  ( .D(n13845), .CK(N28803), .QN(n7314) );
  DFF_X1 \CACHE_MEM_reg[14][172]  ( .D(n13844), .CK(N28803), .QN(n7330) );
  DFF_X1 \CACHE_MEM_reg[14][171]  ( .D(n13843), .CK(N28803), .QN(n7346) );
  DFF_X1 \CACHE_MEM_reg[14][170]  ( .D(n13842), .CK(N28803), .QN(n7362) );
  DFF_X1 \CACHE_MEM_reg[14][169]  ( .D(n13841), .CK(N28803), .QN(n7378) );
  DFF_X1 \CACHE_MEM_reg[14][168]  ( .D(n13840), .CK(N28803), .QN(n7394) );
  DFF_X1 \CACHE_MEM_reg[14][167]  ( .D(n13839), .CK(N28803), .QN(n7410) );
  DFF_X1 \CACHE_MEM_reg[14][166]  ( .D(n13838), .CK(N28803), .QN(n7426) );
  DFF_X1 \CACHE_MEM_reg[14][165]  ( .D(n13837), .CK(N28803), .QN(n7442) );
  DFF_X1 \CACHE_MEM_reg[14][164]  ( .D(n13836), .CK(N28803), .QN(n7458) );
  DFF_X1 \CACHE_MEM_reg[14][163]  ( .D(n13835), .CK(N28803), .QN(n7474) );
  DFF_X1 \CACHE_MEM_reg[14][162]  ( .D(n13834), .CK(N28803), .QN(n7490) );
  DFF_X1 \CACHE_MEM_reg[14][161]  ( .D(n13833), .CK(N28803), .QN(n7506) );
  DFF_X1 \CACHE_MEM_reg[14][160]  ( .D(n13832), .CK(N28803), .QN(n7522) );
  DFF_X1 \CACHE_MEM_reg[14][159]  ( .D(n13831), .CK(N28803), .QN(n7538) );
  DFF_X1 \CACHE_MEM_reg[14][158]  ( .D(n13830), .CK(N28803), .QN(n7554) );
  DFF_X1 \CACHE_MEM_reg[14][157]  ( .D(n13829), .CK(N28803), .QN(n7570) );
  DFF_X1 \CACHE_MEM_reg[14][156]  ( .D(n13828), .CK(N28803), .QN(n7586) );
  DFF_X1 \CACHE_MEM_reg[14][155]  ( .D(n13827), .CK(N28803), .QN(n7602) );
  DFF_X1 \CACHE_MEM_reg[14][154]  ( .D(n13826), .CK(N28803), .QN(n7618) );
  DFF_X1 \CACHE_MEM_reg[14][153]  ( .D(n13825), .CK(N28803), .QN(n7634) );
  DFF_X1 \CACHE_MEM_reg[14][152]  ( .D(n13824), .CK(N28803), .QN(n7650) );
  DFF_X1 \CACHE_MEM_reg[14][151]  ( .D(n13823), .CK(N28803), .QN(n7666) );
  DFF_X1 \CACHE_MEM_reg[14][150]  ( .D(n13822), .CK(N28803), .QN(n7682) );
  DFF_X1 \CACHE_MEM_reg[14][149]  ( .D(n13821), .CK(N28803), .QN(n7698) );
  DFF_X1 \CACHE_MEM_reg[14][148]  ( .D(n13820), .CK(N28803), .QN(n7714) );
  DFF_X1 \CACHE_MEM_reg[14][147]  ( .D(n13819), .CK(N28803), .QN(n7730) );
  DFF_X1 \CACHE_MEM_reg[14][146]  ( .D(n13818), .CK(N28803), .QN(n7746) );
  DFF_X1 \CACHE_MEM_reg[14][145]  ( .D(n13817), .CK(N28803), .QN(n7762) );
  DFF_X1 \CACHE_MEM_reg[14][144]  ( .D(n13816), .CK(N28803), .QN(n7778) );
  DFF_X1 \CACHE_MEM_reg[14][143]  ( .D(n13815), .CK(N28803), .QN(n7794) );
  DFF_X1 \CACHE_MEM_reg[14][142]  ( .D(n13814), .CK(N28803), .QN(n7810) );
  DFF_X1 \CACHE_MEM_reg[14][141]  ( .D(n13813), .CK(N28803), .QN(n7826) );
  DFF_X1 \CACHE_MEM_reg[14][140]  ( .D(n13812), .CK(N28803), .QN(n7842) );
  DFF_X1 \CACHE_MEM_reg[14][139]  ( .D(n13811), .CK(N28803), .QN(n7858) );
  DFF_X1 \CACHE_MEM_reg[14][138]  ( .D(n13810), .CK(N28803), .QN(n7874) );
  DFF_X1 \CACHE_MEM_reg[14][137]  ( .D(n13809), .CK(N28803), .QN(n7890) );
  DFF_X1 \CACHE_MEM_reg[14][136]  ( .D(n13808), .CK(N28803), .QN(n7906) );
  DFF_X1 \CACHE_MEM_reg[14][135]  ( .D(n13807), .CK(N28803), .QN(n7922) );
  DFF_X1 \CACHE_MEM_reg[14][134]  ( .D(n13806), .CK(N28803), .QN(n7938) );
  DFF_X1 \CACHE_MEM_reg[14][133]  ( .D(n13805), .CK(N28803), .QN(n7954) );
  DFF_X1 \CACHE_MEM_reg[14][132]  ( .D(n13804), .CK(N28803), .QN(n7970) );
  DFF_X1 \CACHE_MEM_reg[14][131]  ( .D(n13803), .CK(N28803), .QN(n7986) );
  DFF_X1 \CACHE_MEM_reg[14][130]  ( .D(n13802), .CK(N28803), .QN(n8002) );
  DFF_X1 \CACHE_MEM_reg[14][129]  ( .D(n13801), .CK(N28803), .QN(n8018) );
  DFF_X1 \CACHE_MEM_reg[14][128]  ( .D(n13800), .CK(N28803), .QN(n8034) );
  DFF_X1 \CACHE_MEM_reg[14][127]  ( .D(n13799), .CK(N28803), .QN(n8050) );
  DFF_X1 \CACHE_MEM_reg[14][126]  ( .D(n13798), .CK(N28803), .QN(n8066) );
  DFF_X1 \CACHE_MEM_reg[14][125]  ( .D(n13797), .CK(N28803), .QN(n8082) );
  DFF_X1 \CACHE_MEM_reg[14][124]  ( .D(n13796), .CK(N28803), .QN(n8098) );
  DFF_X1 \CACHE_MEM_reg[14][123]  ( .D(n13795), .CK(N28803), .QN(n8114) );
  DFF_X1 \CACHE_MEM_reg[14][122]  ( .D(n13794), .CK(N28803), .QN(n8130) );
  DFF_X1 \CACHE_MEM_reg[14][121]  ( .D(n13793), .CK(N28803), .QN(n8146) );
  DFF_X1 \CACHE_MEM_reg[14][120]  ( .D(n13792), .CK(N28803), .QN(n8162) );
  DFF_X1 \CACHE_MEM_reg[14][119]  ( .D(n13791), .CK(N28803), .QN(n8178) );
  DFF_X1 \CACHE_MEM_reg[14][118]  ( .D(n13790), .CK(N28803), .QN(n8194) );
  DFF_X1 \CACHE_MEM_reg[14][117]  ( .D(n13789), .CK(N28803), .QN(n8210) );
  DFF_X1 \CACHE_MEM_reg[14][116]  ( .D(n13788), .CK(N28803), .QN(n8226) );
  DFF_X1 \CACHE_MEM_reg[14][115]  ( .D(n13787), .CK(N28803), .QN(n8242) );
  DFF_X1 \CACHE_MEM_reg[14][114]  ( .D(n13786), .CK(N28803), .QN(n8258) );
  DFF_X1 \CACHE_MEM_reg[14][113]  ( .D(n13785), .CK(N28803), .QN(n8274) );
  DFF_X1 \CACHE_MEM_reg[14][112]  ( .D(n13784), .CK(N28803), .QN(n8290) );
  DFF_X1 \CACHE_MEM_reg[14][111]  ( .D(n13783), .CK(N28803), .QN(n8306) );
  DFF_X1 \CACHE_MEM_reg[14][110]  ( .D(n13782), .CK(N28803), .QN(n8322) );
  DFF_X1 \CACHE_MEM_reg[14][109]  ( .D(n13781), .CK(N28803), .QN(n8338) );
  DFF_X1 \CACHE_MEM_reg[14][108]  ( .D(n13780), .CK(N28803), .QN(n8354) );
  DFF_X1 \CACHE_MEM_reg[14][107]  ( .D(n13779), .CK(N28803), .QN(n8370) );
  DFF_X1 \CACHE_MEM_reg[14][106]  ( .D(n13778), .CK(N28803), .QN(n8386) );
  DFF_X1 \CACHE_MEM_reg[14][105]  ( .D(n13777), .CK(N28803), .QN(n8402) );
  DFF_X1 \CACHE_MEM_reg[14][104]  ( .D(n13776), .CK(N28803), .QN(n8418) );
  DFF_X1 \CACHE_MEM_reg[14][103]  ( .D(n13775), .CK(N28803), .QN(n8434) );
  DFF_X1 \CACHE_MEM_reg[14][102]  ( .D(n13774), .CK(N28803), .QN(n8450) );
  DFF_X1 \CACHE_MEM_reg[14][101]  ( .D(n13773), .CK(N28803), .QN(n8466) );
  DFF_X1 \CACHE_MEM_reg[14][100]  ( .D(n13772), .CK(N28803), .QN(n8482) );
  DFF_X1 \CACHE_MEM_reg[14][99]  ( .D(n13771), .CK(N28803), .QN(n8498) );
  DFF_X1 \CACHE_MEM_reg[14][98]  ( .D(n13770), .CK(N28803), .QN(n8514) );
  DFF_X1 \CACHE_MEM_reg[14][97]  ( .D(n13769), .CK(N28803), .QN(n8530) );
  DFF_X1 \CACHE_MEM_reg[14][96]  ( .D(n13768), .CK(N28803), .QN(n8546) );
  DFF_X1 \CACHE_MEM_reg[14][95]  ( .D(n13767), .CK(N28803), .QN(n8562) );
  DFF_X1 \CACHE_MEM_reg[14][94]  ( .D(n13766), .CK(N28803), .QN(n8578) );
  DFF_X1 \CACHE_MEM_reg[14][93]  ( .D(n13765), .CK(N28803), .QN(n8594) );
  DFF_X1 \CACHE_MEM_reg[14][92]  ( .D(n13764), .CK(N28803), .QN(n8610) );
  DFF_X1 \CACHE_MEM_reg[14][91]  ( .D(n13763), .CK(N28803), .QN(n8626) );
  DFF_X1 \CACHE_MEM_reg[14][90]  ( .D(n13762), .CK(N28803), .QN(n8642) );
  DFF_X1 \CACHE_MEM_reg[14][89]  ( .D(n13761), .CK(N28803), .QN(n8658) );
  DFF_X1 \CACHE_MEM_reg[14][88]  ( .D(n13760), .CK(N28803), .QN(n8674) );
  DFF_X1 \CACHE_MEM_reg[14][87]  ( .D(n13759), .CK(N28803), .QN(n8690) );
  DFF_X1 \CACHE_MEM_reg[14][86]  ( .D(n13758), .CK(N28803), .QN(n8706) );
  DFF_X1 \CACHE_MEM_reg[14][85]  ( .D(n13757), .CK(N28803), .QN(n8722) );
  DFF_X1 \CACHE_MEM_reg[14][84]  ( .D(n13756), .CK(N28803), .QN(n8738) );
  DFF_X1 \CACHE_MEM_reg[14][83]  ( .D(n13755), .CK(N28803), .QN(n8754) );
  DFF_X1 \CACHE_MEM_reg[14][82]  ( .D(n13754), .CK(N28803), .QN(n8770) );
  DFF_X1 \CACHE_MEM_reg[14][81]  ( .D(n13753), .CK(N28803), .QN(n8786) );
  DFF_X1 \CACHE_MEM_reg[14][80]  ( .D(n13752), .CK(N28803), .QN(n8802) );
  DFF_X1 \CACHE_MEM_reg[14][79]  ( .D(n13751), .CK(N28803), .QN(n8818) );
  DFF_X1 \CACHE_MEM_reg[14][78]  ( .D(n13750), .CK(N28803), .QN(n8834) );
  DFF_X1 \CACHE_MEM_reg[14][77]  ( .D(n13749), .CK(N28803), .QN(n8850) );
  DFF_X1 \CACHE_MEM_reg[14][76]  ( .D(n13748), .CK(N28803), .QN(n8866) );
  DFF_X1 \CACHE_MEM_reg[14][75]  ( .D(n13747), .CK(N28803), .QN(n8882) );
  DFF_X1 \CACHE_MEM_reg[14][74]  ( .D(n13746), .CK(N28803), .QN(n8898) );
  DFF_X1 \CACHE_MEM_reg[14][73]  ( .D(n13745), .CK(N28803), .QN(n8914) );
  DFF_X1 \CACHE_MEM_reg[14][72]  ( .D(n13744), .CK(N28803), .QN(n8930) );
  DFF_X1 \CACHE_MEM_reg[14][71]  ( .D(n13743), .CK(N28803), .QN(n8946) );
  DFF_X1 \CACHE_MEM_reg[14][70]  ( .D(n13742), .CK(N28803), .QN(n8962) );
  DFF_X1 \CACHE_MEM_reg[14][69]  ( .D(n13741), .CK(N28803), .QN(n8978) );
  DFF_X1 \CACHE_MEM_reg[14][68]  ( .D(n13740), .CK(N28803), .QN(n8994) );
  DFF_X1 \CACHE_MEM_reg[14][67]  ( .D(n13739), .CK(N28803), .QN(n9010) );
  DFF_X1 \CACHE_MEM_reg[14][66]  ( .D(n13738), .CK(N28803), .QN(n9026) );
  DFF_X1 \CACHE_MEM_reg[14][65]  ( .D(n13737), .CK(N28803), .QN(n9042) );
  DFF_X1 \CACHE_MEM_reg[14][64]  ( .D(n13736), .CK(N28803), .QN(n9058) );
  DFF_X1 \CACHE_MEM_reg[14][63]  ( .D(n13735), .CK(N28803), .QN(n9074) );
  DFF_X1 \CACHE_MEM_reg[14][62]  ( .D(n13734), .CK(N28803), .QN(n9090) );
  DFF_X1 \CACHE_MEM_reg[14][61]  ( .D(n13733), .CK(N28803), .QN(n9106) );
  DFF_X1 \CACHE_MEM_reg[14][60]  ( .D(n13732), .CK(N28803), .QN(n9122) );
  DFF_X1 \CACHE_MEM_reg[14][59]  ( .D(n13731), .CK(N28803), .QN(n9138) );
  DFF_X1 \CACHE_MEM_reg[14][58]  ( .D(n13730), .CK(N28803), .QN(n9154) );
  DFF_X1 \CACHE_MEM_reg[14][57]  ( .D(n13729), .CK(N28803), .QN(n9170) );
  DFF_X1 \CACHE_MEM_reg[14][56]  ( .D(n13728), .CK(N28803), .QN(n9186) );
  DFF_X1 \CACHE_MEM_reg[14][55]  ( .D(n13727), .CK(N28803), .QN(n9202) );
  DFF_X1 \CACHE_MEM_reg[14][54]  ( .D(n13726), .CK(N28803), .QN(n9218) );
  DFF_X1 \CACHE_MEM_reg[14][53]  ( .D(n13725), .CK(N28803), .QN(n9234) );
  DFF_X1 \CACHE_MEM_reg[14][52]  ( .D(n13724), .CK(N28803), .QN(n9250) );
  DFF_X1 \CACHE_MEM_reg[14][51]  ( .D(n13723), .CK(N28803), .QN(n9266) );
  DFF_X1 \CACHE_MEM_reg[14][50]  ( .D(n13722), .CK(N28803), .QN(n9282) );
  DFF_X1 \CACHE_MEM_reg[14][49]  ( .D(n13721), .CK(N28803), .QN(n9298) );
  DFF_X1 \CACHE_MEM_reg[14][48]  ( .D(n13720), .CK(N28803), .QN(n9314) );
  DFF_X1 \CACHE_MEM_reg[14][47]  ( .D(n13719), .CK(N28803), .QN(n9330) );
  DFF_X1 \CACHE_MEM_reg[14][46]  ( .D(n13718), .CK(N28803), .QN(n9346) );
  DFF_X1 \CACHE_MEM_reg[14][45]  ( .D(n13717), .CK(N28803), .QN(n9362) );
  DFF_X1 \CACHE_MEM_reg[14][44]  ( .D(n13716), .CK(N28803), .QN(n9378) );
  DFF_X1 \CACHE_MEM_reg[14][43]  ( .D(n13715), .CK(N28803), .QN(n9394) );
  DFF_X1 \CACHE_MEM_reg[14][42]  ( .D(n13714), .CK(N28803), .QN(n9410) );
  DFF_X1 \CACHE_MEM_reg[14][41]  ( .D(n13713), .CK(N28803), .QN(n9426) );
  DFF_X1 \CACHE_MEM_reg[14][40]  ( .D(n13712), .CK(N28803), .QN(n9442) );
  DFF_X1 \CACHE_MEM_reg[14][39]  ( .D(n13711), .CK(N28803), .QN(n9458) );
  DFF_X1 \CACHE_MEM_reg[14][38]  ( .D(n13710), .CK(N28803), .QN(n9474) );
  DFF_X1 \CACHE_MEM_reg[14][37]  ( .D(n13709), .CK(N28803), .QN(n9490) );
  DFF_X1 \CACHE_MEM_reg[14][36]  ( .D(n13708), .CK(N28803), .QN(n9506) );
  DFF_X1 \CACHE_MEM_reg[14][35]  ( .D(n13707), .CK(N28803), .QN(n9522) );
  DFF_X1 \CACHE_MEM_reg[14][34]  ( .D(n13706), .CK(N28803), .QN(n9538) );
  DFF_X1 \CACHE_MEM_reg[14][33]  ( .D(n13705), .CK(N28803), .QN(n9554) );
  DFF_X1 \CACHE_MEM_reg[14][32]  ( .D(n13704), .CK(N28803), .QN(n9570) );
  DFF_X1 \CACHE_MEM_reg[14][31]  ( .D(n13703), .CK(N28803), .QN(n9586) );
  DFF_X1 \CACHE_MEM_reg[14][30]  ( .D(n13702), .CK(N28803), .QN(n9602) );
  DFF_X1 \CACHE_MEM_reg[14][29]  ( .D(n13701), .CK(N28803), .QN(n9618) );
  DFF_X1 \CACHE_MEM_reg[14][28]  ( .D(n13700), .CK(N28803), .QN(n9634) );
  DFF_X1 \CACHE_MEM_reg[14][27]  ( .D(n13699), .CK(N28803), .QN(n9650) );
  DFF_X1 \CACHE_MEM_reg[14][26]  ( .D(n13698), .CK(N28803), .QN(n9666) );
  DFF_X1 \CACHE_MEM_reg[14][25]  ( .D(n13697), .CK(N28803), .QN(n9682) );
  DFF_X1 \CACHE_MEM_reg[14][24]  ( .D(n13696), .CK(N28803), .QN(n9698) );
  DFF_X1 \CACHE_MEM_reg[14][23]  ( .D(n13695), .CK(N28803), .QN(n9714) );
  DFF_X1 \CACHE_MEM_reg[14][22]  ( .D(n13694), .CK(N28803), .QN(n9730) );
  DFF_X1 \CACHE_MEM_reg[14][21]  ( .D(n13693), .CK(N28803), .QN(n9746) );
  DFF_X1 \CACHE_MEM_reg[14][20]  ( .D(n13692), .CK(N28803), .QN(n9762) );
  DFF_X1 \CACHE_MEM_reg[14][19]  ( .D(n13691), .CK(N28803), .QN(n9778) );
  DFF_X1 \CACHE_MEM_reg[14][18]  ( .D(n13690), .CK(N28803), .QN(n9794) );
  DFF_X1 \CACHE_MEM_reg[14][17]  ( .D(n13689), .CK(N28803), .QN(n9810) );
  DFF_X1 \CACHE_MEM_reg[14][16]  ( .D(n13688), .CK(N28803), .QN(n9826) );
  DFF_X1 \CACHE_MEM_reg[14][15]  ( .D(n13687), .CK(N28803), .QN(n9842) );
  DFF_X1 \CACHE_MEM_reg[14][14]  ( .D(n13686), .CK(N28803), .QN(n9858) );
  DFF_X1 \CACHE_MEM_reg[14][13]  ( .D(n13685), .CK(N28803), .QN(n9874) );
  DFF_X1 \CACHE_MEM_reg[14][12]  ( .D(n13684), .CK(N28803), .QN(n9890) );
  DFF_X1 \CACHE_MEM_reg[14][11]  ( .D(n13683), .CK(N28803), .QN(n9906) );
  DFF_X1 \CACHE_MEM_reg[14][10]  ( .D(n13682), .CK(N28803), .QN(n9922) );
  DFF_X1 \CACHE_MEM_reg[14][9]  ( .D(n13681), .CK(N28803), .QN(n9938) );
  DFF_X1 \CACHE_MEM_reg[14][8]  ( .D(n13680), .CK(N28803), .QN(n9954) );
  DFF_X1 \CACHE_MEM_reg[14][7]  ( .D(n13679), .CK(N28803), .QN(n9970) );
  DFF_X1 \CACHE_MEM_reg[14][6]  ( .D(n13678), .CK(N28803), .QN(n9986) );
  DFF_X1 \CACHE_MEM_reg[14][5]  ( .D(n13677), .CK(N28803), .QN(n10002) );
  DFF_X1 \CACHE_MEM_reg[14][4]  ( .D(n13676), .CK(N28803), .QN(n10018) );
  DFF_X1 \CACHE_MEM_reg[14][3]  ( .D(n13675), .CK(N28803), .QN(n10034) );
  DFF_X1 \CACHE_MEM_reg[14][2]  ( .D(n13674), .CK(N28803), .QN(n10050) );
  DFF_X1 \CACHE_MEM_reg[14][1]  ( .D(n13673), .CK(N28803), .QN(n10066) );
  DFF_X1 \CACHE_MEM_reg[14][0]  ( .D(n13672), .CK(N28803), .QN(n10082) );
  DFF_X1 \CACHE_MEM_reg[13][255]  ( .D(n13671), .CK(N28803), .Q(n3563), .QN(
        n5998) );
  DFF_X1 \CACHE_MEM_reg[13][254]  ( .D(n13670), .CK(N28803), .Q(n3555), .QN(
        n6014) );
  DFF_X1 \CACHE_MEM_reg[13][253]  ( .D(n13669), .CK(N28803), .Q(n3548), .QN(
        n6030) );
  DFF_X1 \CACHE_MEM_reg[13][252]  ( .D(n13668), .CK(N28803), .Q(n3542), .QN(
        n6046) );
  DFF_X1 \CACHE_MEM_reg[13][251]  ( .D(n13667), .CK(N28803), .Q(n3531), .QN(
        n6062) );
  DFF_X1 \CACHE_MEM_reg[13][250]  ( .D(n13666), .CK(N28803), .Q(n3527), .QN(
        n6078) );
  DFF_X1 \CACHE_MEM_reg[13][249]  ( .D(n13665), .CK(N28803), .Q(n3520), .QN(
        n6094) );
  DFF_X1 \CACHE_MEM_reg[13][248]  ( .D(n13664), .CK(N28803), .Q(n3514), .QN(
        n6110) );
  DFF_X1 \CACHE_MEM_reg[13][247]  ( .D(n13663), .CK(N28803), .Q(n3507), .QN(
        n6126) );
  DFF_X1 \CACHE_MEM_reg[13][246]  ( .D(n13662), .CK(N28803), .Q(n3503), .QN(
        n6142) );
  DFF_X1 \CACHE_MEM_reg[13][245]  ( .D(n13661), .CK(N28803), .Q(n3492), .QN(
        n6158) );
  DFF_X1 \CACHE_MEM_reg[13][244]  ( .D(n13660), .CK(N28803), .Q(n3486), .QN(
        n6174) );
  DFF_X1 \CACHE_MEM_reg[13][243]  ( .D(n13659), .CK(N28803), .Q(n3479), .QN(
        n6190) );
  DFF_X1 \CACHE_MEM_reg[13][242]  ( .D(n13658), .CK(N28803), .Q(n3475), .QN(
        n6206) );
  DFF_X1 \CACHE_MEM_reg[13][241]  ( .D(n13657), .CK(N28803), .Q(n3468), .QN(
        n6222) );
  DFF_X1 \CACHE_MEM_reg[13][240]  ( .D(n13656), .CK(N28803), .Q(n3458), .QN(
        n6238) );
  DFF_X1 \CACHE_MEM_reg[13][239]  ( .D(n13655), .CK(N28803), .Q(n3451), .QN(
        n6254) );
  DFF_X1 \CACHE_MEM_reg[13][238]  ( .D(n13654), .CK(N28803), .Q(n3447), .QN(
        n6270) );
  DFF_X1 \CACHE_MEM_reg[13][237]  ( .D(n13653), .CK(N28803), .Q(n3440), .QN(
        n6286) );
  DFF_X1 \CACHE_MEM_reg[13][236]  ( .D(n13652), .CK(N28803), .Q(n3434), .QN(
        n6302) );
  DFF_X1 \CACHE_MEM_reg[13][235]  ( .D(n13651), .CK(N28803), .Q(n3418), .QN(
        n6318) );
  DFF_X1 \CACHE_MEM_reg[13][234]  ( .D(n13650), .CK(N28803), .Q(n3414), .QN(
        n6334) );
  DFF_X1 \CACHE_MEM_reg[13][233]  ( .D(n13649), .CK(N28803), .Q(n3407), .QN(
        n6350) );
  DFF_X1 \CACHE_MEM_reg[13][232]  ( .D(n13648), .CK(N28803), .Q(n3401), .QN(
        n6366) );
  DFF_X1 \CACHE_MEM_reg[13][231]  ( .D(n13647), .CK(N28803), .Q(n3394), .QN(
        n6382) );
  DFF_X1 \CACHE_MEM_reg[13][230]  ( .D(n13646), .CK(N28803), .Q(n3390), .QN(
        n6398) );
  DFF_X1 \CACHE_MEM_reg[13][229]  ( .D(n13645), .CK(N28803), .Q(n3379), .QN(
        n6414) );
  DFF_X1 \CACHE_MEM_reg[13][228]  ( .D(n13644), .CK(N28803), .Q(n3373), .QN(
        n6430) );
  DFF_X1 \CACHE_MEM_reg[13][227]  ( .D(n13643), .CK(N28803), .Q(n3366), .QN(
        n6446) );
  DFF_X1 \CACHE_MEM_reg[13][226]  ( .D(n13642), .CK(N28803), .Q(n3362), .QN(
        n6462) );
  DFF_X1 \CACHE_MEM_reg[13][225]  ( .D(n13641), .CK(N28803), .Q(n3355), .QN(
        n6478) );
  DFF_X1 \CACHE_MEM_reg[13][224]  ( .D(n13640), .CK(N28803), .Q(n3345), .QN(
        n6494) );
  DFF_X1 \CACHE_MEM_reg[13][223]  ( .D(n13639), .CK(N28803), .Q(n5263), .QN(
        n6510) );
  DFF_X1 \CACHE_MEM_reg[13][222]  ( .D(n13638), .CK(N28803), .Q(n5246), .QN(
        n6526) );
  DFF_X1 \CACHE_MEM_reg[13][221]  ( .D(n13637), .CK(N28803), .Q(n5235), .QN(
        n6542) );
  DFF_X1 \CACHE_MEM_reg[13][220]  ( .D(n13636), .CK(N28803), .Q(n5222), .QN(
        n6558) );
  DFF_X1 \CACHE_MEM_reg[13][219]  ( .D(n13635), .CK(N28803), .Q(n5202), .QN(
        n6574) );
  DFF_X1 \CACHE_MEM_reg[13][218]  ( .D(n13634), .CK(N28803), .Q(n5189), .QN(
        n6590) );
  DFF_X1 \CACHE_MEM_reg[13][217]  ( .D(n13633), .CK(N28803), .Q(n5178), .QN(
        n6606) );
  DFF_X1 \CACHE_MEM_reg[13][216]  ( .D(n13632), .CK(N28803), .Q(n5161), .QN(
        n6622) );
  DFF_X1 \CACHE_MEM_reg[13][215]  ( .D(n13631), .CK(N28803), .Q(n5150), .QN(
        n6638) );
  DFF_X1 \CACHE_MEM_reg[13][214]  ( .D(n13630), .CK(N28803), .Q(n5133), .QN(
        n6654) );
  DFF_X1 \CACHE_MEM_reg[13][213]  ( .D(n13629), .CK(N28803), .Q(n5122), .QN(
        n6670) );
  DFF_X1 \CACHE_MEM_reg[13][212]  ( .D(n13628), .CK(N28803), .Q(n5109), .QN(
        n6686) );
  DFF_X1 \CACHE_MEM_reg[13][211]  ( .D(n13627), .CK(N28803), .Q(n5094), .QN(
        n6702) );
  DFF_X1 \CACHE_MEM_reg[13][210]  ( .D(n13626), .CK(N28803), .Q(n5081), .QN(
        n6718) );
  DFF_X1 \CACHE_MEM_reg[13][209]  ( .D(n13625), .CK(N28803), .Q(n5070), .QN(
        n6734) );
  DFF_X1 \CACHE_MEM_reg[13][208]  ( .D(n13624), .CK(N28803), .Q(n5053), .QN(
        n6750) );
  DFF_X1 \CACHE_MEM_reg[13][207]  ( .D(n13623), .CK(N28803), .Q(n5040), .QN(
        n6766) );
  DFF_X1 \CACHE_MEM_reg[13][206]  ( .D(n13622), .CK(N28803), .Q(n5029), .QN(
        n6782) );
  DFF_X1 \CACHE_MEM_reg[13][205]  ( .D(n13621), .CK(N28803), .Q(n5012), .QN(
        n6798) );
  DFF_X1 \CACHE_MEM_reg[13][204]  ( .D(n13620), .CK(N28803), .Q(n5001), .QN(
        n6814) );
  DFF_X1 \CACHE_MEM_reg[13][203]  ( .D(n13619), .CK(N28803), .Q(n4984), .QN(
        n6830) );
  DFF_X1 \CACHE_MEM_reg[13][202]  ( .D(n13618), .CK(N28803), .Q(n4973), .QN(
        n6846) );
  DFF_X1 \CACHE_MEM_reg[13][201]  ( .D(n13617), .CK(N28803), .Q(n4960), .QN(
        n6862) );
  DFF_X1 \CACHE_MEM_reg[13][200]  ( .D(n13616), .CK(N28803), .Q(n4945), .QN(
        n6878) );
  DFF_X1 \CACHE_MEM_reg[13][199]  ( .D(n13615), .CK(N28803), .Q(n4932), .QN(
        n6894) );
  DFF_X1 \CACHE_MEM_reg[13][198]  ( .D(n13614), .CK(N28803), .Q(n4921), .QN(
        n6910) );
  DFF_X1 \CACHE_MEM_reg[13][197]  ( .D(n13613), .CK(N28803), .Q(n4899), .QN(
        n6926) );
  DFF_X1 \CACHE_MEM_reg[13][196]  ( .D(n13612), .CK(N28803), .Q(n4888), .QN(
        n6942) );
  DFF_X1 \CACHE_MEM_reg[13][195]  ( .D(n13611), .CK(N28803), .Q(n4871), .QN(
        n6958) );
  DFF_X1 \CACHE_MEM_reg[13][194]  ( .D(n13610), .CK(N28803), .Q(n4860), .QN(
        n6974) );
  DFF_X1 \CACHE_MEM_reg[13][193]  ( .D(n13609), .CK(N28803), .Q(n4847), .QN(
        n6990) );
  DFF_X1 \CACHE_MEM_reg[13][192]  ( .D(n13608), .CK(N28803), .Q(n4832), .QN(
        n7006) );
  DFF_X1 \CACHE_MEM_reg[13][191]  ( .D(n13607), .CK(N28803), .Q(n5705), .QN(
        n7022) );
  DFF_X1 \CACHE_MEM_reg[13][190]  ( .D(n13606), .CK(N28803), .Q(n3556), .QN(
        n7038) );
  DFF_X1 \CACHE_MEM_reg[13][189]  ( .D(n13605), .CK(N28803), .Q(n3550), .QN(
        n7054) );
  DFF_X1 \CACHE_MEM_reg[13][188]  ( .D(n13604), .CK(N28803), .Q(n3543), .QN(
        n7070) );
  DFF_X1 \CACHE_MEM_reg[13][187]  ( .D(n13603), .CK(N28803), .Q(n3539), .QN(
        n7086) );
  DFF_X1 \CACHE_MEM_reg[13][186]  ( .D(n13602), .CK(N28803), .Q(n3528), .QN(
        n7102) );
  DFF_X1 \CACHE_MEM_reg[13][185]  ( .D(n13601), .CK(N28803), .Q(n3522), .QN(
        n7118) );
  DFF_X1 \CACHE_MEM_reg[13][184]  ( .D(n13600), .CK(N28803), .Q(n3515), .QN(
        n7134) );
  DFF_X1 \CACHE_MEM_reg[13][183]  ( .D(n13599), .CK(N28803), .Q(n3511), .QN(
        n7150) );
  DFF_X1 \CACHE_MEM_reg[13][182]  ( .D(n13598), .CK(N28803), .Q(n3504), .QN(
        n7166) );
  DFF_X1 \CACHE_MEM_reg[13][181]  ( .D(n13597), .CK(N28803), .Q(n3494), .QN(
        n7182) );
  DFF_X1 \CACHE_MEM_reg[13][180]  ( .D(n13596), .CK(N28803), .Q(n3487), .QN(
        n7198) );
  DFF_X1 \CACHE_MEM_reg[13][179]  ( .D(n13595), .CK(N28803), .Q(n3483), .QN(
        n7214) );
  DFF_X1 \CACHE_MEM_reg[13][178]  ( .D(n13594), .CK(N28803), .Q(n3476), .QN(
        n7230) );
  DFF_X1 \CACHE_MEM_reg[13][177]  ( .D(n13593), .CK(N28803), .Q(n3470), .QN(
        n7246) );
  DFF_X1 \CACHE_MEM_reg[13][176]  ( .D(n13592), .CK(N28803), .Q(n3459), .QN(
        n7262) );
  DFF_X1 \CACHE_MEM_reg[13][175]  ( .D(n13591), .CK(N28803), .Q(n3455), .QN(
        n7278) );
  DFF_X1 \CACHE_MEM_reg[13][174]  ( .D(n13590), .CK(N28803), .Q(n3448), .QN(
        n7294) );
  DFF_X1 \CACHE_MEM_reg[13][173]  ( .D(n13589), .CK(N28803), .Q(n3442), .QN(
        n7310) );
  DFF_X1 \CACHE_MEM_reg[13][172]  ( .D(n13588), .CK(N28803), .Q(n3435), .QN(
        n7326) );
  DFF_X1 \CACHE_MEM_reg[13][171]  ( .D(n13587), .CK(N28803), .Q(n3431), .QN(
        n7342) );
  DFF_X1 \CACHE_MEM_reg[13][170]  ( .D(n13586), .CK(N28803), .Q(n3415), .QN(
        n7358) );
  DFF_X1 \CACHE_MEM_reg[13][169]  ( .D(n13585), .CK(N28803), .Q(n3409), .QN(
        n7374) );
  DFF_X1 \CACHE_MEM_reg[13][168]  ( .D(n13584), .CK(N28803), .Q(n3402), .QN(
        n7390) );
  DFF_X1 \CACHE_MEM_reg[13][167]  ( .D(n13583), .CK(N28803), .Q(n3398), .QN(
        n7406) );
  DFF_X1 \CACHE_MEM_reg[13][166]  ( .D(n13582), .CK(N28803), .Q(n3391), .QN(
        n7422) );
  DFF_X1 \CACHE_MEM_reg[13][165]  ( .D(n13581), .CK(N28803), .Q(n3381), .QN(
        n7438) );
  DFF_X1 \CACHE_MEM_reg[13][164]  ( .D(n13580), .CK(N28803), .Q(n3374), .QN(
        n7454) );
  DFF_X1 \CACHE_MEM_reg[13][163]  ( .D(n13579), .CK(N28803), .Q(n3370), .QN(
        n7470) );
  DFF_X1 \CACHE_MEM_reg[13][162]  ( .D(n13578), .CK(N28803), .Q(n3363), .QN(
        n7486) );
  DFF_X1 \CACHE_MEM_reg[13][161]  ( .D(n13577), .CK(N28803), .Q(n3357), .QN(
        n7502) );
  DFF_X1 \CACHE_MEM_reg[13][160]  ( .D(n13576), .CK(N28803), .Q(n3346), .QN(
        n7518) );
  DFF_X1 \CACHE_MEM_reg[13][159]  ( .D(n13575), .CK(N28803), .Q(n5710), .QN(
        n7534) );
  DFF_X1 \CACHE_MEM_reg[13][158]  ( .D(n13574), .CK(N28803), .Q(n5693), .QN(
        n7550) );
  DFF_X1 \CACHE_MEM_reg[13][157]  ( .D(n13573), .CK(N28803), .Q(n5682), .QN(
        n7566) );
  DFF_X1 \CACHE_MEM_reg[13][156]  ( .D(n13572), .CK(N28803), .Q(n5669), .QN(
        n7582) );
  DFF_X1 \CACHE_MEM_reg[13][155]  ( .D(n13571), .CK(N28803), .Q(n5649), .QN(
        n7598) );
  DFF_X1 \CACHE_MEM_reg[13][154]  ( .D(n13570), .CK(N28803), .Q(n5636), .QN(
        n7614) );
  DFF_X1 \CACHE_MEM_reg[13][153]  ( .D(n13569), .CK(N28803), .Q(n5625), .QN(
        n7630) );
  DFF_X1 \CACHE_MEM_reg[13][152]  ( .D(n13568), .CK(N28803), .Q(n5608), .QN(
        n7646) );
  DFF_X1 \CACHE_MEM_reg[13][151]  ( .D(n13567), .CK(N28803), .Q(n5597), .QN(
        n7662) );
  DFF_X1 \CACHE_MEM_reg[13][150]  ( .D(n13566), .CK(N28803), .Q(n5580), .QN(
        n7678) );
  DFF_X1 \CACHE_MEM_reg[13][149]  ( .D(n13565), .CK(N28803), .Q(n5569), .QN(
        n7694) );
  DFF_X1 \CACHE_MEM_reg[13][148]  ( .D(n13564), .CK(N28803), .Q(n5556), .QN(
        n7710) );
  DFF_X1 \CACHE_MEM_reg[13][147]  ( .D(n13563), .CK(N28803), .Q(n5541), .QN(
        n7726) );
  DFF_X1 \CACHE_MEM_reg[13][146]  ( .D(n13562), .CK(N28803), .Q(n5528), .QN(
        n7742) );
  DFF_X1 \CACHE_MEM_reg[13][145]  ( .D(n13561), .CK(N28803), .Q(n5517), .QN(
        n7758) );
  DFF_X1 \CACHE_MEM_reg[13][144]  ( .D(n13560), .CK(N28803), .Q(n5495), .QN(
        n7774) );
  DFF_X1 \CACHE_MEM_reg[13][143]  ( .D(n13559), .CK(N28803), .Q(n5484), .QN(
        n7790) );
  DFF_X1 \CACHE_MEM_reg[13][142]  ( .D(n13558), .CK(N28803), .Q(n5467), .QN(
        n7806) );
  DFF_X1 \CACHE_MEM_reg[13][141]  ( .D(n13557), .CK(N28803), .Q(n5456), .QN(
        n7822) );
  DFF_X1 \CACHE_MEM_reg[13][140]  ( .D(n13556), .CK(N28803), .Q(n5443), .QN(
        n7838) );
  DFF_X1 \CACHE_MEM_reg[13][139]  ( .D(n13555), .CK(N28803), .Q(n5428), .QN(
        n7854) );
  DFF_X1 \CACHE_MEM_reg[13][138]  ( .D(n13554), .CK(N28803), .Q(n5415), .QN(
        n7870) );
  DFF_X1 \CACHE_MEM_reg[13][137]  ( .D(n13553), .CK(N28803), .Q(n5404), .QN(
        n7886) );
  DFF_X1 \CACHE_MEM_reg[13][136]  ( .D(n13552), .CK(N28803), .Q(n5387), .QN(
        n7902) );
  DFF_X1 \CACHE_MEM_reg[13][135]  ( .D(n13551), .CK(N28803), .Q(n5376), .QN(
        n7918) );
  DFF_X1 \CACHE_MEM_reg[13][134]  ( .D(n13550), .CK(N28803), .Q(n5354), .QN(
        n7934) );
  DFF_X1 \CACHE_MEM_reg[13][133]  ( .D(n13549), .CK(N28803), .Q(n5343), .QN(
        n7950) );
  DFF_X1 \CACHE_MEM_reg[13][132]  ( .D(n13548), .CK(N28803), .Q(n5330), .QN(
        n7966) );
  DFF_X1 \CACHE_MEM_reg[13][131]  ( .D(n13547), .CK(N28803), .Q(n5315), .QN(
        n7982) );
  DFF_X1 \CACHE_MEM_reg[13][130]  ( .D(n13546), .CK(N28803), .Q(n5302), .QN(
        n7998) );
  DFF_X1 \CACHE_MEM_reg[13][129]  ( .D(n13545), .CK(N28803), .Q(n5291), .QN(
        n8014) );
  DFF_X1 \CACHE_MEM_reg[13][128]  ( .D(n13544), .CK(N28803), .Q(n5274), .QN(
        n8030) );
  DFF_X1 \CACHE_MEM_reg[13][127]  ( .D(n13543), .CK(N28803), .Q(n3558), .QN(
        n8046) );
  DFF_X1 \CACHE_MEM_reg[13][126]  ( .D(n13542), .CK(N28803), .Q(n4352), .QN(
        n8062) );
  DFF_X1 \CACHE_MEM_reg[13][125]  ( .D(n13541), .CK(N28803), .Q(n4336), .QN(
        n8078) );
  DFF_X1 \CACHE_MEM_reg[13][124]  ( .D(n13540), .CK(N28803), .Q(n4311), .QN(
        n8094) );
  DFF_X1 \CACHE_MEM_reg[13][123]  ( .D(n13539), .CK(N28803), .Q(n4295), .QN(
        n8110) );
  DFF_X1 \CACHE_MEM_reg[13][122]  ( .D(n13538), .CK(N28803), .Q(n4275), .QN(
        n8126) );
  DFF_X1 \CACHE_MEM_reg[13][121]  ( .D(n13537), .CK(N28803), .Q(n4259), .QN(
        n8142) );
  DFF_X1 \CACHE_MEM_reg[13][120]  ( .D(n13536), .CK(N28803), .Q(n4239), .QN(
        n8158) );
  DFF_X1 \CACHE_MEM_reg[13][119]  ( .D(n13535), .CK(N28803), .Q(n4223), .QN(
        n8174) );
  DFF_X1 \CACHE_MEM_reg[13][118]  ( .D(n13534), .CK(N28803), .Q(n4203), .QN(
        n8190) );
  DFF_X1 \CACHE_MEM_reg[13][117]  ( .D(n13533), .CK(N28803), .Q(n4187), .QN(
        n8206) );
  DFF_X1 \CACHE_MEM_reg[13][116]  ( .D(n13532), .CK(N28803), .Q(n4162), .QN(
        n8222) );
  DFF_X1 \CACHE_MEM_reg[13][115]  ( .D(n13531), .CK(N28803), .Q(n4146), .QN(
        n8238) );
  DFF_X1 \CACHE_MEM_reg[13][114]  ( .D(n13530), .CK(N28803), .Q(n4126), .QN(
        n8254) );
  DFF_X1 \CACHE_MEM_reg[13][113]  ( .D(n13529), .CK(N28803), .Q(n4110), .QN(
        n8270) );
  DFF_X1 \CACHE_MEM_reg[13][112]  ( .D(n13528), .CK(N28803), .Q(n4090), .QN(
        n8286) );
  DFF_X1 \CACHE_MEM_reg[13][111]  ( .D(n13527), .CK(N28803), .Q(n4074), .QN(
        n8302) );
  DFF_X1 \CACHE_MEM_reg[13][110]  ( .D(n13526), .CK(N28803), .Q(n4054), .QN(
        n8318) );
  DFF_X1 \CACHE_MEM_reg[13][109]  ( .D(n13525), .CK(N28803), .Q(n4038), .QN(
        n8334) );
  DFF_X1 \CACHE_MEM_reg[13][108]  ( .D(n13524), .CK(N28803), .Q(n4013), .QN(
        n8350) );
  DFF_X1 \CACHE_MEM_reg[13][107]  ( .D(n13523), .CK(N28803), .Q(n3997), .QN(
        n8366) );
  DFF_X1 \CACHE_MEM_reg[13][106]  ( .D(n13522), .CK(N28803), .Q(n3977), .QN(
        n8382) );
  DFF_X1 \CACHE_MEM_reg[13][105]  ( .D(n13521), .CK(N28803), .Q(n3961), .QN(
        n8398) );
  DFF_X1 \CACHE_MEM_reg[13][104]  ( .D(n13520), .CK(N28803), .Q(n3941), .QN(
        n8414) );
  DFF_X1 \CACHE_MEM_reg[13][103]  ( .D(n13519), .CK(N28803), .Q(n3925), .QN(
        n8430) );
  DFF_X1 \CACHE_MEM_reg[13][102]  ( .D(n13518), .CK(N28803), .Q(n3905), .QN(
        n8446) );
  DFF_X1 \CACHE_MEM_reg[13][101]  ( .D(n13517), .CK(N28803), .Q(n3889), .QN(
        n8462) );
  DFF_X1 \CACHE_MEM_reg[13][100]  ( .D(n13516), .CK(N28803), .Q(n3864), .QN(
        n8478) );
  DFF_X1 \CACHE_MEM_reg[13][99]  ( .D(n13515), .CK(N28803), .Q(n3848), .QN(
        n8494) );
  DFF_X1 \CACHE_MEM_reg[13][98]  ( .D(n13514), .CK(N28803), .Q(n3828), .QN(
        n8510) );
  DFF_X1 \CACHE_MEM_reg[13][97]  ( .D(n13513), .CK(N28803), .Q(n3812), .QN(
        n8526) );
  DFF_X1 \CACHE_MEM_reg[13][96]  ( .D(n13512), .CK(N28803), .Q(n3792), .QN(
        n8542) );
  DFF_X1 \CACHE_MEM_reg[13][95]  ( .D(n13511), .CK(N28803), .Q(n4372), .QN(
        n8558) );
  DFF_X1 \CACHE_MEM_reg[13][94]  ( .D(n13510), .CK(N28803), .Q(n4361), .QN(
        n8574) );
  DFF_X1 \CACHE_MEM_reg[13][93]  ( .D(n13509), .CK(N28803), .Q(n4341), .QN(
        n8590) );
  DFF_X1 \CACHE_MEM_reg[13][92]  ( .D(n13508), .CK(N28803), .Q(n4325), .QN(
        n8606) );
  DFF_X1 \CACHE_MEM_reg[13][91]  ( .D(n13507), .CK(N28803), .Q(n4300), .QN(
        n8622) );
  DFF_X1 \CACHE_MEM_reg[13][90]  ( .D(n13506), .CK(N28803), .Q(n4284), .QN(
        n8638) );
  DFF_X1 \CACHE_MEM_reg[13][89]  ( .D(n13505), .CK(N28803), .Q(n4264), .QN(
        n8654) );
  DFF_X1 \CACHE_MEM_reg[13][88]  ( .D(n13504), .CK(N28803), .Q(n4248), .QN(
        n8670) );
  DFF_X1 \CACHE_MEM_reg[13][87]  ( .D(n13503), .CK(N28803), .Q(n4228), .QN(
        n8686) );
  DFF_X1 \CACHE_MEM_reg[13][86]  ( .D(n13502), .CK(N28803), .Q(n4212), .QN(
        n8702) );
  DFF_X1 \CACHE_MEM_reg[13][85]  ( .D(n13501), .CK(N28803), .Q(n4192), .QN(
        n8718) );
  DFF_X1 \CACHE_MEM_reg[13][84]  ( .D(n13500), .CK(N28803), .Q(n4176), .QN(
        n8734) );
  DFF_X1 \CACHE_MEM_reg[13][83]  ( .D(n13499), .CK(N28803), .Q(n4151), .QN(
        n8750) );
  DFF_X1 \CACHE_MEM_reg[13][82]  ( .D(n13498), .CK(N28803), .Q(n4135), .QN(
        n8766) );
  DFF_X1 \CACHE_MEM_reg[13][81]  ( .D(n13497), .CK(N28803), .Q(n4115), .QN(
        n8782) );
  DFF_X1 \CACHE_MEM_reg[13][80]  ( .D(n13496), .CK(N28803), .Q(n4099), .QN(
        n8798) );
  DFF_X1 \CACHE_MEM_reg[13][79]  ( .D(n13495), .CK(N28803), .Q(n4079), .QN(
        n8814) );
  DFF_X1 \CACHE_MEM_reg[13][78]  ( .D(n13494), .CK(N28803), .Q(n4063), .QN(
        n8830) );
  DFF_X1 \CACHE_MEM_reg[13][77]  ( .D(n13493), .CK(N28803), .Q(n4043), .QN(
        n8846) );
  DFF_X1 \CACHE_MEM_reg[13][76]  ( .D(n13492), .CK(N28803), .Q(n4027), .QN(
        n8862) );
  DFF_X1 \CACHE_MEM_reg[13][75]  ( .D(n13491), .CK(N28803), .Q(n4002), .QN(
        n8878) );
  DFF_X1 \CACHE_MEM_reg[13][74]  ( .D(n13490), .CK(N28803), .Q(n3986), .QN(
        n8894) );
  DFF_X1 \CACHE_MEM_reg[13][73]  ( .D(n13489), .CK(N28803), .Q(n3966), .QN(
        n8910) );
  DFF_X1 \CACHE_MEM_reg[13][72]  ( .D(n13488), .CK(N28803), .Q(n3950), .QN(
        n8926) );
  DFF_X1 \CACHE_MEM_reg[13][71]  ( .D(n13487), .CK(N28803), .Q(n3930), .QN(
        n8942) );
  DFF_X1 \CACHE_MEM_reg[13][70]  ( .D(n13486), .CK(N28803), .Q(n3914), .QN(
        n8958) );
  DFF_X1 \CACHE_MEM_reg[13][69]  ( .D(n13485), .CK(N28803), .Q(n3894), .QN(
        n8974) );
  DFF_X1 \CACHE_MEM_reg[13][68]  ( .D(n13484), .CK(N28803), .Q(n3878), .QN(
        n8990) );
  DFF_X1 \CACHE_MEM_reg[13][67]  ( .D(n13483), .CK(N28803), .Q(n3853), .QN(
        n9006) );
  DFF_X1 \CACHE_MEM_reg[13][66]  ( .D(n13482), .CK(N28803), .Q(n3837), .QN(
        n9022) );
  DFF_X1 \CACHE_MEM_reg[13][65]  ( .D(n13481), .CK(N28803), .Q(n3817), .QN(
        n9038) );
  DFF_X1 \CACHE_MEM_reg[13][64]  ( .D(n13480), .CK(N28803), .Q(n3801), .QN(
        n9054) );
  DFF_X1 \CACHE_MEM_reg[13][63]  ( .D(n13479), .CK(N28803), .Q(n3559), .QN(
        n9070) );
  DFF_X1 \CACHE_MEM_reg[13][62]  ( .D(n13478), .CK(N28803), .Q(n3551), .QN(
        n9086) );
  DFF_X1 \CACHE_MEM_reg[13][61]  ( .D(n13477), .CK(N28803), .Q(n3547), .QN(
        n9102) );
  DFF_X1 \CACHE_MEM_reg[13][60]  ( .D(n13476), .CK(N28803), .Q(n3540), .QN(
        n9118) );
  DFF_X1 \CACHE_MEM_reg[13][59]  ( .D(n13475), .CK(N28803), .Q(n3530), .QN(
        n9134) );
  DFF_X1 \CACHE_MEM_reg[13][58]  ( .D(n13474), .CK(N28803), .Q(n3523), .QN(
        n9150) );
  DFF_X1 \CACHE_MEM_reg[13][57]  ( .D(n13473), .CK(N28803), .Q(n3519), .QN(
        n9166) );
  DFF_X1 \CACHE_MEM_reg[13][56]  ( .D(n13472), .CK(N28803), .Q(n3512), .QN(
        n9182) );
  DFF_X1 \CACHE_MEM_reg[13][55]  ( .D(n13471), .CK(N28803), .Q(n3506), .QN(
        n9198) );
  DFF_X1 \CACHE_MEM_reg[13][54]  ( .D(n13470), .CK(N28803), .Q(n3495), .QN(
        n9214) );
  DFF_X1 \CACHE_MEM_reg[13][53]  ( .D(n13469), .CK(N28803), .Q(n3491), .QN(
        n9230) );
  DFF_X1 \CACHE_MEM_reg[13][52]  ( .D(n13468), .CK(N28803), .Q(n3484), .QN(
        n9246) );
  DFF_X1 \CACHE_MEM_reg[13][51]  ( .D(n13467), .CK(N28803), .Q(n3478), .QN(
        n9262) );
  DFF_X1 \CACHE_MEM_reg[13][50]  ( .D(n13466), .CK(N28803), .Q(n3471), .QN(
        n9278) );
  DFF_X1 \CACHE_MEM_reg[13][49]  ( .D(n13465), .CK(N28803), .Q(n3467), .QN(
        n9294) );
  DFF_X1 \CACHE_MEM_reg[13][48]  ( .D(n13464), .CK(N28803), .Q(n3456), .QN(
        n9310) );
  DFF_X1 \CACHE_MEM_reg[13][47]  ( .D(n13463), .CK(N28803), .Q(n3450), .QN(
        n9326) );
  DFF_X1 \CACHE_MEM_reg[13][46]  ( .D(n13462), .CK(N28803), .Q(n3443), .QN(
        n9342) );
  DFF_X1 \CACHE_MEM_reg[13][45]  ( .D(n13461), .CK(N28803), .Q(n3439), .QN(
        n9358) );
  DFF_X1 \CACHE_MEM_reg[13][44]  ( .D(n13460), .CK(N28803), .Q(n3432), .QN(
        n9374) );
  DFF_X1 \CACHE_MEM_reg[13][43]  ( .D(n13459), .CK(N28803), .Q(n3417), .QN(
        n9390) );
  DFF_X1 \CACHE_MEM_reg[13][42]  ( .D(n13458), .CK(N28803), .Q(n3410), .QN(
        n9406) );
  DFF_X1 \CACHE_MEM_reg[13][41]  ( .D(n13457), .CK(N28803), .Q(n3406), .QN(
        n9422) );
  DFF_X1 \CACHE_MEM_reg[13][40]  ( .D(n13456), .CK(N28803), .Q(n3399), .QN(
        n9438) );
  DFF_X1 \CACHE_MEM_reg[13][39]  ( .D(n13455), .CK(N28803), .Q(n3393), .QN(
        n9454) );
  DFF_X1 \CACHE_MEM_reg[13][38]  ( .D(n13454), .CK(N28803), .Q(n3382), .QN(
        n9470) );
  DFF_X1 \CACHE_MEM_reg[13][37]  ( .D(n13453), .CK(N28803), .Q(n3378), .QN(
        n9486) );
  DFF_X1 \CACHE_MEM_reg[13][36]  ( .D(n13452), .CK(N28803), .Q(n3371), .QN(
        n9502) );
  DFF_X1 \CACHE_MEM_reg[13][35]  ( .D(n13451), .CK(N28803), .Q(n3365), .QN(
        n9518) );
  DFF_X1 \CACHE_MEM_reg[13][34]  ( .D(n13450), .CK(N28803), .Q(n3358), .QN(
        n9534) );
  DFF_X1 \CACHE_MEM_reg[13][33]  ( .D(n13449), .CK(N28803), .Q(n3354), .QN(
        n9550) );
  DFF_X1 \CACHE_MEM_reg[13][32]  ( .D(n13448), .CK(N28803), .Q(n3343), .QN(
        n9566) );
  DFF_X1 \CACHE_MEM_reg[13][31]  ( .D(n13447), .CK(N28803), .Q(n4819), .QN(
        n9582) );
  DFF_X1 \CACHE_MEM_reg[13][30]  ( .D(n13446), .CK(N28803), .Q(n4808), .QN(
        n9598) );
  DFF_X1 \CACHE_MEM_reg[13][29]  ( .D(n13445), .CK(N28803), .Q(n4791), .QN(
        n9614) );
  DFF_X1 \CACHE_MEM_reg[13][28]  ( .D(n13444), .CK(N28803), .Q(n4780), .QN(
        n9630) );
  DFF_X1 \CACHE_MEM_reg[13][27]  ( .D(n13443), .CK(N28803), .Q(n4758), .QN(
        n9646) );
  DFF_X1 \CACHE_MEM_reg[13][26]  ( .D(n13442), .CK(N28803), .Q(n4747), .QN(
        n9662) );
  DFF_X1 \CACHE_MEM_reg[13][25]  ( .D(n13441), .CK(N28803), .Q(n4734), .QN(
        n9678) );
  DFF_X1 \CACHE_MEM_reg[13][24]  ( .D(n13440), .CK(N28803), .Q(n4719), .QN(
        n9694) );
  DFF_X1 \CACHE_MEM_reg[13][23]  ( .D(n13439), .CK(N28803), .Q(n4706), .QN(
        n9710) );
  DFF_X1 \CACHE_MEM_reg[13][22]  ( .D(n13438), .CK(N28803), .Q(n4695), .QN(
        n9726) );
  DFF_X1 \CACHE_MEM_reg[13][21]  ( .D(n13437), .CK(N28803), .Q(n4678), .QN(
        n9742) );
  DFF_X1 \CACHE_MEM_reg[13][20]  ( .D(n13436), .CK(N28803), .Q(n4667), .QN(
        n9758) );
  DFF_X1 \CACHE_MEM_reg[13][19]  ( .D(n13435), .CK(N28803), .Q(n4650), .QN(
        n9774) );
  DFF_X1 \CACHE_MEM_reg[13][18]  ( .D(n13434), .CK(N28803), .Q(n4639), .QN(
        n9790) );
  DFF_X1 \CACHE_MEM_reg[13][17]  ( .D(n13433), .CK(N28803), .Q(n4626), .QN(
        n9806) );
  DFF_X1 \CACHE_MEM_reg[13][16]  ( .D(n13432), .CK(N28803), .Q(n4606), .QN(
        n9822) );
  DFF_X1 \CACHE_MEM_reg[13][15]  ( .D(n13431), .CK(N28803), .Q(n4593), .QN(
        n9838) );
  DFF_X1 \CACHE_MEM_reg[13][14]  ( .D(n13430), .CK(N28803), .Q(n4582), .QN(
        n9854) );
  DFF_X1 \CACHE_MEM_reg[13][13]  ( .D(n13429), .CK(N28803), .Q(n4565), .QN(
        n9870) );
  DFF_X1 \CACHE_MEM_reg[13][12]  ( .D(n13428), .CK(N28803), .Q(n4554), .QN(
        n9886) );
  DFF_X1 \CACHE_MEM_reg[13][11]  ( .D(n13427), .CK(N28803), .Q(n4537), .QN(
        n9902) );
  DFF_X1 \CACHE_MEM_reg[13][10]  ( .D(n13426), .CK(N28803), .Q(n4526), .QN(
        n9918) );
  DFF_X1 \CACHE_MEM_reg[13][9]  ( .D(n13425), .CK(N28803), .Q(n4513), .QN(
        n9934) );
  DFF_X1 \CACHE_MEM_reg[13][8]  ( .D(n13424), .CK(N28803), .Q(n4498), .QN(
        n9950) );
  DFF_X1 \CACHE_MEM_reg[13][7]  ( .D(n13423), .CK(N28803), .Q(n4485), .QN(
        n9966) );
  DFF_X1 \CACHE_MEM_reg[13][6]  ( .D(n13422), .CK(N28803), .Q(n4474), .QN(
        n9982) );
  DFF_X1 \CACHE_MEM_reg[13][5]  ( .D(n13421), .CK(N28803), .Q(n4452), .QN(
        n9998) );
  DFF_X1 \CACHE_MEM_reg[13][4]  ( .D(n13420), .CK(N28803), .Q(n4441), .QN(
        n10014) );
  DFF_X1 \CACHE_MEM_reg[13][3]  ( .D(n13419), .CK(N28803), .Q(n4424), .QN(
        n10030) );
  DFF_X1 \CACHE_MEM_reg[13][2]  ( .D(n13418), .CK(N28803), .Q(n4413), .QN(
        n10046) );
  DFF_X1 \CACHE_MEM_reg[13][1]  ( .D(n13417), .CK(N28803), .Q(n4400), .QN(
        n10062) );
  DFF_X1 \CACHE_MEM_reg[13][0]  ( .D(n13416), .CK(N28803), .Q(n4385), .QN(
        n10078) );
  DFF_X1 \CACHE_MEM_reg[12][255]  ( .D(n13415), .CK(N28803), .QN(n5994) );
  DFF_X1 \CACHE_MEM_reg[12][254]  ( .D(n13414), .CK(N28803), .QN(n6010) );
  DFF_X1 \CACHE_MEM_reg[12][253]  ( .D(n13413), .CK(N28803), .QN(n6026) );
  DFF_X1 \CACHE_MEM_reg[12][252]  ( .D(n13412), .CK(N28803), .QN(n6042) );
  DFF_X1 \CACHE_MEM_reg[12][251]  ( .D(n13411), .CK(N28803), .QN(n6058) );
  DFF_X1 \CACHE_MEM_reg[12][250]  ( .D(n13410), .CK(N28803), .QN(n6074) );
  DFF_X1 \CACHE_MEM_reg[12][249]  ( .D(n13409), .CK(N28803), .QN(n6090) );
  DFF_X1 \CACHE_MEM_reg[12][248]  ( .D(n13408), .CK(N28803), .QN(n6106) );
  DFF_X1 \CACHE_MEM_reg[12][247]  ( .D(n13407), .CK(N28803), .QN(n6122) );
  DFF_X1 \CACHE_MEM_reg[12][246]  ( .D(n13406), .CK(N28803), .QN(n6138) );
  DFF_X1 \CACHE_MEM_reg[12][245]  ( .D(n13405), .CK(N28803), .QN(n6154) );
  DFF_X1 \CACHE_MEM_reg[12][244]  ( .D(n13404), .CK(N28803), .QN(n6170) );
  DFF_X1 \CACHE_MEM_reg[12][243]  ( .D(n13403), .CK(N28803), .QN(n6186) );
  DFF_X1 \CACHE_MEM_reg[12][242]  ( .D(n13402), .CK(N28803), .QN(n6202) );
  DFF_X1 \CACHE_MEM_reg[12][241]  ( .D(n13401), .CK(N28803), .QN(n6218) );
  DFF_X1 \CACHE_MEM_reg[12][240]  ( .D(n13400), .CK(N28803), .QN(n6234) );
  DFF_X1 \CACHE_MEM_reg[12][239]  ( .D(n13399), .CK(N28803), .QN(n6250) );
  DFF_X1 \CACHE_MEM_reg[12][238]  ( .D(n13398), .CK(N28803), .QN(n6266) );
  DFF_X1 \CACHE_MEM_reg[12][237]  ( .D(n13397), .CK(N28803), .QN(n6282) );
  DFF_X1 \CACHE_MEM_reg[12][236]  ( .D(n13396), .CK(N28803), .QN(n6298) );
  DFF_X1 \CACHE_MEM_reg[12][235]  ( .D(n13395), .CK(N28803), .QN(n6314) );
  DFF_X1 \CACHE_MEM_reg[12][234]  ( .D(n13394), .CK(N28803), .QN(n6330) );
  DFF_X1 \CACHE_MEM_reg[12][233]  ( .D(n13393), .CK(N28803), .QN(n6346) );
  DFF_X1 \CACHE_MEM_reg[12][232]  ( .D(n13392), .CK(N28803), .QN(n6362) );
  DFF_X1 \CACHE_MEM_reg[12][231]  ( .D(n13391), .CK(N28803), .QN(n6378) );
  DFF_X1 \CACHE_MEM_reg[12][230]  ( .D(n13390), .CK(N28803), .QN(n6394) );
  DFF_X1 \CACHE_MEM_reg[12][229]  ( .D(n13389), .CK(N28803), .QN(n6410) );
  DFF_X1 \CACHE_MEM_reg[12][228]  ( .D(n13388), .CK(N28803), .QN(n6426) );
  DFF_X1 \CACHE_MEM_reg[12][227]  ( .D(n13387), .CK(N28803), .QN(n6442) );
  DFF_X1 \CACHE_MEM_reg[12][226]  ( .D(n13386), .CK(N28803), .QN(n6458) );
  DFF_X1 \CACHE_MEM_reg[12][225]  ( .D(n13385), .CK(N28803), .QN(n6474) );
  DFF_X1 \CACHE_MEM_reg[12][224]  ( .D(n13384), .CK(N28803), .QN(n6490) );
  DFF_X1 \CACHE_MEM_reg[12][223]  ( .D(n13383), .CK(N28803), .QN(n6506) );
  DFF_X1 \CACHE_MEM_reg[12][222]  ( .D(n13382), .CK(N28803), .QN(n6522) );
  DFF_X1 \CACHE_MEM_reg[12][221]  ( .D(n13381), .CK(N28803), .QN(n6538) );
  DFF_X1 \CACHE_MEM_reg[12][220]  ( .D(n13380), .CK(N28803), .QN(n6554) );
  DFF_X1 \CACHE_MEM_reg[12][219]  ( .D(n13379), .CK(N28803), .QN(n6570) );
  DFF_X1 \CACHE_MEM_reg[12][218]  ( .D(n13378), .CK(N28803), .QN(n6586) );
  DFF_X1 \CACHE_MEM_reg[12][217]  ( .D(n13377), .CK(N28803), .QN(n6602) );
  DFF_X1 \CACHE_MEM_reg[12][216]  ( .D(n13376), .CK(N28803), .QN(n6618) );
  DFF_X1 \CACHE_MEM_reg[12][215]  ( .D(n13375), .CK(N28803), .QN(n6634) );
  DFF_X1 \CACHE_MEM_reg[12][214]  ( .D(n13374), .CK(N28803), .QN(n6650) );
  DFF_X1 \CACHE_MEM_reg[12][213]  ( .D(n13373), .CK(N28803), .QN(n6666) );
  DFF_X1 \CACHE_MEM_reg[12][212]  ( .D(n13372), .CK(N28803), .QN(n6682) );
  DFF_X1 \CACHE_MEM_reg[12][211]  ( .D(n13371), .CK(N28803), .QN(n6698) );
  DFF_X1 \CACHE_MEM_reg[12][210]  ( .D(n13370), .CK(N28803), .QN(n6714) );
  DFF_X1 \CACHE_MEM_reg[12][209]  ( .D(n13369), .CK(N28803), .QN(n6730) );
  DFF_X1 \CACHE_MEM_reg[12][208]  ( .D(n13368), .CK(N28803), .QN(n6746) );
  DFF_X1 \CACHE_MEM_reg[12][207]  ( .D(n13367), .CK(N28803), .QN(n6762) );
  DFF_X1 \CACHE_MEM_reg[12][206]  ( .D(n13366), .CK(N28803), .QN(n6778) );
  DFF_X1 \CACHE_MEM_reg[12][205]  ( .D(n13365), .CK(N28803), .QN(n6794) );
  DFF_X1 \CACHE_MEM_reg[12][204]  ( .D(n13364), .CK(N28803), .QN(n6810) );
  DFF_X1 \CACHE_MEM_reg[12][203]  ( .D(n13363), .CK(N28803), .QN(n6826) );
  DFF_X1 \CACHE_MEM_reg[12][202]  ( .D(n13362), .CK(N28803), .QN(n6842) );
  DFF_X1 \CACHE_MEM_reg[12][201]  ( .D(n13361), .CK(N28803), .QN(n6858) );
  DFF_X1 \CACHE_MEM_reg[12][200]  ( .D(n13360), .CK(N28803), .QN(n6874) );
  DFF_X1 \CACHE_MEM_reg[12][199]  ( .D(n13359), .CK(N28803), .QN(n6890) );
  DFF_X1 \CACHE_MEM_reg[12][198]  ( .D(n13358), .CK(N28803), .QN(n6906) );
  DFF_X1 \CACHE_MEM_reg[12][197]  ( .D(n13357), .CK(N28803), .QN(n6922) );
  DFF_X1 \CACHE_MEM_reg[12][196]  ( .D(n13356), .CK(N28803), .QN(n6938) );
  DFF_X1 \CACHE_MEM_reg[12][195]  ( .D(n13355), .CK(N28803), .QN(n6954) );
  DFF_X1 \CACHE_MEM_reg[12][194]  ( .D(n13354), .CK(N28803), .QN(n6970) );
  DFF_X1 \CACHE_MEM_reg[12][193]  ( .D(n13353), .CK(N28803), .QN(n6986) );
  DFF_X1 \CACHE_MEM_reg[12][192]  ( .D(n13352), .CK(N28803), .QN(n7002) );
  DFF_X1 \CACHE_MEM_reg[12][191]  ( .D(n13351), .CK(N28803), .QN(n7018) );
  DFF_X1 \CACHE_MEM_reg[12][190]  ( .D(n13350), .CK(N28803), .QN(n7034) );
  DFF_X1 \CACHE_MEM_reg[12][189]  ( .D(n13349), .CK(N28803), .QN(n7050) );
  DFF_X1 \CACHE_MEM_reg[12][188]  ( .D(n13348), .CK(N28803), .QN(n7066) );
  DFF_X1 \CACHE_MEM_reg[12][187]  ( .D(n13347), .CK(N28803), .QN(n7082) );
  DFF_X1 \CACHE_MEM_reg[12][186]  ( .D(n13346), .CK(N28803), .QN(n7098) );
  DFF_X1 \CACHE_MEM_reg[12][185]  ( .D(n13345), .CK(N28803), .QN(n7114) );
  DFF_X1 \CACHE_MEM_reg[12][184]  ( .D(n13344), .CK(N28803), .QN(n7130) );
  DFF_X1 \CACHE_MEM_reg[12][183]  ( .D(n13343), .CK(N28803), .QN(n7146) );
  DFF_X1 \CACHE_MEM_reg[12][182]  ( .D(n13342), .CK(N28803), .QN(n7162) );
  DFF_X1 \CACHE_MEM_reg[12][181]  ( .D(n13341), .CK(N28803), .QN(n7178) );
  DFF_X1 \CACHE_MEM_reg[12][180]  ( .D(n13340), .CK(N28803), .QN(n7194) );
  DFF_X1 \CACHE_MEM_reg[12][179]  ( .D(n13339), .CK(N28803), .QN(n7210) );
  DFF_X1 \CACHE_MEM_reg[12][178]  ( .D(n13338), .CK(N28803), .QN(n7226) );
  DFF_X1 \CACHE_MEM_reg[12][177]  ( .D(n13337), .CK(N28803), .QN(n7242) );
  DFF_X1 \CACHE_MEM_reg[12][176]  ( .D(n13336), .CK(N28803), .QN(n7258) );
  DFF_X1 \CACHE_MEM_reg[12][175]  ( .D(n13335), .CK(N28803), .QN(n7274) );
  DFF_X1 \CACHE_MEM_reg[12][174]  ( .D(n13334), .CK(N28803), .QN(n7290) );
  DFF_X1 \CACHE_MEM_reg[12][173]  ( .D(n13333), .CK(N28803), .QN(n7306) );
  DFF_X1 \CACHE_MEM_reg[12][172]  ( .D(n13332), .CK(N28803), .QN(n7322) );
  DFF_X1 \CACHE_MEM_reg[12][171]  ( .D(n13331), .CK(N28803), .QN(n7338) );
  DFF_X1 \CACHE_MEM_reg[12][170]  ( .D(n13330), .CK(N28803), .QN(n7354) );
  DFF_X1 \CACHE_MEM_reg[12][169]  ( .D(n13329), .CK(N28803), .QN(n7370) );
  DFF_X1 \CACHE_MEM_reg[12][168]  ( .D(n13328), .CK(N28803), .QN(n7386) );
  DFF_X1 \CACHE_MEM_reg[12][167]  ( .D(n13327), .CK(N28803), .QN(n7402) );
  DFF_X1 \CACHE_MEM_reg[12][166]  ( .D(n13326), .CK(N28803), .QN(n7418) );
  DFF_X1 \CACHE_MEM_reg[12][165]  ( .D(n13325), .CK(N28803), .QN(n7434) );
  DFF_X1 \CACHE_MEM_reg[12][164]  ( .D(n13324), .CK(N28803), .QN(n7450) );
  DFF_X1 \CACHE_MEM_reg[12][163]  ( .D(n13323), .CK(N28803), .QN(n7466) );
  DFF_X1 \CACHE_MEM_reg[12][162]  ( .D(n13322), .CK(N28803), .QN(n7482) );
  DFF_X1 \CACHE_MEM_reg[12][161]  ( .D(n13321), .CK(N28803), .QN(n7498) );
  DFF_X1 \CACHE_MEM_reg[12][160]  ( .D(n13320), .CK(N28803), .QN(n7514) );
  DFF_X1 \CACHE_MEM_reg[12][159]  ( .D(n13319), .CK(N28803), .QN(n7530) );
  DFF_X1 \CACHE_MEM_reg[12][158]  ( .D(n13318), .CK(N28803), .QN(n7546) );
  DFF_X1 \CACHE_MEM_reg[12][157]  ( .D(n13317), .CK(N28803), .QN(n7562) );
  DFF_X1 \CACHE_MEM_reg[12][156]  ( .D(n13316), .CK(N28803), .QN(n7578) );
  DFF_X1 \CACHE_MEM_reg[12][155]  ( .D(n13315), .CK(N28803), .QN(n7594) );
  DFF_X1 \CACHE_MEM_reg[12][154]  ( .D(n13314), .CK(N28803), .QN(n7610) );
  DFF_X1 \CACHE_MEM_reg[12][153]  ( .D(n13313), .CK(N28803), .QN(n7626) );
  DFF_X1 \CACHE_MEM_reg[12][152]  ( .D(n13312), .CK(N28803), .QN(n7642) );
  DFF_X1 \CACHE_MEM_reg[12][151]  ( .D(n13311), .CK(N28803), .QN(n7658) );
  DFF_X1 \CACHE_MEM_reg[12][150]  ( .D(n13310), .CK(N28803), .QN(n7674) );
  DFF_X1 \CACHE_MEM_reg[12][149]  ( .D(n13309), .CK(N28803), .QN(n7690) );
  DFF_X1 \CACHE_MEM_reg[12][148]  ( .D(n13308), .CK(N28803), .QN(n7706) );
  DFF_X1 \CACHE_MEM_reg[12][147]  ( .D(n13307), .CK(N28803), .QN(n7722) );
  DFF_X1 \CACHE_MEM_reg[12][146]  ( .D(n13306), .CK(N28803), .QN(n7738) );
  DFF_X1 \CACHE_MEM_reg[12][145]  ( .D(n13305), .CK(N28803), .QN(n7754) );
  DFF_X1 \CACHE_MEM_reg[12][144]  ( .D(n13304), .CK(N28803), .QN(n7770) );
  DFF_X1 \CACHE_MEM_reg[12][143]  ( .D(n13303), .CK(N28803), .QN(n7786) );
  DFF_X1 \CACHE_MEM_reg[12][142]  ( .D(n13302), .CK(N28803), .QN(n7802) );
  DFF_X1 \CACHE_MEM_reg[12][141]  ( .D(n13301), .CK(N28803), .QN(n7818) );
  DFF_X1 \CACHE_MEM_reg[12][140]  ( .D(n13300), .CK(N28803), .QN(n7834) );
  DFF_X1 \CACHE_MEM_reg[12][139]  ( .D(n13299), .CK(N28803), .QN(n7850) );
  DFF_X1 \CACHE_MEM_reg[12][138]  ( .D(n13298), .CK(N28803), .QN(n7866) );
  DFF_X1 \CACHE_MEM_reg[12][137]  ( .D(n13297), .CK(N28803), .QN(n7882) );
  DFF_X1 \CACHE_MEM_reg[12][136]  ( .D(n13296), .CK(N28803), .QN(n7898) );
  DFF_X1 \CACHE_MEM_reg[12][135]  ( .D(n13295), .CK(N28803), .QN(n7914) );
  DFF_X1 \CACHE_MEM_reg[12][134]  ( .D(n13294), .CK(N28803), .QN(n7930) );
  DFF_X1 \CACHE_MEM_reg[12][133]  ( .D(n13293), .CK(N28803), .QN(n7946) );
  DFF_X1 \CACHE_MEM_reg[12][132]  ( .D(n13292), .CK(N28803), .QN(n7962) );
  DFF_X1 \CACHE_MEM_reg[12][131]  ( .D(n13291), .CK(N28803), .QN(n7978) );
  DFF_X1 \CACHE_MEM_reg[12][130]  ( .D(n13290), .CK(N28803), .QN(n7994) );
  DFF_X1 \CACHE_MEM_reg[12][129]  ( .D(n13289), .CK(N28803), .QN(n8010) );
  DFF_X1 \CACHE_MEM_reg[12][128]  ( .D(n13288), .CK(N28803), .QN(n8026) );
  DFF_X1 \CACHE_MEM_reg[12][127]  ( .D(n13287), .CK(N28803), .QN(n8042) );
  DFF_X1 \CACHE_MEM_reg[12][126]  ( .D(n13286), .CK(N28803), .QN(n8058) );
  DFF_X1 \CACHE_MEM_reg[12][125]  ( .D(n13285), .CK(N28803), .QN(n8074) );
  DFF_X1 \CACHE_MEM_reg[12][124]  ( .D(n13284), .CK(N28803), .QN(n8090) );
  DFF_X1 \CACHE_MEM_reg[12][123]  ( .D(n13283), .CK(N28803), .QN(n8106) );
  DFF_X1 \CACHE_MEM_reg[12][122]  ( .D(n13282), .CK(N28803), .QN(n8122) );
  DFF_X1 \CACHE_MEM_reg[12][121]  ( .D(n13281), .CK(N28803), .QN(n8138) );
  DFF_X1 \CACHE_MEM_reg[12][120]  ( .D(n13280), .CK(N28803), .QN(n8154) );
  DFF_X1 \CACHE_MEM_reg[12][119]  ( .D(n13279), .CK(N28803), .QN(n8170) );
  DFF_X1 \CACHE_MEM_reg[12][118]  ( .D(n13278), .CK(N28803), .QN(n8186) );
  DFF_X1 \CACHE_MEM_reg[12][117]  ( .D(n13277), .CK(N28803), .QN(n8202) );
  DFF_X1 \CACHE_MEM_reg[12][116]  ( .D(n13276), .CK(N28803), .QN(n8218) );
  DFF_X1 \CACHE_MEM_reg[12][115]  ( .D(n13275), .CK(N28803), .QN(n8234) );
  DFF_X1 \CACHE_MEM_reg[12][114]  ( .D(n13274), .CK(N28803), .QN(n8250) );
  DFF_X1 \CACHE_MEM_reg[12][113]  ( .D(n13273), .CK(N28803), .QN(n8266) );
  DFF_X1 \CACHE_MEM_reg[12][112]  ( .D(n13272), .CK(N28803), .QN(n8282) );
  DFF_X1 \CACHE_MEM_reg[12][111]  ( .D(n13271), .CK(N28803), .QN(n8298) );
  DFF_X1 \CACHE_MEM_reg[12][110]  ( .D(n13270), .CK(N28803), .QN(n8314) );
  DFF_X1 \CACHE_MEM_reg[12][109]  ( .D(n13269), .CK(N28803), .QN(n8330) );
  DFF_X1 \CACHE_MEM_reg[12][108]  ( .D(n13268), .CK(N28803), .QN(n8346) );
  DFF_X1 \CACHE_MEM_reg[12][107]  ( .D(n13267), .CK(N28803), .QN(n8362) );
  DFF_X1 \CACHE_MEM_reg[12][106]  ( .D(n13266), .CK(N28803), .QN(n8378) );
  DFF_X1 \CACHE_MEM_reg[12][105]  ( .D(n13265), .CK(N28803), .QN(n8394) );
  DFF_X1 \CACHE_MEM_reg[12][104]  ( .D(n13264), .CK(N28803), .QN(n8410) );
  DFF_X1 \CACHE_MEM_reg[12][103]  ( .D(n13263), .CK(N28803), .QN(n8426) );
  DFF_X1 \CACHE_MEM_reg[12][102]  ( .D(n13262), .CK(N28803), .QN(n8442) );
  DFF_X1 \CACHE_MEM_reg[12][101]  ( .D(n13261), .CK(N28803), .QN(n8458) );
  DFF_X1 \CACHE_MEM_reg[12][100]  ( .D(n13260), .CK(N28803), .QN(n8474) );
  DFF_X1 \CACHE_MEM_reg[12][99]  ( .D(n13259), .CK(N28803), .QN(n8490) );
  DFF_X1 \CACHE_MEM_reg[12][98]  ( .D(n13258), .CK(N28803), .QN(n8506) );
  DFF_X1 \CACHE_MEM_reg[12][97]  ( .D(n13257), .CK(N28803), .QN(n8522) );
  DFF_X1 \CACHE_MEM_reg[12][96]  ( .D(n13256), .CK(N28803), .QN(n8538) );
  DFF_X1 \CACHE_MEM_reg[12][95]  ( .D(n13255), .CK(N28803), .QN(n8554) );
  DFF_X1 \CACHE_MEM_reg[12][94]  ( .D(n13254), .CK(N28803), .QN(n8570) );
  DFF_X1 \CACHE_MEM_reg[12][93]  ( .D(n13253), .CK(N28803), .QN(n8586) );
  DFF_X1 \CACHE_MEM_reg[12][92]  ( .D(n13252), .CK(N28803), .QN(n8602) );
  DFF_X1 \CACHE_MEM_reg[12][91]  ( .D(n13251), .CK(N28803), .QN(n8618) );
  DFF_X1 \CACHE_MEM_reg[12][90]  ( .D(n13250), .CK(N28803), .QN(n8634) );
  DFF_X1 \CACHE_MEM_reg[12][89]  ( .D(n13249), .CK(N28803), .QN(n8650) );
  DFF_X1 \CACHE_MEM_reg[12][88]  ( .D(n13248), .CK(N28803), .QN(n8666) );
  DFF_X1 \CACHE_MEM_reg[12][87]  ( .D(n13247), .CK(N28803), .QN(n8682) );
  DFF_X1 \CACHE_MEM_reg[12][86]  ( .D(n13246), .CK(N28803), .QN(n8698) );
  DFF_X1 \CACHE_MEM_reg[12][85]  ( .D(n13245), .CK(N28803), .QN(n8714) );
  DFF_X1 \CACHE_MEM_reg[12][84]  ( .D(n13244), .CK(N28803), .QN(n8730) );
  DFF_X1 \CACHE_MEM_reg[12][83]  ( .D(n13243), .CK(N28803), .QN(n8746) );
  DFF_X1 \CACHE_MEM_reg[12][82]  ( .D(n13242), .CK(N28803), .QN(n8762) );
  DFF_X1 \CACHE_MEM_reg[12][81]  ( .D(n13241), .CK(N28803), .QN(n8778) );
  DFF_X1 \CACHE_MEM_reg[12][80]  ( .D(n13240), .CK(N28803), .QN(n8794) );
  DFF_X1 \CACHE_MEM_reg[12][79]  ( .D(n13239), .CK(N28803), .QN(n8810) );
  DFF_X1 \CACHE_MEM_reg[12][78]  ( .D(n13238), .CK(N28803), .QN(n8826) );
  DFF_X1 \CACHE_MEM_reg[12][77]  ( .D(n13237), .CK(N28803), .QN(n8842) );
  DFF_X1 \CACHE_MEM_reg[12][76]  ( .D(n13236), .CK(N28803), .QN(n8858) );
  DFF_X1 \CACHE_MEM_reg[12][75]  ( .D(n13235), .CK(N28803), .QN(n8874) );
  DFF_X1 \CACHE_MEM_reg[12][74]  ( .D(n13234), .CK(N28803), .QN(n8890) );
  DFF_X1 \CACHE_MEM_reg[12][73]  ( .D(n13233), .CK(N28803), .QN(n8906) );
  DFF_X1 \CACHE_MEM_reg[12][72]  ( .D(n13232), .CK(N28803), .QN(n8922) );
  DFF_X1 \CACHE_MEM_reg[12][71]  ( .D(n13231), .CK(N28803), .QN(n8938) );
  DFF_X1 \CACHE_MEM_reg[12][70]  ( .D(n13230), .CK(N28803), .QN(n8954) );
  DFF_X1 \CACHE_MEM_reg[12][69]  ( .D(n13229), .CK(N28803), .QN(n8970) );
  DFF_X1 \CACHE_MEM_reg[12][68]  ( .D(n13228), .CK(N28803), .QN(n8986) );
  DFF_X1 \CACHE_MEM_reg[12][67]  ( .D(n13227), .CK(N28803), .QN(n9002) );
  DFF_X1 \CACHE_MEM_reg[12][66]  ( .D(n13226), .CK(N28803), .QN(n9018) );
  DFF_X1 \CACHE_MEM_reg[12][65]  ( .D(n13225), .CK(N28803), .QN(n9034) );
  DFF_X1 \CACHE_MEM_reg[12][64]  ( .D(n13224), .CK(N28803), .QN(n9050) );
  DFF_X1 \CACHE_MEM_reg[12][63]  ( .D(n13223), .CK(N28803), .QN(n9066) );
  DFF_X1 \CACHE_MEM_reg[12][62]  ( .D(n13222), .CK(N28803), .QN(n9082) );
  DFF_X1 \CACHE_MEM_reg[12][61]  ( .D(n13221), .CK(N28803), .QN(n9098) );
  DFF_X1 \CACHE_MEM_reg[12][60]  ( .D(n13220), .CK(N28803), .QN(n9114) );
  DFF_X1 \CACHE_MEM_reg[12][59]  ( .D(n13219), .CK(N28803), .QN(n9130) );
  DFF_X1 \CACHE_MEM_reg[12][58]  ( .D(n13218), .CK(N28803), .QN(n9146) );
  DFF_X1 \CACHE_MEM_reg[12][57]  ( .D(n13217), .CK(N28803), .QN(n9162) );
  DFF_X1 \CACHE_MEM_reg[12][56]  ( .D(n13216), .CK(N28803), .QN(n9178) );
  DFF_X1 \CACHE_MEM_reg[12][55]  ( .D(n13215), .CK(N28803), .QN(n9194) );
  DFF_X1 \CACHE_MEM_reg[12][54]  ( .D(n13214), .CK(N28803), .QN(n9210) );
  DFF_X1 \CACHE_MEM_reg[12][53]  ( .D(n13213), .CK(N28803), .QN(n9226) );
  DFF_X1 \CACHE_MEM_reg[12][52]  ( .D(n13212), .CK(N28803), .QN(n9242) );
  DFF_X1 \CACHE_MEM_reg[12][51]  ( .D(n13211), .CK(N28803), .QN(n9258) );
  DFF_X1 \CACHE_MEM_reg[12][50]  ( .D(n13210), .CK(N28803), .QN(n9274) );
  DFF_X1 \CACHE_MEM_reg[12][49]  ( .D(n13209), .CK(N28803), .QN(n9290) );
  DFF_X1 \CACHE_MEM_reg[12][48]  ( .D(n13208), .CK(N28803), .QN(n9306) );
  DFF_X1 \CACHE_MEM_reg[12][47]  ( .D(n13207), .CK(N28803), .QN(n9322) );
  DFF_X1 \CACHE_MEM_reg[12][46]  ( .D(n13206), .CK(N28803), .QN(n9338) );
  DFF_X1 \CACHE_MEM_reg[12][45]  ( .D(n13205), .CK(N28803), .QN(n9354) );
  DFF_X1 \CACHE_MEM_reg[12][44]  ( .D(n13204), .CK(N28803), .QN(n9370) );
  DFF_X1 \CACHE_MEM_reg[12][43]  ( .D(n13203), .CK(N28803), .QN(n9386) );
  DFF_X1 \CACHE_MEM_reg[12][42]  ( .D(n13202), .CK(N28803), .QN(n9402) );
  DFF_X1 \CACHE_MEM_reg[12][41]  ( .D(n13201), .CK(N28803), .QN(n9418) );
  DFF_X1 \CACHE_MEM_reg[12][40]  ( .D(n13200), .CK(N28803), .QN(n9434) );
  DFF_X1 \CACHE_MEM_reg[12][39]  ( .D(n13199), .CK(N28803), .QN(n9450) );
  DFF_X1 \CACHE_MEM_reg[12][38]  ( .D(n13198), .CK(N28803), .QN(n9466) );
  DFF_X1 \CACHE_MEM_reg[12][37]  ( .D(n13197), .CK(N28803), .QN(n9482) );
  DFF_X1 \CACHE_MEM_reg[12][36]  ( .D(n13196), .CK(N28803), .QN(n9498) );
  DFF_X1 \CACHE_MEM_reg[12][35]  ( .D(n13195), .CK(N28803), .QN(n9514) );
  DFF_X1 \CACHE_MEM_reg[12][34]  ( .D(n13194), .CK(N28803), .QN(n9530) );
  DFF_X1 \CACHE_MEM_reg[12][33]  ( .D(n13193), .CK(N28803), .QN(n9546) );
  DFF_X1 \CACHE_MEM_reg[12][32]  ( .D(n13192), .CK(N28803), .QN(n9562) );
  DFF_X1 \CACHE_MEM_reg[12][31]  ( .D(n13191), .CK(N28803), .QN(n9578) );
  DFF_X1 \CACHE_MEM_reg[12][30]  ( .D(n13190), .CK(N28803), .QN(n9594) );
  DFF_X1 \CACHE_MEM_reg[12][29]  ( .D(n13189), .CK(N28803), .QN(n9610) );
  DFF_X1 \CACHE_MEM_reg[12][28]  ( .D(n13188), .CK(N28803), .QN(n9626) );
  DFF_X1 \CACHE_MEM_reg[12][27]  ( .D(n13187), .CK(N28803), .QN(n9642) );
  DFF_X1 \CACHE_MEM_reg[12][26]  ( .D(n13186), .CK(N28803), .QN(n9658) );
  DFF_X1 \CACHE_MEM_reg[12][25]  ( .D(n13185), .CK(N28803), .QN(n9674) );
  DFF_X1 \CACHE_MEM_reg[12][24]  ( .D(n13184), .CK(N28803), .QN(n9690) );
  DFF_X1 \CACHE_MEM_reg[12][23]  ( .D(n13183), .CK(N28803), .QN(n9706) );
  DFF_X1 \CACHE_MEM_reg[12][22]  ( .D(n13182), .CK(N28803), .QN(n9722) );
  DFF_X1 \CACHE_MEM_reg[12][21]  ( .D(n13181), .CK(N28803), .QN(n9738) );
  DFF_X1 \CACHE_MEM_reg[12][20]  ( .D(n13180), .CK(N28803), .QN(n9754) );
  DFF_X1 \CACHE_MEM_reg[12][19]  ( .D(n13179), .CK(N28803), .QN(n9770) );
  DFF_X1 \CACHE_MEM_reg[12][18]  ( .D(n13178), .CK(N28803), .QN(n9786) );
  DFF_X1 \CACHE_MEM_reg[12][17]  ( .D(n13177), .CK(N28803), .QN(n9802) );
  DFF_X1 \CACHE_MEM_reg[12][16]  ( .D(n13176), .CK(N28803), .QN(n9818) );
  DFF_X1 \CACHE_MEM_reg[12][15]  ( .D(n13175), .CK(N28803), .QN(n9834) );
  DFF_X1 \CACHE_MEM_reg[12][14]  ( .D(n13174), .CK(N28803), .QN(n9850) );
  DFF_X1 \CACHE_MEM_reg[12][13]  ( .D(n13173), .CK(N28803), .QN(n9866) );
  DFF_X1 \CACHE_MEM_reg[12][12]  ( .D(n13172), .CK(N28803), .QN(n9882) );
  DFF_X1 \CACHE_MEM_reg[12][11]  ( .D(n13171), .CK(N28803), .QN(n9898) );
  DFF_X1 \CACHE_MEM_reg[12][10]  ( .D(n13170), .CK(N28803), .QN(n9914) );
  DFF_X1 \CACHE_MEM_reg[12][9]  ( .D(n13169), .CK(N28803), .QN(n9930) );
  DFF_X1 \CACHE_MEM_reg[12][8]  ( .D(n13168), .CK(N28803), .QN(n9946) );
  DFF_X1 \CACHE_MEM_reg[12][7]  ( .D(n13167), .CK(N28803), .QN(n9962) );
  DFF_X1 \CACHE_MEM_reg[12][6]  ( .D(n13166), .CK(N28803), .QN(n9978) );
  DFF_X1 \CACHE_MEM_reg[12][5]  ( .D(n13165), .CK(N28803), .QN(n9994) );
  DFF_X1 \CACHE_MEM_reg[12][4]  ( .D(n13164), .CK(N28803), .QN(n10010) );
  DFF_X1 \CACHE_MEM_reg[12][3]  ( .D(n13163), .CK(N28803), .QN(n10026) );
  DFF_X1 \CACHE_MEM_reg[12][2]  ( .D(n13162), .CK(N28803), .QN(n10042) );
  DFF_X1 \CACHE_MEM_reg[12][1]  ( .D(n13161), .CK(N28803), .QN(n10058) );
  DFF_X1 \CACHE_MEM_reg[12][0]  ( .D(n13160), .CK(N28803), .QN(n10074) );
  DFF_X1 \CACHE_MEM_reg[11][255]  ( .D(n13159), .CK(N28803), .Q(n5264), .QN(
        n6004) );
  DFF_X1 \CACHE_MEM_reg[11][254]  ( .D(n13158), .CK(N28803), .Q(n5247), .QN(
        n6020) );
  DFF_X1 \CACHE_MEM_reg[11][253]  ( .D(n13157), .CK(N28803), .Q(n5236), .QN(
        n6036) );
  DFF_X1 \CACHE_MEM_reg[11][252]  ( .D(n13156), .CK(N28803), .Q(n5223), .QN(
        n6052) );
  DFF_X1 \CACHE_MEM_reg[11][251]  ( .D(n13155), .CK(N28803), .Q(n5203), .QN(
        n6068) );
  DFF_X1 \CACHE_MEM_reg[11][250]  ( .D(n13154), .CK(N28803), .Q(n5190), .QN(
        n6084) );
  DFF_X1 \CACHE_MEM_reg[11][249]  ( .D(n13153), .CK(N28803), .Q(n5179), .QN(
        n6100) );
  DFF_X1 \CACHE_MEM_reg[11][248]  ( .D(n13152), .CK(N28803), .Q(n5162), .QN(
        n6116) );
  DFF_X1 \CACHE_MEM_reg[11][247]  ( .D(n13151), .CK(N28803), .Q(n5151), .QN(
        n6132) );
  DFF_X1 \CACHE_MEM_reg[11][246]  ( .D(n13150), .CK(N28803), .Q(n5134), .QN(
        n6148) );
  DFF_X1 \CACHE_MEM_reg[11][245]  ( .D(n13149), .CK(N28803), .Q(n5123), .QN(
        n6164) );
  DFF_X1 \CACHE_MEM_reg[11][244]  ( .D(n13148), .CK(N28803), .Q(n5110), .QN(
        n6180) );
  DFF_X1 \CACHE_MEM_reg[11][243]  ( .D(n13147), .CK(N28803), .Q(n5095), .QN(
        n6196) );
  DFF_X1 \CACHE_MEM_reg[11][242]  ( .D(n13146), .CK(N28803), .Q(n5082), .QN(
        n6212) );
  DFF_X1 \CACHE_MEM_reg[11][241]  ( .D(n13145), .CK(N28803), .Q(n5071), .QN(
        n6228) );
  DFF_X1 \CACHE_MEM_reg[11][240]  ( .D(n13144), .CK(N28803), .Q(n5719), .QN(
        n6244) );
  DFF_X1 \CACHE_MEM_reg[11][239]  ( .D(n13143), .CK(N28803), .Q(n5041), .QN(
        n6260) );
  DFF_X1 \CACHE_MEM_reg[11][238]  ( .D(n13142), .CK(N28803), .Q(n5030), .QN(
        n6276) );
  DFF_X1 \CACHE_MEM_reg[11][237]  ( .D(n13141), .CK(N28803), .Q(n5013), .QN(
        n6292) );
  DFF_X1 \CACHE_MEM_reg[11][236]  ( .D(n13140), .CK(N28803), .Q(n5002), .QN(
        n6308) );
  DFF_X1 \CACHE_MEM_reg[11][235]  ( .D(n13139), .CK(N28803), .Q(n4985), .QN(
        n6324) );
  DFF_X1 \CACHE_MEM_reg[11][234]  ( .D(n13138), .CK(N28803), .Q(n4974), .QN(
        n6340) );
  DFF_X1 \CACHE_MEM_reg[11][233]  ( .D(n13137), .CK(N28803), .Q(n4961), .QN(
        n6356) );
  DFF_X1 \CACHE_MEM_reg[11][232]  ( .D(n13136), .CK(N28803), .Q(n4946), .QN(
        n6372) );
  DFF_X1 \CACHE_MEM_reg[11][231]  ( .D(n13135), .CK(N28803), .Q(n4933), .QN(
        n6388) );
  DFF_X1 \CACHE_MEM_reg[11][230]  ( .D(n13134), .CK(N28803), .Q(n4922), .QN(
        n6404) );
  DFF_X1 \CACHE_MEM_reg[11][229]  ( .D(n13133), .CK(N28803), .Q(n4900), .QN(
        n6420) );
  DFF_X1 \CACHE_MEM_reg[11][228]  ( .D(n13132), .CK(N28803), .Q(n4889), .QN(
        n6436) );
  DFF_X1 \CACHE_MEM_reg[11][227]  ( .D(n13131), .CK(N28803), .Q(n4872), .QN(
        n6452) );
  DFF_X1 \CACHE_MEM_reg[11][226]  ( .D(n13130), .CK(N28803), .Q(n4861), .QN(
        n6468) );
  DFF_X1 \CACHE_MEM_reg[11][225]  ( .D(n13129), .CK(N28803), .Q(n4848), .QN(
        n6484) );
  DFF_X1 \CACHE_MEM_reg[11][224]  ( .D(n13128), .CK(N28803), .Q(n4833), .QN(
        n6500) );
  DFF_X1 \CACHE_MEM_reg[11][223]  ( .D(n13127), .CK(N28803), .Q(n5267), .QN(
        n6516) );
  DFF_X1 \CACHE_MEM_reg[11][222]  ( .D(n13126), .CK(N28803), .Q(n5256), .QN(
        n6532) );
  DFF_X1 \CACHE_MEM_reg[11][221]  ( .D(n13125), .CK(N28803), .Q(n5239), .QN(
        n6548) );
  DFF_X1 \CACHE_MEM_reg[11][220]  ( .D(n13124), .CK(N28803), .Q(n5228), .QN(
        n6564) );
  DFF_X1 \CACHE_MEM_reg[11][219]  ( .D(n13123), .CK(N28803), .Q(n5206), .QN(
        n6580) );
  DFF_X1 \CACHE_MEM_reg[11][218]  ( .D(n13122), .CK(N28803), .Q(n5195), .QN(
        n6596) );
  DFF_X1 \CACHE_MEM_reg[11][217]  ( .D(n13121), .CK(N28803), .Q(n5182), .QN(
        n6612) );
  DFF_X1 \CACHE_MEM_reg[11][216]  ( .D(n13120), .CK(N28803), .Q(n5167), .QN(
        n6628) );
  DFF_X1 \CACHE_MEM_reg[11][215]  ( .D(n13119), .CK(N28803), .Q(n5154), .QN(
        n6644) );
  DFF_X1 \CACHE_MEM_reg[11][214]  ( .D(n13118), .CK(N28803), .Q(n5143), .QN(
        n6660) );
  DFF_X1 \CACHE_MEM_reg[11][213]  ( .D(n13117), .CK(N28803), .Q(n5126), .QN(
        n6676) );
  DFF_X1 \CACHE_MEM_reg[11][212]  ( .D(n13116), .CK(N28803), .Q(n5115), .QN(
        n6692) );
  DFF_X1 \CACHE_MEM_reg[11][211]  ( .D(n13115), .CK(N28803), .Q(n5098), .QN(
        n6708) );
  DFF_X1 \CACHE_MEM_reg[11][210]  ( .D(n13114), .CK(N28803), .Q(n5087), .QN(
        n6724) );
  DFF_X1 \CACHE_MEM_reg[11][209]  ( .D(n13113), .CK(N28803), .Q(n5074), .QN(
        n6740) );
  DFF_X1 \CACHE_MEM_reg[11][208]  ( .D(n13112), .CK(N28803), .Q(n5054), .QN(
        n6756) );
  DFF_X1 \CACHE_MEM_reg[11][207]  ( .D(n13111), .CK(N28803), .Q(n5046), .QN(
        n6772) );
  DFF_X1 \CACHE_MEM_reg[11][206]  ( .D(n13110), .CK(N28803), .Q(n5033), .QN(
        n6788) );
  DFF_X1 \CACHE_MEM_reg[11][205]  ( .D(n13109), .CK(N28803), .Q(n5018), .QN(
        n6804) );
  DFF_X1 \CACHE_MEM_reg[11][204]  ( .D(n13108), .CK(N28803), .Q(n5005), .QN(
        n6820) );
  DFF_X1 \CACHE_MEM_reg[11][203]  ( .D(n13107), .CK(N28803), .Q(n4994), .QN(
        n6836) );
  DFF_X1 \CACHE_MEM_reg[11][202]  ( .D(n13106), .CK(N28803), .Q(n4977), .QN(
        n6852) );
  DFF_X1 \CACHE_MEM_reg[11][201]  ( .D(n13105), .CK(N28803), .Q(n4966), .QN(
        n6868) );
  DFF_X1 \CACHE_MEM_reg[11][200]  ( .D(n13104), .CK(N28803), .Q(n4949), .QN(
        n6884) );
  DFF_X1 \CACHE_MEM_reg[11][199]  ( .D(n13103), .CK(N28803), .Q(n4938), .QN(
        n6900) );
  DFF_X1 \CACHE_MEM_reg[11][198]  ( .D(n13102), .CK(N28803), .Q(n4925), .QN(
        n6916) );
  DFF_X1 \CACHE_MEM_reg[11][197]  ( .D(n13101), .CK(N28803), .Q(n4905), .QN(
        n6932) );
  DFF_X1 \CACHE_MEM_reg[11][196]  ( .D(n13100), .CK(N28803), .Q(n4892), .QN(
        n6948) );
  DFF_X1 \CACHE_MEM_reg[11][195]  ( .D(n13099), .CK(N28803), .Q(n4881), .QN(
        n6964) );
  DFF_X1 \CACHE_MEM_reg[11][194]  ( .D(n13098), .CK(N28803), .Q(n4864), .QN(
        n6980) );
  DFF_X1 \CACHE_MEM_reg[11][193]  ( .D(n13097), .CK(N28803), .Q(n4853), .QN(
        n6996) );
  DFF_X1 \CACHE_MEM_reg[11][192]  ( .D(n13096), .CK(N28803), .Q(n4836), .QN(
        n7012) );
  DFF_X1 \CACHE_MEM_reg[11][191]  ( .D(n13095), .CK(N28803), .Q(n5711), .QN(
        n7028) );
  DFF_X1 \CACHE_MEM_reg[11][190]  ( .D(n13094), .CK(N28803), .Q(n5694), .QN(
        n7044) );
  DFF_X1 \CACHE_MEM_reg[11][189]  ( .D(n13093), .CK(N28803), .Q(n5683), .QN(
        n7060) );
  DFF_X1 \CACHE_MEM_reg[11][188]  ( .D(n13092), .CK(N28803), .Q(n5670), .QN(
        n7076) );
  DFF_X1 \CACHE_MEM_reg[11][187]  ( .D(n13091), .CK(N28803), .Q(n5650), .QN(
        n7092) );
  DFF_X1 \CACHE_MEM_reg[11][186]  ( .D(n13090), .CK(N28803), .Q(n5637), .QN(
        n7108) );
  DFF_X1 \CACHE_MEM_reg[11][185]  ( .D(n13089), .CK(N28803), .Q(n5626), .QN(
        n7124) );
  DFF_X1 \CACHE_MEM_reg[11][184]  ( .D(n13088), .CK(N28803), .Q(n5609), .QN(
        n7140) );
  DFF_X1 \CACHE_MEM_reg[11][183]  ( .D(n13087), .CK(N28803), .Q(n5598), .QN(
        n7156) );
  DFF_X1 \CACHE_MEM_reg[11][182]  ( .D(n13086), .CK(N28803), .Q(n5581), .QN(
        n7172) );
  DFF_X1 \CACHE_MEM_reg[11][181]  ( .D(n13085), .CK(N28803), .Q(n5570), .QN(
        n7188) );
  DFF_X1 \CACHE_MEM_reg[11][180]  ( .D(n13084), .CK(N28803), .Q(n5557), .QN(
        n7204) );
  DFF_X1 \CACHE_MEM_reg[11][179]  ( .D(n13083), .CK(N28803), .Q(n5542), .QN(
        n7220) );
  DFF_X1 \CACHE_MEM_reg[11][178]  ( .D(n13082), .CK(N28803), .Q(n5529), .QN(
        n7236) );
  DFF_X1 \CACHE_MEM_reg[11][177]  ( .D(n13081), .CK(N28803), .Q(n5518), .QN(
        n7252) );
  DFF_X1 \CACHE_MEM_reg[11][176]  ( .D(n13080), .CK(N28803), .Q(n5496), .QN(
        n7268) );
  DFF_X1 \CACHE_MEM_reg[11][175]  ( .D(n13079), .CK(N28803), .Q(n5485), .QN(
        n7284) );
  DFF_X1 \CACHE_MEM_reg[11][174]  ( .D(n13078), .CK(N28803), .Q(n5468), .QN(
        n7300) );
  DFF_X1 \CACHE_MEM_reg[11][173]  ( .D(n13077), .CK(N28803), .Q(n5457), .QN(
        n7316) );
  DFF_X1 \CACHE_MEM_reg[11][172]  ( .D(n13076), .CK(N28803), .Q(n5444), .QN(
        n7332) );
  DFF_X1 \CACHE_MEM_reg[11][171]  ( .D(n13075), .CK(N28803), .Q(n5429), .QN(
        n7348) );
  DFF_X1 \CACHE_MEM_reg[11][170]  ( .D(n13074), .CK(N28803), .Q(n5416), .QN(
        n7364) );
  DFF_X1 \CACHE_MEM_reg[11][169]  ( .D(n13073), .CK(N28803), .Q(n5405), .QN(
        n7380) );
  DFF_X1 \CACHE_MEM_reg[11][168]  ( .D(n13072), .CK(N28803), .Q(n5388), .QN(
        n7396) );
  DFF_X1 \CACHE_MEM_reg[11][167]  ( .D(n13071), .CK(N28803), .Q(n5377), .QN(
        n7412) );
  DFF_X1 \CACHE_MEM_reg[11][166]  ( .D(n13070), .CK(N28803), .Q(n5355), .QN(
        n7428) );
  DFF_X1 \CACHE_MEM_reg[11][165]  ( .D(n13069), .CK(N28803), .Q(n5344), .QN(
        n7444) );
  DFF_X1 \CACHE_MEM_reg[11][164]  ( .D(n13068), .CK(N28803), .Q(n5331), .QN(
        n7460) );
  DFF_X1 \CACHE_MEM_reg[11][163]  ( .D(n13067), .CK(N28803), .Q(n5316), .QN(
        n7476) );
  DFF_X1 \CACHE_MEM_reg[11][162]  ( .D(n13066), .CK(N28803), .Q(n5303), .QN(
        n7492) );
  DFF_X1 \CACHE_MEM_reg[11][161]  ( .D(n13065), .CK(N28803), .Q(n5292), .QN(
        n7508) );
  DFF_X1 \CACHE_MEM_reg[11][160]  ( .D(n13064), .CK(N28803), .Q(n5275), .QN(
        n7524) );
  DFF_X1 \CACHE_MEM_reg[11][159]  ( .D(n13063), .CK(N28803), .Q(n5714), .QN(
        n7540) );
  DFF_X1 \CACHE_MEM_reg[11][158]  ( .D(n13062), .CK(N28803), .Q(n5722), .QN(
        n7556) );
  DFF_X1 \CACHE_MEM_reg[11][157]  ( .D(n13061), .CK(N28803), .Q(n5686), .QN(
        n7572) );
  DFF_X1 \CACHE_MEM_reg[11][156]  ( .D(n13060), .CK(N28803), .Q(n5675), .QN(
        n7588) );
  DFF_X1 \CACHE_MEM_reg[11][155]  ( .D(n13059), .CK(N28803), .Q(n5653), .QN(
        n7604) );
  DFF_X1 \CACHE_MEM_reg[11][154]  ( .D(n13058), .CK(N28803), .Q(n5642), .QN(
        n7620) );
  DFF_X1 \CACHE_MEM_reg[11][153]  ( .D(n13057), .CK(N28803), .Q(n5629), .QN(
        n7636) );
  DFF_X1 \CACHE_MEM_reg[11][152]  ( .D(n13056), .CK(N28803), .Q(n5614), .QN(
        n7652) );
  DFF_X1 \CACHE_MEM_reg[11][151]  ( .D(n13055), .CK(N28803), .Q(n5601), .QN(
        n7668) );
  DFF_X1 \CACHE_MEM_reg[11][150]  ( .D(n13054), .CK(N28803), .Q(n5590), .QN(
        n7684) );
  DFF_X1 \CACHE_MEM_reg[11][149]  ( .D(n13053), .CK(N28803), .Q(n5573), .QN(
        n7700) );
  DFF_X1 \CACHE_MEM_reg[11][148]  ( .D(n13052), .CK(N28803), .Q(n5562), .QN(
        n7716) );
  DFF_X1 \CACHE_MEM_reg[11][147]  ( .D(n13051), .CK(N28803), .Q(n5545), .QN(
        n7732) );
  DFF_X1 \CACHE_MEM_reg[11][146]  ( .D(n13050), .CK(N28803), .Q(n5534), .QN(
        n7748) );
  DFF_X1 \CACHE_MEM_reg[11][145]  ( .D(n13049), .CK(N28803), .Q(n5521), .QN(
        n7764) );
  DFF_X1 \CACHE_MEM_reg[11][144]  ( .D(n13048), .CK(N28803), .Q(n5501), .QN(
        n7780) );
  DFF_X1 \CACHE_MEM_reg[11][143]  ( .D(n13047), .CK(N28803), .Q(n5488), .QN(
        n7796) );
  DFF_X1 \CACHE_MEM_reg[11][142]  ( .D(n13046), .CK(N28803), .Q(n5477), .QN(
        n7812) );
  DFF_X1 \CACHE_MEM_reg[11][141]  ( .D(n13045), .CK(N28803), .Q(n5460), .QN(
        n7828) );
  DFF_X1 \CACHE_MEM_reg[11][140]  ( .D(n13044), .CK(N28803), .Q(n5449), .QN(
        n7844) );
  DFF_X1 \CACHE_MEM_reg[11][139]  ( .D(n13043), .CK(N28803), .Q(n5432), .QN(
        n7860) );
  DFF_X1 \CACHE_MEM_reg[11][138]  ( .D(n13042), .CK(N28803), .Q(n5421), .QN(
        n7876) );
  DFF_X1 \CACHE_MEM_reg[11][137]  ( .D(n13041), .CK(N28803), .Q(n5408), .QN(
        n7892) );
  DFF_X1 \CACHE_MEM_reg[11][136]  ( .D(n13040), .CK(N28803), .Q(n5393), .QN(
        n7908) );
  DFF_X1 \CACHE_MEM_reg[11][135]  ( .D(n13039), .CK(N28803), .Q(n5380), .QN(
        n7924) );
  DFF_X1 \CACHE_MEM_reg[11][134]  ( .D(n13038), .CK(N28803), .Q(n5369), .QN(
        n7940) );
  DFF_X1 \CACHE_MEM_reg[11][133]  ( .D(n13037), .CK(N28803), .Q(n5347), .QN(
        n7956) );
  DFF_X1 \CACHE_MEM_reg[11][132]  ( .D(n13036), .CK(N28803), .Q(n5336), .QN(
        n7972) );
  DFF_X1 \CACHE_MEM_reg[11][131]  ( .D(n13035), .CK(N28803), .Q(n5319), .QN(
        n7988) );
  DFF_X1 \CACHE_MEM_reg[11][130]  ( .D(n13034), .CK(N28803), .Q(n5308), .QN(
        n8004) );
  DFF_X1 \CACHE_MEM_reg[11][129]  ( .D(n13033), .CK(N28803), .Q(n5295), .QN(
        n8020) );
  DFF_X1 \CACHE_MEM_reg[11][128]  ( .D(n13032), .CK(N28803), .Q(n5280), .QN(
        n8036) );
  DFF_X1 \CACHE_MEM_reg[11][127]  ( .D(n13031), .CK(N28803), .Q(n4373), .QN(
        n8052) );
  DFF_X1 \CACHE_MEM_reg[11][126]  ( .D(n13030), .CK(N28803), .Q(n4362), .QN(
        n8068) );
  DFF_X1 \CACHE_MEM_reg[11][125]  ( .D(n13029), .CK(N28803), .Q(n4342), .QN(
        n8084) );
  DFF_X1 \CACHE_MEM_reg[11][124]  ( .D(n13028), .CK(N28803), .Q(n4326), .QN(
        n8100) );
  DFF_X1 \CACHE_MEM_reg[11][123]  ( .D(n13027), .CK(N28803), .Q(n4301), .QN(
        n8116) );
  DFF_X1 \CACHE_MEM_reg[11][122]  ( .D(n13026), .CK(N28803), .Q(n4285), .QN(
        n8132) );
  DFF_X1 \CACHE_MEM_reg[11][121]  ( .D(n13025), .CK(N28803), .Q(n4265), .QN(
        n8148) );
  DFF_X1 \CACHE_MEM_reg[11][120]  ( .D(n13024), .CK(N28803), .Q(n4249), .QN(
        n8164) );
  DFF_X1 \CACHE_MEM_reg[11][119]  ( .D(n13023), .CK(N28803), .Q(n4229), .QN(
        n8180) );
  DFF_X1 \CACHE_MEM_reg[11][118]  ( .D(n13022), .CK(N28803), .Q(n4213), .QN(
        n8196) );
  DFF_X1 \CACHE_MEM_reg[11][117]  ( .D(n13021), .CK(N28803), .Q(n4193), .QN(
        n8212) );
  DFF_X1 \CACHE_MEM_reg[11][116]  ( .D(n13020), .CK(N28803), .Q(n4177), .QN(
        n8228) );
  DFF_X1 \CACHE_MEM_reg[11][115]  ( .D(n13019), .CK(N28803), .Q(n4152), .QN(
        n8244) );
  DFF_X1 \CACHE_MEM_reg[11][114]  ( .D(n13018), .CK(N28803), .Q(n4136), .QN(
        n8260) );
  DFF_X1 \CACHE_MEM_reg[11][113]  ( .D(n13017), .CK(N28803), .Q(n4116), .QN(
        n8276) );
  DFF_X1 \CACHE_MEM_reg[11][112]  ( .D(n13016), .CK(N28803), .Q(n4100), .QN(
        n8292) );
  DFF_X1 \CACHE_MEM_reg[11][111]  ( .D(n13015), .CK(N28803), .Q(n4080), .QN(
        n8308) );
  DFF_X1 \CACHE_MEM_reg[11][110]  ( .D(n13014), .CK(N28803), .Q(n4064), .QN(
        n8324) );
  DFF_X1 \CACHE_MEM_reg[11][109]  ( .D(n13013), .CK(N28803), .Q(n4044), .QN(
        n8340) );
  DFF_X1 \CACHE_MEM_reg[11][108]  ( .D(n13012), .CK(N28803), .Q(n4028), .QN(
        n8356) );
  DFF_X1 \CACHE_MEM_reg[11][107]  ( .D(n13011), .CK(N28803), .Q(n4003), .QN(
        n8372) );
  DFF_X1 \CACHE_MEM_reg[11][106]  ( .D(n13010), .CK(N28803), .Q(n3987), .QN(
        n8388) );
  DFF_X1 \CACHE_MEM_reg[11][105]  ( .D(n13009), .CK(N28803), .Q(n3967), .QN(
        n8404) );
  DFF_X1 \CACHE_MEM_reg[11][104]  ( .D(n13008), .CK(N28803), .Q(n3951), .QN(
        n8420) );
  DFF_X1 \CACHE_MEM_reg[11][103]  ( .D(n13007), .CK(N28803), .Q(n3931), .QN(
        n8436) );
  DFF_X1 \CACHE_MEM_reg[11][102]  ( .D(n13006), .CK(N28803), .Q(n3915), .QN(
        n8452) );
  DFF_X1 \CACHE_MEM_reg[11][101]  ( .D(n13005), .CK(N28803), .Q(n3895), .QN(
        n8468) );
  DFF_X1 \CACHE_MEM_reg[11][100]  ( .D(n13004), .CK(N28803), .Q(n3879), .QN(
        n8484) );
  DFF_X1 \CACHE_MEM_reg[11][99]  ( .D(n13003), .CK(N28803), .Q(n3854), .QN(
        n8500) );
  DFF_X1 \CACHE_MEM_reg[11][98]  ( .D(n13002), .CK(N28803), .Q(n3838), .QN(
        n8516) );
  DFF_X1 \CACHE_MEM_reg[11][97]  ( .D(n13001), .CK(N28803), .Q(n3818), .QN(
        n8532) );
  DFF_X1 \CACHE_MEM_reg[11][96]  ( .D(n13000), .CK(N28803), .Q(n3802), .QN(
        n8548) );
  DFF_X1 \CACHE_MEM_reg[11][95]  ( .D(n12999), .CK(N28803), .Q(n4378), .QN(
        n8564) );
  DFF_X1 \CACHE_MEM_reg[11][94]  ( .D(n12998), .CK(N28803), .Q(n4365), .QN(
        n8580) );
  DFF_X1 \CACHE_MEM_reg[11][93]  ( .D(n12997), .CK(N28803), .Q(n4345), .QN(
        n8596) );
  DFF_X1 \CACHE_MEM_reg[11][92]  ( .D(n12996), .CK(N28803), .Q(n4329), .QN(
        n8612) );
  DFF_X1 \CACHE_MEM_reg[11][91]  ( .D(n12995), .CK(N28803), .Q(n4304), .QN(
        n8628) );
  DFF_X1 \CACHE_MEM_reg[11][90]  ( .D(n12994), .CK(N28803), .Q(n4288), .QN(
        n8644) );
  DFF_X1 \CACHE_MEM_reg[11][89]  ( .D(n12993), .CK(N28803), .Q(n4268), .QN(
        n8660) );
  DFF_X1 \CACHE_MEM_reg[11][88]  ( .D(n12992), .CK(N28803), .Q(n4252), .QN(
        n8676) );
  DFF_X1 \CACHE_MEM_reg[11][87]  ( .D(n12991), .CK(N28803), .Q(n4232), .QN(
        n8692) );
  DFF_X1 \CACHE_MEM_reg[11][86]  ( .D(n12990), .CK(N28803), .Q(n4216), .QN(
        n8708) );
  DFF_X1 \CACHE_MEM_reg[11][85]  ( .D(n12989), .CK(N28803), .Q(n4196), .QN(
        n8724) );
  DFF_X1 \CACHE_MEM_reg[11][84]  ( .D(n12988), .CK(N28803), .Q(n4180), .QN(
        n8740) );
  DFF_X1 \CACHE_MEM_reg[11][83]  ( .D(n12987), .CK(N28803), .Q(n4155), .QN(
        n8756) );
  DFF_X1 \CACHE_MEM_reg[11][82]  ( .D(n12986), .CK(N28803), .Q(n4139), .QN(
        n8772) );
  DFF_X1 \CACHE_MEM_reg[11][81]  ( .D(n12985), .CK(N28803), .Q(n4119), .QN(
        n8788) );
  DFF_X1 \CACHE_MEM_reg[11][80]  ( .D(n12984), .CK(N28803), .Q(n4103), .QN(
        n8804) );
  DFF_X1 \CACHE_MEM_reg[11][79]  ( .D(n12983), .CK(N28803), .Q(n4083), .QN(
        n8820) );
  DFF_X1 \CACHE_MEM_reg[11][78]  ( .D(n12982), .CK(N28803), .Q(n4067), .QN(
        n8836) );
  DFF_X1 \CACHE_MEM_reg[11][77]  ( .D(n12981), .CK(N28803), .Q(n4047), .QN(
        n8852) );
  DFF_X1 \CACHE_MEM_reg[11][76]  ( .D(n12980), .CK(N28803), .Q(n4031), .QN(
        n8868) );
  DFF_X1 \CACHE_MEM_reg[11][75]  ( .D(n12979), .CK(N28803), .Q(n4006), .QN(
        n8884) );
  DFF_X1 \CACHE_MEM_reg[11][74]  ( .D(n12978), .CK(N28803), .Q(n3990), .QN(
        n8900) );
  DFF_X1 \CACHE_MEM_reg[11][73]  ( .D(n12977), .CK(N28803), .Q(n3970), .QN(
        n8916) );
  DFF_X1 \CACHE_MEM_reg[11][72]  ( .D(n12976), .CK(N28803), .Q(n3954), .QN(
        n8932) );
  DFF_X1 \CACHE_MEM_reg[11][71]  ( .D(n12975), .CK(N28803), .Q(n3934), .QN(
        n8948) );
  DFF_X1 \CACHE_MEM_reg[11][70]  ( .D(n12974), .CK(N28803), .Q(n3918), .QN(
        n8964) );
  DFF_X1 \CACHE_MEM_reg[11][69]  ( .D(n12973), .CK(N28803), .Q(n3898), .QN(
        n8980) );
  DFF_X1 \CACHE_MEM_reg[11][68]  ( .D(n12972), .CK(N28803), .Q(n3882), .QN(
        n8996) );
  DFF_X1 \CACHE_MEM_reg[11][67]  ( .D(n12971), .CK(N28803), .Q(n3857), .QN(
        n9012) );
  DFF_X1 \CACHE_MEM_reg[11][66]  ( .D(n12970), .CK(N28803), .Q(n3841), .QN(
        n9028) );
  DFF_X1 \CACHE_MEM_reg[11][65]  ( .D(n12969), .CK(N28803), .Q(n3821), .QN(
        n9044) );
  DFF_X1 \CACHE_MEM_reg[11][64]  ( .D(n12968), .CK(N28803), .Q(n3805), .QN(
        n9060) );
  DFF_X1 \CACHE_MEM_reg[11][63]  ( .D(n12967), .CK(N28803), .Q(n4820), .QN(
        n9076) );
  DFF_X1 \CACHE_MEM_reg[11][62]  ( .D(n12966), .CK(N28803), .Q(n4809), .QN(
        n9092) );
  DFF_X1 \CACHE_MEM_reg[11][61]  ( .D(n12965), .CK(N28803), .Q(n4792), .QN(
        n9108) );
  DFF_X1 \CACHE_MEM_reg[11][60]  ( .D(n12964), .CK(N28803), .Q(n4781), .QN(
        n9124) );
  DFF_X1 \CACHE_MEM_reg[11][59]  ( .D(n12963), .CK(N28803), .Q(n4759), .QN(
        n9140) );
  DFF_X1 \CACHE_MEM_reg[11][58]  ( .D(n12962), .CK(N28803), .Q(n4748), .QN(
        n9156) );
  DFF_X1 \CACHE_MEM_reg[11][57]  ( .D(n12961), .CK(N28803), .Q(n4735), .QN(
        n9172) );
  DFF_X1 \CACHE_MEM_reg[11][56]  ( .D(n12960), .CK(N28803), .Q(n4720), .QN(
        n9188) );
  DFF_X1 \CACHE_MEM_reg[11][55]  ( .D(n12959), .CK(N28803), .Q(n4707), .QN(
        n9204) );
  DFF_X1 \CACHE_MEM_reg[11][54]  ( .D(n12958), .CK(N28803), .Q(n4696), .QN(
        n9220) );
  DFF_X1 \CACHE_MEM_reg[11][53]  ( .D(n12957), .CK(N28803), .Q(n4679), .QN(
        n9236) );
  DFF_X1 \CACHE_MEM_reg[11][52]  ( .D(n12956), .CK(N28803), .Q(n4668), .QN(
        n9252) );
  DFF_X1 \CACHE_MEM_reg[11][51]  ( .D(n12955), .CK(N28803), .Q(n4651), .QN(
        n9268) );
  DFF_X1 \CACHE_MEM_reg[11][50]  ( .D(n12954), .CK(N28803), .Q(n4640), .QN(
        n9284) );
  DFF_X1 \CACHE_MEM_reg[11][49]  ( .D(n12953), .CK(N28803), .Q(n4627), .QN(
        n9300) );
  DFF_X1 \CACHE_MEM_reg[11][48]  ( .D(n12952), .CK(N28803), .Q(n4607), .QN(
        n9316) );
  DFF_X1 \CACHE_MEM_reg[11][47]  ( .D(n12951), .CK(N28803), .Q(n4594), .QN(
        n9332) );
  DFF_X1 \CACHE_MEM_reg[11][46]  ( .D(n12950), .CK(N28803), .Q(n4583), .QN(
        n9348) );
  DFF_X1 \CACHE_MEM_reg[11][45]  ( .D(n12949), .CK(N28803), .Q(n4566), .QN(
        n9364) );
  DFF_X1 \CACHE_MEM_reg[11][44]  ( .D(n12948), .CK(N28803), .Q(n4555), .QN(
        n9380) );
  DFF_X1 \CACHE_MEM_reg[11][43]  ( .D(n12947), .CK(N28803), .Q(n4538), .QN(
        n9396) );
  DFF_X1 \CACHE_MEM_reg[11][42]  ( .D(n12946), .CK(N28803), .Q(n4527), .QN(
        n9412) );
  DFF_X1 \CACHE_MEM_reg[11][41]  ( .D(n12945), .CK(N28803), .Q(n4514), .QN(
        n9428) );
  DFF_X1 \CACHE_MEM_reg[11][40]  ( .D(n12944), .CK(N28803), .Q(n4499), .QN(
        n9444) );
  DFF_X1 \CACHE_MEM_reg[11][39]  ( .D(n12943), .CK(N28803), .Q(n4486), .QN(
        n9460) );
  DFF_X1 \CACHE_MEM_reg[11][38]  ( .D(n12942), .CK(N28803), .Q(n4475), .QN(
        n9476) );
  DFF_X1 \CACHE_MEM_reg[11][37]  ( .D(n12941), .CK(N28803), .Q(n4453), .QN(
        n9492) );
  DFF_X1 \CACHE_MEM_reg[11][36]  ( .D(n12940), .CK(N28803), .Q(n4442), .QN(
        n9508) );
  DFF_X1 \CACHE_MEM_reg[11][35]  ( .D(n12939), .CK(N28803), .Q(n4425), .QN(
        n9524) );
  DFF_X1 \CACHE_MEM_reg[11][34]  ( .D(n12938), .CK(N28803), .Q(n4414), .QN(
        n9540) );
  DFF_X1 \CACHE_MEM_reg[11][33]  ( .D(n12937), .CK(N28803), .Q(n4401), .QN(
        n9556) );
  DFF_X1 \CACHE_MEM_reg[11][32]  ( .D(n12936), .CK(N28803), .Q(n4386), .QN(
        n9572) );
  DFF_X1 \CACHE_MEM_reg[11][31]  ( .D(n12935), .CK(N28803), .Q(n4825), .QN(
        n9588) );
  DFF_X1 \CACHE_MEM_reg[11][30]  ( .D(n12934), .CK(N28803), .Q(n4812), .QN(
        n9604) );
  DFF_X1 \CACHE_MEM_reg[11][29]  ( .D(n12933), .CK(N28803), .Q(n4797), .QN(
        n9620) );
  DFF_X1 \CACHE_MEM_reg[11][28]  ( .D(n12932), .CK(N28803), .Q(n4784), .QN(
        n9636) );
  DFF_X1 \CACHE_MEM_reg[11][27]  ( .D(n12931), .CK(N28803), .Q(n4773), .QN(
        n9652) );
  DFF_X1 \CACHE_MEM_reg[11][26]  ( .D(n12930), .CK(N28803), .Q(n4751), .QN(
        n9668) );
  DFF_X1 \CACHE_MEM_reg[11][25]  ( .D(n12929), .CK(N28803), .Q(n4740), .QN(
        n9684) );
  DFF_X1 \CACHE_MEM_reg[11][24]  ( .D(n12928), .CK(N28803), .Q(n4723), .QN(
        n9700) );
  DFF_X1 \CACHE_MEM_reg[11][23]  ( .D(n12927), .CK(N28803), .Q(n4712), .QN(
        n9716) );
  DFF_X1 \CACHE_MEM_reg[11][22]  ( .D(n12926), .CK(N28803), .Q(n4699), .QN(
        n9732) );
  DFF_X1 \CACHE_MEM_reg[11][21]  ( .D(n12925), .CK(N28803), .Q(n4684), .QN(
        n9748) );
  DFF_X1 \CACHE_MEM_reg[11][20]  ( .D(n12924), .CK(N28803), .Q(n4671), .QN(
        n9764) );
  DFF_X1 \CACHE_MEM_reg[11][19]  ( .D(n12923), .CK(N28803), .Q(n4660), .QN(
        n9780) );
  DFF_X1 \CACHE_MEM_reg[11][18]  ( .D(n12922), .CK(N28803), .Q(n4643), .QN(
        n9796) );
  DFF_X1 \CACHE_MEM_reg[11][17]  ( .D(n12921), .CK(N28803), .Q(n4632), .QN(
        n9812) );
  DFF_X1 \CACHE_MEM_reg[11][16]  ( .D(n12920), .CK(N28803), .Q(n4610), .QN(
        n9828) );
  DFF_X1 \CACHE_MEM_reg[11][15]  ( .D(n12919), .CK(N28803), .Q(n4599), .QN(
        n9844) );
  DFF_X1 \CACHE_MEM_reg[11][14]  ( .D(n12918), .CK(N28803), .Q(n4586), .QN(
        n9860) );
  DFF_X1 \CACHE_MEM_reg[11][13]  ( .D(n12917), .CK(N28803), .Q(n4571), .QN(
        n9876) );
  DFF_X1 \CACHE_MEM_reg[11][12]  ( .D(n12916), .CK(N28803), .Q(n4558), .QN(
        n9892) );
  DFF_X1 \CACHE_MEM_reg[11][11]  ( .D(n12915), .CK(N28803), .Q(n4547), .QN(
        n9908) );
  DFF_X1 \CACHE_MEM_reg[11][10]  ( .D(n12914), .CK(N28803), .Q(n4530), .QN(
        n9924) );
  DFF_X1 \CACHE_MEM_reg[11][9]  ( .D(n12913), .CK(N28803), .Q(n4519), .QN(
        n9940) );
  DFF_X1 \CACHE_MEM_reg[11][8]  ( .D(n12912), .CK(N28803), .Q(n4502), .QN(
        n9956) );
  DFF_X1 \CACHE_MEM_reg[11][7]  ( .D(n12911), .CK(N28803), .Q(n4491), .QN(
        n9972) );
  DFF_X1 \CACHE_MEM_reg[11][6]  ( .D(n12910), .CK(N28803), .Q(n4478), .QN(
        n9988) );
  DFF_X1 \CACHE_MEM_reg[11][5]  ( .D(n12909), .CK(N28803), .Q(n4458), .QN(
        n10004) );
  DFF_X1 \CACHE_MEM_reg[11][4]  ( .D(n12908), .CK(N28803), .Q(n4445), .QN(
        n10020) );
  DFF_X1 \CACHE_MEM_reg[11][3]  ( .D(n12907), .CK(N28803), .Q(n4434), .QN(
        n10036) );
  DFF_X1 \CACHE_MEM_reg[11][2]  ( .D(n12906), .CK(N28803), .Q(n4417), .QN(
        n10052) );
  DFF_X1 \CACHE_MEM_reg[11][1]  ( .D(n12905), .CK(N28803), .Q(n4406), .QN(
        n10068) );
  DFF_X1 \CACHE_MEM_reg[11][0]  ( .D(n12904), .CK(N28803), .Q(n4389), .QN(
        n10084) );
  DFF_X1 \CACHE_MEM_reg[10][255]  ( .D(n12903), .CK(N28803), .Q(n2880), .QN(
        n6000) );
  DFF_X1 \CACHE_MEM_reg[10][254]  ( .D(n12902), .CK(N28803), .Q(n2863), .QN(
        n6016) );
  DFF_X1 \CACHE_MEM_reg[10][253]  ( .D(n12901), .CK(N28803), .Q(n2852), .QN(
        n6032) );
  DFF_X1 \CACHE_MEM_reg[10][252]  ( .D(n12900), .CK(N28803), .Q(n2839), .QN(
        n6048) );
  DFF_X1 \CACHE_MEM_reg[10][251]  ( .D(n12899), .CK(N28803), .Q(n2819), .QN(
        n6064) );
  DFF_X1 \CACHE_MEM_reg[10][250]  ( .D(n12898), .CK(N28803), .Q(n2806), .QN(
        n6080) );
  DFF_X1 \CACHE_MEM_reg[10][249]  ( .D(n12897), .CK(N28803), .Q(n2795), .QN(
        n6096) );
  DFF_X1 \CACHE_MEM_reg[10][248]  ( .D(n12896), .CK(N28803), .Q(n2778), .QN(
        n6112) );
  DFF_X1 \CACHE_MEM_reg[10][247]  ( .D(n12895), .CK(N28803), .Q(n2767), .QN(
        n6128) );
  DFF_X1 \CACHE_MEM_reg[10][246]  ( .D(n12894), .CK(N28803), .Q(n2750), .QN(
        n6144) );
  DFF_X1 \CACHE_MEM_reg[10][245]  ( .D(n12893), .CK(N28803), .Q(n2739), .QN(
        n6160) );
  DFF_X1 \CACHE_MEM_reg[10][244]  ( .D(n12892), .CK(N28803), .Q(n2726), .QN(
        n6176) );
  DFF_X1 \CACHE_MEM_reg[10][243]  ( .D(n12891), .CK(N28803), .Q(n2711), .QN(
        n6192) );
  DFF_X1 \CACHE_MEM_reg[10][242]  ( .D(n12890), .CK(N28803), .Q(n2698), .QN(
        n6208) );
  DFF_X1 \CACHE_MEM_reg[10][241]  ( .D(n12889), .CK(N28803), .Q(n2687), .QN(
        n6224) );
  DFF_X1 \CACHE_MEM_reg[10][240]  ( .D(n12888), .CK(N28803), .Q(n3335), .QN(
        n6240) );
  DFF_X1 \CACHE_MEM_reg[10][239]  ( .D(n12887), .CK(N28803), .Q(n2657), .QN(
        n6256) );
  DFF_X1 \CACHE_MEM_reg[10][238]  ( .D(n12886), .CK(N28803), .Q(n2646), .QN(
        n6272) );
  DFF_X1 \CACHE_MEM_reg[10][237]  ( .D(n12885), .CK(N28803), .Q(n2629), .QN(
        n6288) );
  DFF_X1 \CACHE_MEM_reg[10][236]  ( .D(n12884), .CK(N28803), .Q(n2618), .QN(
        n6304) );
  DFF_X1 \CACHE_MEM_reg[10][235]  ( .D(n12883), .CK(N28803), .Q(n2601), .QN(
        n6320) );
  DFF_X1 \CACHE_MEM_reg[10][234]  ( .D(n12882), .CK(N28803), .Q(n2590), .QN(
        n6336) );
  DFF_X1 \CACHE_MEM_reg[10][233]  ( .D(n12881), .CK(N28803), .Q(n2577), .QN(
        n6352) );
  DFF_X1 \CACHE_MEM_reg[10][232]  ( .D(n12880), .CK(N28803), .Q(n2562), .QN(
        n6368) );
  DFF_X1 \CACHE_MEM_reg[10][231]  ( .D(n12879), .CK(N28803), .Q(n2549), .QN(
        n6384) );
  DFF_X1 \CACHE_MEM_reg[10][230]  ( .D(n12878), .CK(N28803), .Q(n2538), .QN(
        n6400) );
  DFF_X1 \CACHE_MEM_reg[10][229]  ( .D(n12877), .CK(N28803), .Q(n2516), .QN(
        n6416) );
  DFF_X1 \CACHE_MEM_reg[10][228]  ( .D(n12876), .CK(N28803), .Q(n2505), .QN(
        n6432) );
  DFF_X1 \CACHE_MEM_reg[10][227]  ( .D(n12875), .CK(N28803), .Q(n2488), .QN(
        n6448) );
  DFF_X1 \CACHE_MEM_reg[10][226]  ( .D(n12874), .CK(N28803), .Q(n2477), .QN(
        n6464) );
  DFF_X1 \CACHE_MEM_reg[10][225]  ( .D(n12873), .CK(N28803), .Q(n2464), .QN(
        n6480) );
  DFF_X1 \CACHE_MEM_reg[10][224]  ( .D(n12872), .CK(N28803), .Q(n2449), .QN(
        n6496) );
  DFF_X1 \CACHE_MEM_reg[10][223]  ( .D(n12871), .CK(N28803), .Q(n2883), .QN(
        n6512) );
  DFF_X1 \CACHE_MEM_reg[10][222]  ( .D(n12870), .CK(N28803), .Q(n2872), .QN(
        n6528) );
  DFF_X1 \CACHE_MEM_reg[10][221]  ( .D(n12869), .CK(N28803), .Q(n2855), .QN(
        n6544) );
  DFF_X1 \CACHE_MEM_reg[10][220]  ( .D(n12868), .CK(N28803), .Q(n2844), .QN(
        n6560) );
  DFF_X1 \CACHE_MEM_reg[10][219]  ( .D(n12867), .CK(N28803), .Q(n2822), .QN(
        n6576) );
  DFF_X1 \CACHE_MEM_reg[10][218]  ( .D(n12866), .CK(N28803), .Q(n2811), .QN(
        n6592) );
  DFF_X1 \CACHE_MEM_reg[10][217]  ( .D(n12865), .CK(N28803), .Q(n2798), .QN(
        n6608) );
  DFF_X1 \CACHE_MEM_reg[10][216]  ( .D(n12864), .CK(N28803), .Q(n2783), .QN(
        n6624) );
  DFF_X1 \CACHE_MEM_reg[10][215]  ( .D(n12863), .CK(N28803), .Q(n2770), .QN(
        n6640) );
  DFF_X1 \CACHE_MEM_reg[10][214]  ( .D(n12862), .CK(N28803), .Q(n2759), .QN(
        n6656) );
  DFF_X1 \CACHE_MEM_reg[10][213]  ( .D(n12861), .CK(N28803), .Q(n2742), .QN(
        n6672) );
  DFF_X1 \CACHE_MEM_reg[10][212]  ( .D(n12860), .CK(N28803), .Q(n2731), .QN(
        n6688) );
  DFF_X1 \CACHE_MEM_reg[10][211]  ( .D(n12859), .CK(N28803), .Q(n2714), .QN(
        n6704) );
  DFF_X1 \CACHE_MEM_reg[10][210]  ( .D(n12858), .CK(N28803), .Q(n2703), .QN(
        n6720) );
  DFF_X1 \CACHE_MEM_reg[10][209]  ( .D(n12857), .CK(N28803), .Q(n2690), .QN(
        n6736) );
  DFF_X1 \CACHE_MEM_reg[10][208]  ( .D(n12856), .CK(N28803), .Q(n2670), .QN(
        n6752) );
  DFF_X1 \CACHE_MEM_reg[10][207]  ( .D(n12855), .CK(N28803), .Q(n2662), .QN(
        n6768) );
  DFF_X1 \CACHE_MEM_reg[10][206]  ( .D(n12854), .CK(N28803), .Q(n2649), .QN(
        n6784) );
  DFF_X1 \CACHE_MEM_reg[10][205]  ( .D(n12853), .CK(N28803), .Q(n2634), .QN(
        n6800) );
  DFF_X1 \CACHE_MEM_reg[10][204]  ( .D(n12852), .CK(N28803), .Q(n2621), .QN(
        n6816) );
  DFF_X1 \CACHE_MEM_reg[10][203]  ( .D(n12851), .CK(N28803), .Q(n2610), .QN(
        n6832) );
  DFF_X1 \CACHE_MEM_reg[10][202]  ( .D(n12850), .CK(N28803), .Q(n2593), .QN(
        n6848) );
  DFF_X1 \CACHE_MEM_reg[10][201]  ( .D(n12849), .CK(N28803), .Q(n2582), .QN(
        n6864) );
  DFF_X1 \CACHE_MEM_reg[10][200]  ( .D(n12848), .CK(N28803), .Q(n2565), .QN(
        n6880) );
  DFF_X1 \CACHE_MEM_reg[10][199]  ( .D(n12847), .CK(N28803), .Q(n2554), .QN(
        n6896) );
  DFF_X1 \CACHE_MEM_reg[10][198]  ( .D(n12846), .CK(N28803), .Q(n2541), .QN(
        n6912) );
  DFF_X1 \CACHE_MEM_reg[10][197]  ( .D(n12845), .CK(N28803), .Q(n2521), .QN(
        n6928) );
  DFF_X1 \CACHE_MEM_reg[10][196]  ( .D(n12844), .CK(N28803), .Q(n2508), .QN(
        n6944) );
  DFF_X1 \CACHE_MEM_reg[10][195]  ( .D(n12843), .CK(N28803), .Q(n2497), .QN(
        n6960) );
  DFF_X1 \CACHE_MEM_reg[10][194]  ( .D(n12842), .CK(N28803), .Q(n2480), .QN(
        n6976) );
  DFF_X1 \CACHE_MEM_reg[10][193]  ( .D(n12841), .CK(N28803), .Q(n2469), .QN(
        n6992) );
  DFF_X1 \CACHE_MEM_reg[10][192]  ( .D(n12840), .CK(N28803), .Q(n2452), .QN(
        n7008) );
  DFF_X1 \CACHE_MEM_reg[10][191]  ( .D(n12839), .CK(N28803), .Q(n3327), .QN(
        n7024) );
  DFF_X1 \CACHE_MEM_reg[10][190]  ( .D(n12838), .CK(N28803), .Q(n3310), .QN(
        n7040) );
  DFF_X1 \CACHE_MEM_reg[10][189]  ( .D(n12837), .CK(N28803), .Q(n3299), .QN(
        n7056) );
  DFF_X1 \CACHE_MEM_reg[10][188]  ( .D(n12836), .CK(N28803), .Q(n3286), .QN(
        n7072) );
  DFF_X1 \CACHE_MEM_reg[10][187]  ( .D(n12835), .CK(N28803), .Q(n3266), .QN(
        n7088) );
  DFF_X1 \CACHE_MEM_reg[10][186]  ( .D(n12834), .CK(N28803), .Q(n3253), .QN(
        n7104) );
  DFF_X1 \CACHE_MEM_reg[10][185]  ( .D(n12833), .CK(N28803), .Q(n3242), .QN(
        n7120) );
  DFF_X1 \CACHE_MEM_reg[10][184]  ( .D(n12832), .CK(N28803), .Q(n3225), .QN(
        n7136) );
  DFF_X1 \CACHE_MEM_reg[10][183]  ( .D(n12831), .CK(N28803), .Q(n3214), .QN(
        n7152) );
  DFF_X1 \CACHE_MEM_reg[10][182]  ( .D(n12830), .CK(N28803), .Q(n3197), .QN(
        n7168) );
  DFF_X1 \CACHE_MEM_reg[10][181]  ( .D(n12829), .CK(N28803), .Q(n3186), .QN(
        n7184) );
  DFF_X1 \CACHE_MEM_reg[10][180]  ( .D(n12828), .CK(N28803), .Q(n3173), .QN(
        n7200) );
  DFF_X1 \CACHE_MEM_reg[10][179]  ( .D(n12827), .CK(N28803), .Q(n3158), .QN(
        n7216) );
  DFF_X1 \CACHE_MEM_reg[10][178]  ( .D(n12826), .CK(N28803), .Q(n3145), .QN(
        n7232) );
  DFF_X1 \CACHE_MEM_reg[10][177]  ( .D(n12825), .CK(N28803), .Q(n3134), .QN(
        n7248) );
  DFF_X1 \CACHE_MEM_reg[10][176]  ( .D(n12824), .CK(N28803), .Q(n3112), .QN(
        n7264) );
  DFF_X1 \CACHE_MEM_reg[10][175]  ( .D(n12823), .CK(N28803), .Q(n3101), .QN(
        n7280) );
  DFF_X1 \CACHE_MEM_reg[10][174]  ( .D(n12822), .CK(N28803), .Q(n3084), .QN(
        n7296) );
  DFF_X1 \CACHE_MEM_reg[10][173]  ( .D(n12821), .CK(N28803), .Q(n3073), .QN(
        n7312) );
  DFF_X1 \CACHE_MEM_reg[10][172]  ( .D(n12820), .CK(N28803), .Q(n3060), .QN(
        n7328) );
  DFF_X1 \CACHE_MEM_reg[10][171]  ( .D(n12819), .CK(N28803), .Q(n3045), .QN(
        n7344) );
  DFF_X1 \CACHE_MEM_reg[10][170]  ( .D(n12818), .CK(N28803), .Q(n3032), .QN(
        n7360) );
  DFF_X1 \CACHE_MEM_reg[10][169]  ( .D(n12817), .CK(N28803), .Q(n3021), .QN(
        n7376) );
  DFF_X1 \CACHE_MEM_reg[10][168]  ( .D(n12816), .CK(N28803), .Q(n3004), .QN(
        n7392) );
  DFF_X1 \CACHE_MEM_reg[10][167]  ( .D(n12815), .CK(N28803), .Q(n2993), .QN(
        n7408) );
  DFF_X1 \CACHE_MEM_reg[10][166]  ( .D(n12814), .CK(N28803), .Q(n2971), .QN(
        n7424) );
  DFF_X1 \CACHE_MEM_reg[10][165]  ( .D(n12813), .CK(N28803), .Q(n2960), .QN(
        n7440) );
  DFF_X1 \CACHE_MEM_reg[10][164]  ( .D(n12812), .CK(N28803), .Q(n2947), .QN(
        n7456) );
  DFF_X1 \CACHE_MEM_reg[10][163]  ( .D(n12811), .CK(N28803), .Q(n2932), .QN(
        n7472) );
  DFF_X1 \CACHE_MEM_reg[10][162]  ( .D(n12810), .CK(N28803), .Q(n2919), .QN(
        n7488) );
  DFF_X1 \CACHE_MEM_reg[10][161]  ( .D(n12809), .CK(N28803), .Q(n2908), .QN(
        n7504) );
  DFF_X1 \CACHE_MEM_reg[10][160]  ( .D(n12808), .CK(N28803), .Q(n2891), .QN(
        n7520) );
  DFF_X1 \CACHE_MEM_reg[10][159]  ( .D(n12807), .CK(N28803), .Q(n3330), .QN(
        n7536) );
  DFF_X1 \CACHE_MEM_reg[10][158]  ( .D(n12806), .CK(N28803), .Q(n3338), .QN(
        n7552) );
  DFF_X1 \CACHE_MEM_reg[10][157]  ( .D(n12805), .CK(N28803), .Q(n3302), .QN(
        n7568) );
  DFF_X1 \CACHE_MEM_reg[10][156]  ( .D(n12804), .CK(N28803), .Q(n3291), .QN(
        n7584) );
  DFF_X1 \CACHE_MEM_reg[10][155]  ( .D(n12803), .CK(N28803), .Q(n3269), .QN(
        n7600) );
  DFF_X1 \CACHE_MEM_reg[10][154]  ( .D(n12802), .CK(N28803), .Q(n3258), .QN(
        n7616) );
  DFF_X1 \CACHE_MEM_reg[10][153]  ( .D(n12801), .CK(N28803), .Q(n3245), .QN(
        n7632) );
  DFF_X1 \CACHE_MEM_reg[10][152]  ( .D(n12800), .CK(N28803), .Q(n3230), .QN(
        n7648) );
  DFF_X1 \CACHE_MEM_reg[10][151]  ( .D(n12799), .CK(N28803), .Q(n3217), .QN(
        n7664) );
  DFF_X1 \CACHE_MEM_reg[10][150]  ( .D(n12798), .CK(N28803), .Q(n3206), .QN(
        n7680) );
  DFF_X1 \CACHE_MEM_reg[10][149]  ( .D(n12797), .CK(N28803), .Q(n3189), .QN(
        n7696) );
  DFF_X1 \CACHE_MEM_reg[10][148]  ( .D(n12796), .CK(N28803), .Q(n3178), .QN(
        n7712) );
  DFF_X1 \CACHE_MEM_reg[10][147]  ( .D(n12795), .CK(N28803), .Q(n3161), .QN(
        n7728) );
  DFF_X1 \CACHE_MEM_reg[10][146]  ( .D(n12794), .CK(N28803), .Q(n3150), .QN(
        n7744) );
  DFF_X1 \CACHE_MEM_reg[10][145]  ( .D(n12793), .CK(N28803), .Q(n3137), .QN(
        n7760) );
  DFF_X1 \CACHE_MEM_reg[10][144]  ( .D(n12792), .CK(N28803), .Q(n3117), .QN(
        n7776) );
  DFF_X1 \CACHE_MEM_reg[10][143]  ( .D(n12791), .CK(N28803), .Q(n3104), .QN(
        n7792) );
  DFF_X1 \CACHE_MEM_reg[10][142]  ( .D(n12790), .CK(N28803), .Q(n3093), .QN(
        n7808) );
  DFF_X1 \CACHE_MEM_reg[10][141]  ( .D(n12789), .CK(N28803), .Q(n3076), .QN(
        n7824) );
  DFF_X1 \CACHE_MEM_reg[10][140]  ( .D(n12788), .CK(N28803), .Q(n3065), .QN(
        n7840) );
  DFF_X1 \CACHE_MEM_reg[10][139]  ( .D(n12787), .CK(N28803), .Q(n3048), .QN(
        n7856) );
  DFF_X1 \CACHE_MEM_reg[10][138]  ( .D(n12786), .CK(N28803), .Q(n3037), .QN(
        n7872) );
  DFF_X1 \CACHE_MEM_reg[10][137]  ( .D(n12785), .CK(N28803), .Q(n3024), .QN(
        n7888) );
  DFF_X1 \CACHE_MEM_reg[10][136]  ( .D(n12784), .CK(N28803), .Q(n3009), .QN(
        n7904) );
  DFF_X1 \CACHE_MEM_reg[10][135]  ( .D(n12783), .CK(N28803), .Q(n2996), .QN(
        n7920) );
  DFF_X1 \CACHE_MEM_reg[10][134]  ( .D(n12782), .CK(N28803), .Q(n2985), .QN(
        n7936) );
  DFF_X1 \CACHE_MEM_reg[10][133]  ( .D(n12781), .CK(N28803), .Q(n2963), .QN(
        n7952) );
  DFF_X1 \CACHE_MEM_reg[10][132]  ( .D(n12780), .CK(N28803), .Q(n2952), .QN(
        n7968) );
  DFF_X1 \CACHE_MEM_reg[10][131]  ( .D(n12779), .CK(N28803), .Q(n2935), .QN(
        n7984) );
  DFF_X1 \CACHE_MEM_reg[10][130]  ( .D(n12778), .CK(N28803), .Q(n2924), .QN(
        n8000) );
  DFF_X1 \CACHE_MEM_reg[10][129]  ( .D(n12777), .CK(N28803), .Q(n2911), .QN(
        n8016) );
  DFF_X1 \CACHE_MEM_reg[10][128]  ( .D(n12776), .CK(N28803), .Q(n2896), .QN(
        n8032) );
  DFF_X1 \CACHE_MEM_reg[10][127]  ( .D(n12775), .CK(N28803), .Q(n1989), .QN(
        n8048) );
  DFF_X1 \CACHE_MEM_reg[10][126]  ( .D(n12774), .CK(N28803), .Q(n1978), .QN(
        n8064) );
  DFF_X1 \CACHE_MEM_reg[10][125]  ( .D(n12773), .CK(N28803), .Q(n1958), .QN(
        n8080) );
  DFF_X1 \CACHE_MEM_reg[10][124]  ( .D(n12772), .CK(N28803), .Q(n1942), .QN(
        n8096) );
  DFF_X1 \CACHE_MEM_reg[10][123]  ( .D(n12771), .CK(N28803), .Q(n1917), .QN(
        n8112) );
  DFF_X1 \CACHE_MEM_reg[10][122]  ( .D(n12770), .CK(N28803), .Q(n1901), .QN(
        n8128) );
  DFF_X1 \CACHE_MEM_reg[10][121]  ( .D(n12769), .CK(N28803), .Q(n1881), .QN(
        n8144) );
  DFF_X1 \CACHE_MEM_reg[10][120]  ( .D(n12768), .CK(N28803), .Q(n1865), .QN(
        n8160) );
  DFF_X1 \CACHE_MEM_reg[10][119]  ( .D(n12767), .CK(N28803), .Q(n1845), .QN(
        n8176) );
  DFF_X1 \CACHE_MEM_reg[10][118]  ( .D(n12766), .CK(N28803), .Q(n1829), .QN(
        n8192) );
  DFF_X1 \CACHE_MEM_reg[10][117]  ( .D(n12765), .CK(N28803), .Q(n1809), .QN(
        n8208) );
  DFF_X1 \CACHE_MEM_reg[10][116]  ( .D(n12764), .CK(N28803), .Q(n1793), .QN(
        n8224) );
  DFF_X1 \CACHE_MEM_reg[10][115]  ( .D(n12763), .CK(N28803), .Q(n1768), .QN(
        n8240) );
  DFF_X1 \CACHE_MEM_reg[10][114]  ( .D(n12762), .CK(N28803), .Q(n1752), .QN(
        n8256) );
  DFF_X1 \CACHE_MEM_reg[10][113]  ( .D(n12761), .CK(N28803), .Q(n1732), .QN(
        n8272) );
  DFF_X1 \CACHE_MEM_reg[10][112]  ( .D(n12760), .CK(N28803), .Q(n1716), .QN(
        n8288) );
  DFF_X1 \CACHE_MEM_reg[10][111]  ( .D(n12759), .CK(N28803), .Q(n1696), .QN(
        n8304) );
  DFF_X1 \CACHE_MEM_reg[10][110]  ( .D(n12758), .CK(N28803), .Q(n1680), .QN(
        n8320) );
  DFF_X1 \CACHE_MEM_reg[10][109]  ( .D(n12757), .CK(N28803), .Q(n1660), .QN(
        n8336) );
  DFF_X1 \CACHE_MEM_reg[10][108]  ( .D(n12756), .CK(N28803), .Q(n1644), .QN(
        n8352) );
  DFF_X1 \CACHE_MEM_reg[10][107]  ( .D(n12755), .CK(N28803), .Q(n1619), .QN(
        n8368) );
  DFF_X1 \CACHE_MEM_reg[10][106]  ( .D(n12754), .CK(N28803), .Q(n1603), .QN(
        n8384) );
  DFF_X1 \CACHE_MEM_reg[10][105]  ( .D(n12753), .CK(N28803), .Q(n1583), .QN(
        n8400) );
  DFF_X1 \CACHE_MEM_reg[10][104]  ( .D(n12752), .CK(N28803), .Q(n1567), .QN(
        n8416) );
  DFF_X1 \CACHE_MEM_reg[10][103]  ( .D(n12751), .CK(N28803), .Q(n1547), .QN(
        n8432) );
  DFF_X1 \CACHE_MEM_reg[10][102]  ( .D(n12750), .CK(N28803), .Q(n1531), .QN(
        n8448) );
  DFF_X1 \CACHE_MEM_reg[10][101]  ( .D(n12749), .CK(N28803), .Q(n1511), .QN(
        n8464) );
  DFF_X1 \CACHE_MEM_reg[10][100]  ( .D(n12748), .CK(N28803), .Q(n1495), .QN(
        n8480) );
  DFF_X1 \CACHE_MEM_reg[10][99]  ( .D(n12747), .CK(N28803), .Q(n1470), .QN(
        n8496) );
  DFF_X1 \CACHE_MEM_reg[10][98]  ( .D(n12746), .CK(N28803), .Q(n1454), .QN(
        n8512) );
  DFF_X1 \CACHE_MEM_reg[10][97]  ( .D(n12745), .CK(N28803), .Q(n1434), .QN(
        n8528) );
  DFF_X1 \CACHE_MEM_reg[10][96]  ( .D(n12744), .CK(N28803), .Q(n1418), .QN(
        n8544) );
  DFF_X1 \CACHE_MEM_reg[10][95]  ( .D(n12743), .CK(N28803), .Q(n1994), .QN(
        n8560) );
  DFF_X1 \CACHE_MEM_reg[10][94]  ( .D(n12742), .CK(N28803), .Q(n1981), .QN(
        n8576) );
  DFF_X1 \CACHE_MEM_reg[10][93]  ( .D(n12741), .CK(N28803), .Q(n1961), .QN(
        n8592) );
  DFF_X1 \CACHE_MEM_reg[10][92]  ( .D(n12740), .CK(N28803), .Q(n1945), .QN(
        n8608) );
  DFF_X1 \CACHE_MEM_reg[10][91]  ( .D(n12739), .CK(N28803), .Q(n1920), .QN(
        n8624) );
  DFF_X1 \CACHE_MEM_reg[10][90]  ( .D(n12738), .CK(N28803), .Q(n1904), .QN(
        n8640) );
  DFF_X1 \CACHE_MEM_reg[10][89]  ( .D(n12737), .CK(N28803), .Q(n1884), .QN(
        n8656) );
  DFF_X1 \CACHE_MEM_reg[10][88]  ( .D(n12736), .CK(N28803), .Q(n1868), .QN(
        n8672) );
  DFF_X1 \CACHE_MEM_reg[10][87]  ( .D(n12735), .CK(N28803), .Q(n1848), .QN(
        n8688) );
  DFF_X1 \CACHE_MEM_reg[10][86]  ( .D(n12734), .CK(N28803), .Q(n1832), .QN(
        n8704) );
  DFF_X1 \CACHE_MEM_reg[10][85]  ( .D(n12733), .CK(N28803), .Q(n1812), .QN(
        n8720) );
  DFF_X1 \CACHE_MEM_reg[10][84]  ( .D(n12732), .CK(N28803), .Q(n1796), .QN(
        n8736) );
  DFF_X1 \CACHE_MEM_reg[10][83]  ( .D(n12731), .CK(N28803), .Q(n1771), .QN(
        n8752) );
  DFF_X1 \CACHE_MEM_reg[10][82]  ( .D(n12730), .CK(N28803), .Q(n1755), .QN(
        n8768) );
  DFF_X1 \CACHE_MEM_reg[10][81]  ( .D(n12729), .CK(N28803), .Q(n1735), .QN(
        n8784) );
  DFF_X1 \CACHE_MEM_reg[10][80]  ( .D(n12728), .CK(N28803), .Q(n1719), .QN(
        n8800) );
  DFF_X1 \CACHE_MEM_reg[10][79]  ( .D(n12727), .CK(N28803), .Q(n1699), .QN(
        n8816) );
  DFF_X1 \CACHE_MEM_reg[10][78]  ( .D(n12726), .CK(N28803), .Q(n1683), .QN(
        n8832) );
  DFF_X1 \CACHE_MEM_reg[10][77]  ( .D(n12725), .CK(N28803), .Q(n1663), .QN(
        n8848) );
  DFF_X1 \CACHE_MEM_reg[10][76]  ( .D(n12724), .CK(N28803), .Q(n1647), .QN(
        n8864) );
  DFF_X1 \CACHE_MEM_reg[10][75]  ( .D(n12723), .CK(N28803), .Q(n1622), .QN(
        n8880) );
  DFF_X1 \CACHE_MEM_reg[10][74]  ( .D(n12722), .CK(N28803), .Q(n1606), .QN(
        n8896) );
  DFF_X1 \CACHE_MEM_reg[10][73]  ( .D(n12721), .CK(N28803), .Q(n1586), .QN(
        n8912) );
  DFF_X1 \CACHE_MEM_reg[10][72]  ( .D(n12720), .CK(N28803), .Q(n1570), .QN(
        n8928) );
  DFF_X1 \CACHE_MEM_reg[10][71]  ( .D(n12719), .CK(N28803), .Q(n1550), .QN(
        n8944) );
  DFF_X1 \CACHE_MEM_reg[10][70]  ( .D(n12718), .CK(N28803), .Q(n1534), .QN(
        n8960) );
  DFF_X1 \CACHE_MEM_reg[10][69]  ( .D(n12717), .CK(N28803), .Q(n1514), .QN(
        n8976) );
  DFF_X1 \CACHE_MEM_reg[10][68]  ( .D(n12716), .CK(N28803), .Q(n1498), .QN(
        n8992) );
  DFF_X1 \CACHE_MEM_reg[10][67]  ( .D(n12715), .CK(N28803), .Q(n1473), .QN(
        n9008) );
  DFF_X1 \CACHE_MEM_reg[10][66]  ( .D(n12714), .CK(N28803), .Q(n1457), .QN(
        n9024) );
  DFF_X1 \CACHE_MEM_reg[10][65]  ( .D(n12713), .CK(N28803), .Q(n1437), .QN(
        n9040) );
  DFF_X1 \CACHE_MEM_reg[10][64]  ( .D(n12712), .CK(N28803), .Q(n1421), .QN(
        n9056) );
  DFF_X1 \CACHE_MEM_reg[10][63]  ( .D(n12711), .CK(N28803), .Q(n2436), .QN(
        n9072) );
  DFF_X1 \CACHE_MEM_reg[10][62]  ( .D(n12710), .CK(N28803), .Q(n2425), .QN(
        n9088) );
  DFF_X1 \CACHE_MEM_reg[10][61]  ( .D(n12709), .CK(N28803), .Q(n2408), .QN(
        n9104) );
  DFF_X1 \CACHE_MEM_reg[10][60]  ( .D(n12708), .CK(N28803), .Q(n2397), .QN(
        n9120) );
  DFF_X1 \CACHE_MEM_reg[10][59]  ( .D(n12707), .CK(N28803), .Q(n2375), .QN(
        n9136) );
  DFF_X1 \CACHE_MEM_reg[10][58]  ( .D(n12706), .CK(N28803), .Q(n2364), .QN(
        n9152) );
  DFF_X1 \CACHE_MEM_reg[10][57]  ( .D(n12705), .CK(N28803), .Q(n2351), .QN(
        n9168) );
  DFF_X1 \CACHE_MEM_reg[10][56]  ( .D(n12704), .CK(N28803), .Q(n2336), .QN(
        n9184) );
  DFF_X1 \CACHE_MEM_reg[10][55]  ( .D(n12703), .CK(N28803), .Q(n2323), .QN(
        n9200) );
  DFF_X1 \CACHE_MEM_reg[10][54]  ( .D(n12702), .CK(N28803), .Q(n2312), .QN(
        n9216) );
  DFF_X1 \CACHE_MEM_reg[10][53]  ( .D(n12701), .CK(N28803), .Q(n2295), .QN(
        n9232) );
  DFF_X1 \CACHE_MEM_reg[10][52]  ( .D(n12700), .CK(N28803), .Q(n2284), .QN(
        n9248) );
  DFF_X1 \CACHE_MEM_reg[10][51]  ( .D(n12699), .CK(N28803), .Q(n2267), .QN(
        n9264) );
  DFF_X1 \CACHE_MEM_reg[10][50]  ( .D(n12698), .CK(N28803), .Q(n2256), .QN(
        n9280) );
  DFF_X1 \CACHE_MEM_reg[10][49]  ( .D(n12697), .CK(N28803), .Q(n2243), .QN(
        n9296) );
  DFF_X1 \CACHE_MEM_reg[10][48]  ( .D(n12696), .CK(N28803), .Q(n2223), .QN(
        n9312) );
  DFF_X1 \CACHE_MEM_reg[10][47]  ( .D(n12695), .CK(N28803), .Q(n2210), .QN(
        n9328) );
  DFF_X1 \CACHE_MEM_reg[10][46]  ( .D(n12694), .CK(N28803), .Q(n2199), .QN(
        n9344) );
  DFF_X1 \CACHE_MEM_reg[10][45]  ( .D(n12693), .CK(N28803), .Q(n2182), .QN(
        n9360) );
  DFF_X1 \CACHE_MEM_reg[10][44]  ( .D(n12692), .CK(N28803), .Q(n2171), .QN(
        n9376) );
  DFF_X1 \CACHE_MEM_reg[10][43]  ( .D(n12691), .CK(N28803), .Q(n2154), .QN(
        n9392) );
  DFF_X1 \CACHE_MEM_reg[10][42]  ( .D(n12690), .CK(N28803), .Q(n2143), .QN(
        n9408) );
  DFF_X1 \CACHE_MEM_reg[10][41]  ( .D(n12689), .CK(N28803), .Q(n2130), .QN(
        n9424) );
  DFF_X1 \CACHE_MEM_reg[10][40]  ( .D(n12688), .CK(N28803), .Q(n2115), .QN(
        n9440) );
  DFF_X1 \CACHE_MEM_reg[10][39]  ( .D(n12687), .CK(N28803), .Q(n2102), .QN(
        n9456) );
  DFF_X1 \CACHE_MEM_reg[10][38]  ( .D(n12686), .CK(N28803), .Q(n2091), .QN(
        n9472) );
  DFF_X1 \CACHE_MEM_reg[10][37]  ( .D(n12685), .CK(N28803), .Q(n2069), .QN(
        n9488) );
  DFF_X1 \CACHE_MEM_reg[10][36]  ( .D(n12684), .CK(N28803), .Q(n2058), .QN(
        n9504) );
  DFF_X1 \CACHE_MEM_reg[10][35]  ( .D(n12683), .CK(N28803), .Q(n2041), .QN(
        n9520) );
  DFF_X1 \CACHE_MEM_reg[10][34]  ( .D(n12682), .CK(N28803), .Q(n2030), .QN(
        n9536) );
  DFF_X1 \CACHE_MEM_reg[10][33]  ( .D(n12681), .CK(N28803), .Q(n2017), .QN(
        n9552) );
  DFF_X1 \CACHE_MEM_reg[10][32]  ( .D(n12680), .CK(N28803), .Q(n2002), .QN(
        n9568) );
  DFF_X1 \CACHE_MEM_reg[10][31]  ( .D(n12679), .CK(N28803), .Q(n2441), .QN(
        n9584) );
  DFF_X1 \CACHE_MEM_reg[10][30]  ( .D(n12678), .CK(N28803), .Q(n2428), .QN(
        n9600) );
  DFF_X1 \CACHE_MEM_reg[10][29]  ( .D(n12677), .CK(N28803), .Q(n2413), .QN(
        n9616) );
  DFF_X1 \CACHE_MEM_reg[10][28]  ( .D(n12676), .CK(N28803), .Q(n2400), .QN(
        n9632) );
  DFF_X1 \CACHE_MEM_reg[10][27]  ( .D(n12675), .CK(N28803), .Q(n2389), .QN(
        n9648) );
  DFF_X1 \CACHE_MEM_reg[10][26]  ( .D(n12674), .CK(N28803), .Q(n2367), .QN(
        n9664) );
  DFF_X1 \CACHE_MEM_reg[10][25]  ( .D(n12673), .CK(N28803), .Q(n2356), .QN(
        n9680) );
  DFF_X1 \CACHE_MEM_reg[10][24]  ( .D(n12672), .CK(N28803), .Q(n2339), .QN(
        n9696) );
  DFF_X1 \CACHE_MEM_reg[10][23]  ( .D(n12671), .CK(N28803), .Q(n2328), .QN(
        n9712) );
  DFF_X1 \CACHE_MEM_reg[10][22]  ( .D(n12670), .CK(N28803), .Q(n2315), .QN(
        n9728) );
  DFF_X1 \CACHE_MEM_reg[10][21]  ( .D(n12669), .CK(N28803), .Q(n2300), .QN(
        n9744) );
  DFF_X1 \CACHE_MEM_reg[10][20]  ( .D(n12668), .CK(N28803), .Q(n2287), .QN(
        n9760) );
  DFF_X1 \CACHE_MEM_reg[10][19]  ( .D(n12667), .CK(N28803), .Q(n2276), .QN(
        n9776) );
  DFF_X1 \CACHE_MEM_reg[10][18]  ( .D(n12666), .CK(N28803), .Q(n2259), .QN(
        n9792) );
  DFF_X1 \CACHE_MEM_reg[10][17]  ( .D(n12665), .CK(N28803), .Q(n2248), .QN(
        n9808) );
  DFF_X1 \CACHE_MEM_reg[10][16]  ( .D(n12664), .CK(N28803), .Q(n2226), .QN(
        n9824) );
  DFF_X1 \CACHE_MEM_reg[10][15]  ( .D(n12663), .CK(N28803), .Q(n2215), .QN(
        n9840) );
  DFF_X1 \CACHE_MEM_reg[10][14]  ( .D(n12662), .CK(N28803), .Q(n2202), .QN(
        n9856) );
  DFF_X1 \CACHE_MEM_reg[10][13]  ( .D(n12661), .CK(N28803), .Q(n2187), .QN(
        n9872) );
  DFF_X1 \CACHE_MEM_reg[10][12]  ( .D(n12660), .CK(N28803), .Q(n2174), .QN(
        n9888) );
  DFF_X1 \CACHE_MEM_reg[10][11]  ( .D(n12659), .CK(N28803), .Q(n2163), .QN(
        n9904) );
  DFF_X1 \CACHE_MEM_reg[10][10]  ( .D(n12658), .CK(N28803), .Q(n2146), .QN(
        n9920) );
  DFF_X1 \CACHE_MEM_reg[10][9]  ( .D(n12657), .CK(N28803), .Q(n2135), .QN(
        n9936) );
  DFF_X1 \CACHE_MEM_reg[10][8]  ( .D(n12656), .CK(N28803), .Q(n2118), .QN(
        n9952) );
  DFF_X1 \CACHE_MEM_reg[10][7]  ( .D(n12655), .CK(N28803), .Q(n2107), .QN(
        n9968) );
  DFF_X1 \CACHE_MEM_reg[10][6]  ( .D(n12654), .CK(N28803), .Q(n2094), .QN(
        n9984) );
  DFF_X1 \CACHE_MEM_reg[10][5]  ( .D(n12653), .CK(N28803), .Q(n2074), .QN(
        n10000) );
  DFF_X1 \CACHE_MEM_reg[10][4]  ( .D(n12652), .CK(N28803), .Q(n2061), .QN(
        n10016) );
  DFF_X1 \CACHE_MEM_reg[10][3]  ( .D(n12651), .CK(N28803), .Q(n2050), .QN(
        n10032) );
  DFF_X1 \CACHE_MEM_reg[10][2]  ( .D(n12650), .CK(N28803), .Q(n2033), .QN(
        n10048) );
  DFF_X1 \CACHE_MEM_reg[10][1]  ( .D(n12649), .CK(N28803), .Q(n2022), .QN(
        n10064) );
  DFF_X1 \CACHE_MEM_reg[10][0]  ( .D(n12648), .CK(N28803), .Q(n2005), .QN(
        n10080) );
  DFF_X1 \CACHE_MEM_reg[9][255]  ( .D(n12647), .CK(N28803), .Q(n3789), .QN(
        n5996) );
  DFF_X1 \CACHE_MEM_reg[9][254]  ( .D(n12646), .CK(N28803), .Q(n3781), .QN(
        n6012) );
  DFF_X1 \CACHE_MEM_reg[9][253]  ( .D(n12645), .CK(N28803), .Q(n3774), .QN(
        n6028) );
  DFF_X1 \CACHE_MEM_reg[9][252]  ( .D(n12644), .CK(N28803), .Q(n3768), .QN(
        n6044) );
  DFF_X1 \CACHE_MEM_reg[9][251]  ( .D(n12643), .CK(N28803), .Q(n3757), .QN(
        n6060) );
  DFF_X1 \CACHE_MEM_reg[9][250]  ( .D(n12642), .CK(N28803), .Q(n3753), .QN(
        n6076) );
  DFF_X1 \CACHE_MEM_reg[9][249]  ( .D(n12641), .CK(N28803), .Q(n3746), .QN(
        n6092) );
  DFF_X1 \CACHE_MEM_reg[9][248]  ( .D(n12640), .CK(N28803), .Q(n3740), .QN(
        n6108) );
  DFF_X1 \CACHE_MEM_reg[9][247]  ( .D(n12639), .CK(N28803), .Q(n3733), .QN(
        n6124) );
  DFF_X1 \CACHE_MEM_reg[9][246]  ( .D(n12638), .CK(N28803), .Q(n3729), .QN(
        n6140) );
  DFF_X1 \CACHE_MEM_reg[9][245]  ( .D(n12637), .CK(N28803), .Q(n3713), .QN(
        n6156) );
  DFF_X1 \CACHE_MEM_reg[9][244]  ( .D(n12636), .CK(N28803), .Q(n3707), .QN(
        n6172) );
  DFF_X1 \CACHE_MEM_reg[9][243]  ( .D(n12635), .CK(N28803), .Q(n3700), .QN(
        n6188) );
  DFF_X1 \CACHE_MEM_reg[9][242]  ( .D(n12634), .CK(N28803), .Q(n3696), .QN(
        n6204) );
  DFF_X1 \CACHE_MEM_reg[9][241]  ( .D(n12633), .CK(N28803), .Q(n3689), .QN(
        n6220) );
  DFF_X1 \CACHE_MEM_reg[9][240]  ( .D(n12632), .CK(N28803), .Q(n3679), .QN(
        n6236) );
  DFF_X1 \CACHE_MEM_reg[9][239]  ( .D(n12631), .CK(N28803), .Q(n3672), .QN(
        n6252) );
  DFF_X1 \CACHE_MEM_reg[9][238]  ( .D(n12630), .CK(N28803), .Q(n3668), .QN(
        n6268) );
  DFF_X1 \CACHE_MEM_reg[9][237]  ( .D(n12629), .CK(N28803), .Q(n3661), .QN(
        n6284) );
  DFF_X1 \CACHE_MEM_reg[9][236]  ( .D(n12628), .CK(N28803), .Q(n3655), .QN(
        n6300) );
  DFF_X1 \CACHE_MEM_reg[9][235]  ( .D(n12627), .CK(N28803), .Q(n3644), .QN(
        n6316) );
  DFF_X1 \CACHE_MEM_reg[9][234]  ( .D(n12626), .CK(N28803), .Q(n3640), .QN(
        n6332) );
  DFF_X1 \CACHE_MEM_reg[9][233]  ( .D(n12625), .CK(N28803), .Q(n3633), .QN(
        n6348) );
  DFF_X1 \CACHE_MEM_reg[9][232]  ( .D(n12624), .CK(N28803), .Q(n3627), .QN(
        n6364) );
  DFF_X1 \CACHE_MEM_reg[9][231]  ( .D(n12623), .CK(N28803), .Q(n3620), .QN(
        n6380) );
  DFF_X1 \CACHE_MEM_reg[9][230]  ( .D(n12622), .CK(N28803), .Q(n3616), .QN(
        n6396) );
  DFF_X1 \CACHE_MEM_reg[9][229]  ( .D(n12621), .CK(N28803), .Q(n3605), .QN(
        n6412) );
  DFF_X1 \CACHE_MEM_reg[9][228]  ( .D(n12620), .CK(N28803), .Q(n3599), .QN(
        n6428) );
  DFF_X1 \CACHE_MEM_reg[9][227]  ( .D(n12619), .CK(N28803), .Q(n3592), .QN(
        n6444) );
  DFF_X1 \CACHE_MEM_reg[9][226]  ( .D(n12618), .CK(N28803), .Q(n3588), .QN(
        n6460) );
  DFF_X1 \CACHE_MEM_reg[9][225]  ( .D(n12617), .CK(N28803), .Q(n3581), .QN(
        n6476) );
  DFF_X1 \CACHE_MEM_reg[9][224]  ( .D(n12616), .CK(N28803), .Q(n3566), .QN(
        n6492) );
  DFF_X1 \CACHE_MEM_reg[9][223]  ( .D(n12615), .CK(N28803), .Q(n5259), .QN(
        n6508) );
  DFF_X1 \CACHE_MEM_reg[9][222]  ( .D(n12614), .CK(N28803), .Q(n5244), .QN(
        n6524) );
  DFF_X1 \CACHE_MEM_reg[9][221]  ( .D(n12613), .CK(N28803), .Q(n5231), .QN(
        n6540) );
  DFF_X1 \CACHE_MEM_reg[9][220]  ( .D(n12612), .CK(N28803), .Q(n5220), .QN(
        n6556) );
  DFF_X1 \CACHE_MEM_reg[9][219]  ( .D(n12611), .CK(N28803), .Q(n5198), .QN(
        n6572) );
  DFF_X1 \CACHE_MEM_reg[9][218]  ( .D(n12610), .CK(N28803), .Q(n5187), .QN(
        n6588) );
  DFF_X1 \CACHE_MEM_reg[9][217]  ( .D(n12609), .CK(N28803), .Q(n5170), .QN(
        n6604) );
  DFF_X1 \CACHE_MEM_reg[9][216]  ( .D(n12608), .CK(N28803), .Q(n5159), .QN(
        n6620) );
  DFF_X1 \CACHE_MEM_reg[9][215]  ( .D(n12607), .CK(N28803), .Q(n5146), .QN(
        n6636) );
  DFF_X1 \CACHE_MEM_reg[9][214]  ( .D(n12606), .CK(N28803), .Q(n5131), .QN(
        n6652) );
  DFF_X1 \CACHE_MEM_reg[9][213]  ( .D(n12605), .CK(N28803), .Q(n5118), .QN(
        n6668) );
  DFF_X1 \CACHE_MEM_reg[9][212]  ( .D(n12604), .CK(N28803), .Q(n5107), .QN(
        n6684) );
  DFF_X1 \CACHE_MEM_reg[9][211]  ( .D(n12603), .CK(N28803), .Q(n5090), .QN(
        n6700) );
  DFF_X1 \CACHE_MEM_reg[9][210]  ( .D(n12602), .CK(N28803), .Q(n5079), .QN(
        n6716) );
  DFF_X1 \CACHE_MEM_reg[9][209]  ( .D(n12601), .CK(N28803), .Q(n5057), .QN(
        n6732) );
  DFF_X1 \CACHE_MEM_reg[9][208]  ( .D(n12600), .CK(N28803), .Q(n5049), .QN(
        n6748) );
  DFF_X1 \CACHE_MEM_reg[9][207]  ( .D(n12599), .CK(N28803), .Q(n5038), .QN(
        n6764) );
  DFF_X1 \CACHE_MEM_reg[9][206]  ( .D(n12598), .CK(N28803), .Q(n5021), .QN(
        n6780) );
  DFF_X1 \CACHE_MEM_reg[9][205]  ( .D(n12597), .CK(N28803), .Q(n5010), .QN(
        n6796) );
  DFF_X1 \CACHE_MEM_reg[9][204]  ( .D(n12596), .CK(N28803), .Q(n4997), .QN(
        n6812) );
  DFF_X1 \CACHE_MEM_reg[9][203]  ( .D(n12595), .CK(N28803), .Q(n4982), .QN(
        n6828) );
  DFF_X1 \CACHE_MEM_reg[9][202]  ( .D(n12594), .CK(N28803), .Q(n4969), .QN(
        n6844) );
  DFF_X1 \CACHE_MEM_reg[9][201]  ( .D(n12593), .CK(N28803), .Q(n4958), .QN(
        n6860) );
  DFF_X1 \CACHE_MEM_reg[9][200]  ( .D(n12592), .CK(N28803), .Q(n4941), .QN(
        n6876) );
  DFF_X1 \CACHE_MEM_reg[9][199]  ( .D(n12591), .CK(N28803), .Q(n4930), .QN(
        n6892) );
  DFF_X1 \CACHE_MEM_reg[9][198]  ( .D(n12590), .CK(N28803), .Q(n4908), .QN(
        n6908) );
  DFF_X1 \CACHE_MEM_reg[9][197]  ( .D(n12589), .CK(N28803), .Q(n4897), .QN(
        n6924) );
  DFF_X1 \CACHE_MEM_reg[9][196]  ( .D(n12588), .CK(N28803), .Q(n4884), .QN(
        n6940) );
  DFF_X1 \CACHE_MEM_reg[9][195]  ( .D(n12587), .CK(N28803), .Q(n4869), .QN(
        n6956) );
  DFF_X1 \CACHE_MEM_reg[9][194]  ( .D(n12586), .CK(N28803), .Q(n4856), .QN(
        n6972) );
  DFF_X1 \CACHE_MEM_reg[9][193]  ( .D(n12585), .CK(N28803), .Q(n4845), .QN(
        n6988) );
  DFF_X1 \CACHE_MEM_reg[9][192]  ( .D(n12584), .CK(N28803), .Q(n4828), .QN(
        n7004) );
  DFF_X1 \CACHE_MEM_reg[9][191]  ( .D(n12583), .CK(N28803), .Q(n5703), .QN(
        n7020) );
  DFF_X1 \CACHE_MEM_reg[9][190]  ( .D(n12582), .CK(N28803), .Q(n3782), .QN(
        n7036) );
  DFF_X1 \CACHE_MEM_reg[9][189]  ( .D(n12581), .CK(N28803), .Q(n3776), .QN(
        n7052) );
  DFF_X1 \CACHE_MEM_reg[9][188]  ( .D(n12580), .CK(N28803), .Q(n3769), .QN(
        n7068) );
  DFF_X1 \CACHE_MEM_reg[9][187]  ( .D(n12579), .CK(N28803), .Q(n3765), .QN(
        n7084) );
  DFF_X1 \CACHE_MEM_reg[9][186]  ( .D(n12578), .CK(N28803), .Q(n3754), .QN(
        n7100) );
  DFF_X1 \CACHE_MEM_reg[9][185]  ( .D(n12577), .CK(N28803), .Q(n3748), .QN(
        n7116) );
  DFF_X1 \CACHE_MEM_reg[9][184]  ( .D(n12576), .CK(N28803), .Q(n3741), .QN(
        n7132) );
  DFF_X1 \CACHE_MEM_reg[9][183]  ( .D(n12575), .CK(N28803), .Q(n3737), .QN(
        n7148) );
  DFF_X1 \CACHE_MEM_reg[9][182]  ( .D(n12574), .CK(N28803), .Q(n3730), .QN(
        n7164) );
  DFF_X1 \CACHE_MEM_reg[9][181]  ( .D(n12573), .CK(N28803), .Q(n3715), .QN(
        n7180) );
  DFF_X1 \CACHE_MEM_reg[9][180]  ( .D(n12572), .CK(N28803), .Q(n3708), .QN(
        n7196) );
  DFF_X1 \CACHE_MEM_reg[9][179]  ( .D(n12571), .CK(N28803), .Q(n3704), .QN(
        n7212) );
  DFF_X1 \CACHE_MEM_reg[9][178]  ( .D(n12570), .CK(N28803), .Q(n3697), .QN(
        n7228) );
  DFF_X1 \CACHE_MEM_reg[9][177]  ( .D(n12569), .CK(N28803), .Q(n3691), .QN(
        n7244) );
  DFF_X1 \CACHE_MEM_reg[9][176]  ( .D(n12568), .CK(N28803), .Q(n3680), .QN(
        n7260) );
  DFF_X1 \CACHE_MEM_reg[9][175]  ( .D(n12567), .CK(N28803), .Q(n3676), .QN(
        n7276) );
  DFF_X1 \CACHE_MEM_reg[9][174]  ( .D(n12566), .CK(N28803), .Q(n3669), .QN(
        n7292) );
  DFF_X1 \CACHE_MEM_reg[9][173]  ( .D(n12565), .CK(N28803), .Q(n3663), .QN(
        n7308) );
  DFF_X1 \CACHE_MEM_reg[9][172]  ( .D(n12564), .CK(N28803), .Q(n3656), .QN(
        n7324) );
  DFF_X1 \CACHE_MEM_reg[9][171]  ( .D(n12563), .CK(N28803), .Q(n3652), .QN(
        n7340) );
  DFF_X1 \CACHE_MEM_reg[9][170]  ( .D(n12562), .CK(N28803), .Q(n3641), .QN(
        n7356) );
  DFF_X1 \CACHE_MEM_reg[9][169]  ( .D(n12561), .CK(N28803), .Q(n3635), .QN(
        n7372) );
  DFF_X1 \CACHE_MEM_reg[9][168]  ( .D(n12560), .CK(N28803), .Q(n3628), .QN(
        n7388) );
  DFF_X1 \CACHE_MEM_reg[9][167]  ( .D(n12559), .CK(N28803), .Q(n3624), .QN(
        n7404) );
  DFF_X1 \CACHE_MEM_reg[9][166]  ( .D(n12558), .CK(N28803), .Q(n3617), .QN(
        n7420) );
  DFF_X1 \CACHE_MEM_reg[9][165]  ( .D(n12557), .CK(N28803), .Q(n3607), .QN(
        n7436) );
  DFF_X1 \CACHE_MEM_reg[9][164]  ( .D(n12556), .CK(N28803), .Q(n3600), .QN(
        n7452) );
  DFF_X1 \CACHE_MEM_reg[9][163]  ( .D(n12555), .CK(N28803), .Q(n3596), .QN(
        n7468) );
  DFF_X1 \CACHE_MEM_reg[9][162]  ( .D(n12554), .CK(N28803), .Q(n3589), .QN(
        n7484) );
  DFF_X1 \CACHE_MEM_reg[9][161]  ( .D(n12553), .CK(N28803), .Q(n3583), .QN(
        n7500) );
  DFF_X1 \CACHE_MEM_reg[9][160]  ( .D(n12552), .CK(N28803), .Q(n3567), .QN(
        n7516) );
  DFF_X1 \CACHE_MEM_reg[9][159]  ( .D(n12551), .CK(N28803), .Q(n5706), .QN(
        n7532) );
  DFF_X1 \CACHE_MEM_reg[9][158]  ( .D(n12550), .CK(N28803), .Q(n5691), .QN(
        n7548) );
  DFF_X1 \CACHE_MEM_reg[9][157]  ( .D(n12549), .CK(N28803), .Q(n5678), .QN(
        n7564) );
  DFF_X1 \CACHE_MEM_reg[9][156]  ( .D(n12548), .CK(N28803), .Q(n5667), .QN(
        n7580) );
  DFF_X1 \CACHE_MEM_reg[9][155]  ( .D(n12547), .CK(N28803), .Q(n5645), .QN(
        n7596) );
  DFF_X1 \CACHE_MEM_reg[9][154]  ( .D(n12546), .CK(N28803), .Q(n5634), .QN(
        n7612) );
  DFF_X1 \CACHE_MEM_reg[9][153]  ( .D(n12545), .CK(N28803), .Q(n5617), .QN(
        n7628) );
  DFF_X1 \CACHE_MEM_reg[9][152]  ( .D(n12544), .CK(N28803), .Q(n5606), .QN(
        n7644) );
  DFF_X1 \CACHE_MEM_reg[9][151]  ( .D(n12543), .CK(N28803), .Q(n5593), .QN(
        n7660) );
  DFF_X1 \CACHE_MEM_reg[9][150]  ( .D(n12542), .CK(N28803), .Q(n5578), .QN(
        n7676) );
  DFF_X1 \CACHE_MEM_reg[9][149]  ( .D(n12541), .CK(N28803), .Q(n5565), .QN(
        n7692) );
  DFF_X1 \CACHE_MEM_reg[9][148]  ( .D(n12540), .CK(N28803), .Q(n5554), .QN(
        n7708) );
  DFF_X1 \CACHE_MEM_reg[9][147]  ( .D(n12539), .CK(N28803), .Q(n5537), .QN(
        n7724) );
  DFF_X1 \CACHE_MEM_reg[9][146]  ( .D(n12538), .CK(N28803), .Q(n5526), .QN(
        n7740) );
  DFF_X1 \CACHE_MEM_reg[9][145]  ( .D(n12537), .CK(N28803), .Q(n5504), .QN(
        n7756) );
  DFF_X1 \CACHE_MEM_reg[9][144]  ( .D(n12536), .CK(N28803), .Q(n5493), .QN(
        n7772) );
  DFF_X1 \CACHE_MEM_reg[9][143]  ( .D(n12535), .CK(N28803), .Q(n5480), .QN(
        n7788) );
  DFF_X1 \CACHE_MEM_reg[9][142]  ( .D(n12534), .CK(N28803), .Q(n5465), .QN(
        n7804) );
  DFF_X1 \CACHE_MEM_reg[9][141]  ( .D(n12533), .CK(N28803), .Q(n5452), .QN(
        n7820) );
  DFF_X1 \CACHE_MEM_reg[9][140]  ( .D(n12532), .CK(N28803), .Q(n5441), .QN(
        n7836) );
  DFF_X1 \CACHE_MEM_reg[9][139]  ( .D(n12531), .CK(N28803), .Q(n5424), .QN(
        n7852) );
  DFF_X1 \CACHE_MEM_reg[9][138]  ( .D(n12530), .CK(N28803), .Q(n5413), .QN(
        n7868) );
  DFF_X1 \CACHE_MEM_reg[9][137]  ( .D(n12529), .CK(N28803), .Q(n5396), .QN(
        n7884) );
  DFF_X1 \CACHE_MEM_reg[9][136]  ( .D(n12528), .CK(N28803), .Q(n5385), .QN(
        n7900) );
  DFF_X1 \CACHE_MEM_reg[9][135]  ( .D(n12527), .CK(N28803), .Q(n5372), .QN(
        n7916) );
  DFF_X1 \CACHE_MEM_reg[9][134]  ( .D(n12526), .CK(N28803), .Q(n5352), .QN(
        n7932) );
  DFF_X1 \CACHE_MEM_reg[9][133]  ( .D(n12525), .CK(N28803), .Q(n5339), .QN(
        n7948) );
  DFF_X1 \CACHE_MEM_reg[9][132]  ( .D(n12524), .CK(N28803), .Q(n5328), .QN(
        n7964) );
  DFF_X1 \CACHE_MEM_reg[9][131]  ( .D(n12523), .CK(N28803), .Q(n5311), .QN(
        n7980) );
  DFF_X1 \CACHE_MEM_reg[9][130]  ( .D(n12522), .CK(N28803), .Q(n5300), .QN(
        n7996) );
  DFF_X1 \CACHE_MEM_reg[9][129]  ( .D(n12521), .CK(N28803), .Q(n5283), .QN(
        n8012) );
  DFF_X1 \CACHE_MEM_reg[9][128]  ( .D(n12520), .CK(N28803), .Q(n5272), .QN(
        n8028) );
  DFF_X1 \CACHE_MEM_reg[9][127]  ( .D(n12519), .CK(N28803), .Q(n3784), .QN(
        n8044) );
  DFF_X1 \CACHE_MEM_reg[9][126]  ( .D(n12518), .CK(N28803), .Q(n4350), .QN(
        n8060) );
  DFF_X1 \CACHE_MEM_reg[9][125]  ( .D(n12517), .CK(N28803), .Q(n4334), .QN(
        n8076) );
  DFF_X1 \CACHE_MEM_reg[9][124]  ( .D(n12516), .CK(N28803), .Q(n4309), .QN(
        n8092) );
  DFF_X1 \CACHE_MEM_reg[9][123]  ( .D(n12515), .CK(N28803), .Q(n4293), .QN(
        n8108) );
  DFF_X1 \CACHE_MEM_reg[9][122]  ( .D(n12514), .CK(N28803), .Q(n4273), .QN(
        n8124) );
  DFF_X1 \CACHE_MEM_reg[9][121]  ( .D(n12513), .CK(N28803), .Q(n4257), .QN(
        n8140) );
  DFF_X1 \CACHE_MEM_reg[9][120]  ( .D(n12512), .CK(N28803), .Q(n4237), .QN(
        n8156) );
  DFF_X1 \CACHE_MEM_reg[9][119]  ( .D(n12511), .CK(N28803), .Q(n4221), .QN(
        n8172) );
  DFF_X1 \CACHE_MEM_reg[9][118]  ( .D(n12510), .CK(N28803), .Q(n4201), .QN(
        n8188) );
  DFF_X1 \CACHE_MEM_reg[9][117]  ( .D(n12509), .CK(N28803), .Q(n4185), .QN(
        n8204) );
  DFF_X1 \CACHE_MEM_reg[9][116]  ( .D(n12508), .CK(N28803), .Q(n4160), .QN(
        n8220) );
  DFF_X1 \CACHE_MEM_reg[9][115]  ( .D(n12507), .CK(N28803), .Q(n4144), .QN(
        n8236) );
  DFF_X1 \CACHE_MEM_reg[9][114]  ( .D(n12506), .CK(N28803), .Q(n4124), .QN(
        n8252) );
  DFF_X1 \CACHE_MEM_reg[9][113]  ( .D(n12505), .CK(N28803), .Q(n4108), .QN(
        n8268) );
  DFF_X1 \CACHE_MEM_reg[9][112]  ( .D(n12504), .CK(N28803), .Q(n4088), .QN(
        n8284) );
  DFF_X1 \CACHE_MEM_reg[9][111]  ( .D(n12503), .CK(N28803), .Q(n4072), .QN(
        n8300) );
  DFF_X1 \CACHE_MEM_reg[9][110]  ( .D(n12502), .CK(N28803), .Q(n4052), .QN(
        n8316) );
  DFF_X1 \CACHE_MEM_reg[9][109]  ( .D(n12501), .CK(N28803), .Q(n4036), .QN(
        n8332) );
  DFF_X1 \CACHE_MEM_reg[9][108]  ( .D(n12500), .CK(N28803), .Q(n4011), .QN(
        n8348) );
  DFF_X1 \CACHE_MEM_reg[9][107]  ( .D(n12499), .CK(N28803), .Q(n3995), .QN(
        n8364) );
  DFF_X1 \CACHE_MEM_reg[9][106]  ( .D(n12498), .CK(N28803), .Q(n3975), .QN(
        n8380) );
  DFF_X1 \CACHE_MEM_reg[9][105]  ( .D(n12497), .CK(N28803), .Q(n3959), .QN(
        n8396) );
  DFF_X1 \CACHE_MEM_reg[9][104]  ( .D(n12496), .CK(N28803), .Q(n3939), .QN(
        n8412) );
  DFF_X1 \CACHE_MEM_reg[9][103]  ( .D(n12495), .CK(N28803), .Q(n3923), .QN(
        n8428) );
  DFF_X1 \CACHE_MEM_reg[9][102]  ( .D(n12494), .CK(N28803), .Q(n3903), .QN(
        n8444) );
  DFF_X1 \CACHE_MEM_reg[9][101]  ( .D(n12493), .CK(N28803), .Q(n3887), .QN(
        n8460) );
  DFF_X1 \CACHE_MEM_reg[9][100]  ( .D(n12492), .CK(N28803), .Q(n3862), .QN(
        n8476) );
  DFF_X1 \CACHE_MEM_reg[9][99]  ( .D(n12491), .CK(N28803), .Q(n3846), .QN(
        n8492) );
  DFF_X1 \CACHE_MEM_reg[9][98]  ( .D(n12490), .CK(N28803), .Q(n3826), .QN(
        n8508) );
  DFF_X1 \CACHE_MEM_reg[9][97]  ( .D(n12489), .CK(N28803), .Q(n3810), .QN(
        n8524) );
  DFF_X1 \CACHE_MEM_reg[9][96]  ( .D(n12488), .CK(N28803), .Q(n3790), .QN(
        n8540) );
  DFF_X1 \CACHE_MEM_reg[9][95]  ( .D(n12487), .CK(N28803), .Q(n4370), .QN(
        n8556) );
  DFF_X1 \CACHE_MEM_reg[9][94]  ( .D(n12486), .CK(N28803), .Q(n4353), .QN(
        n8572) );
  DFF_X1 \CACHE_MEM_reg[9][93]  ( .D(n12485), .CK(N28803), .Q(n4337), .QN(
        n8588) );
  DFF_X1 \CACHE_MEM_reg[9][92]  ( .D(n12484), .CK(N28803), .Q(n4312), .QN(
        n8604) );
  DFF_X1 \CACHE_MEM_reg[9][91]  ( .D(n12483), .CK(N28803), .Q(n4296), .QN(
        n8620) );
  DFF_X1 \CACHE_MEM_reg[9][90]  ( .D(n12482), .CK(N28803), .Q(n4276), .QN(
        n8636) );
  DFF_X1 \CACHE_MEM_reg[9][89]  ( .D(n12481), .CK(N28803), .Q(n4260), .QN(
        n8652) );
  DFF_X1 \CACHE_MEM_reg[9][88]  ( .D(n12480), .CK(N28803), .Q(n4240), .QN(
        n8668) );
  DFF_X1 \CACHE_MEM_reg[9][87]  ( .D(n12479), .CK(N28803), .Q(n4224), .QN(
        n8684) );
  DFF_X1 \CACHE_MEM_reg[9][86]  ( .D(n12478), .CK(N28803), .Q(n4204), .QN(
        n8700) );
  DFF_X1 \CACHE_MEM_reg[9][85]  ( .D(n12477), .CK(N28803), .Q(n4188), .QN(
        n8716) );
  DFF_X1 \CACHE_MEM_reg[9][84]  ( .D(n12476), .CK(N28803), .Q(n4163), .QN(
        n8732) );
  DFF_X1 \CACHE_MEM_reg[9][83]  ( .D(n12475), .CK(N28803), .Q(n4147), .QN(
        n8748) );
  DFF_X1 \CACHE_MEM_reg[9][82]  ( .D(n12474), .CK(N28803), .Q(n4127), .QN(
        n8764) );
  DFF_X1 \CACHE_MEM_reg[9][81]  ( .D(n12473), .CK(N28803), .Q(n4111), .QN(
        n8780) );
  DFF_X1 \CACHE_MEM_reg[9][80]  ( .D(n12472), .CK(N28803), .Q(n4091), .QN(
        n8796) );
  DFF_X1 \CACHE_MEM_reg[9][79]  ( .D(n12471), .CK(N28803), .Q(n4075), .QN(
        n8812) );
  DFF_X1 \CACHE_MEM_reg[9][78]  ( .D(n12470), .CK(N28803), .Q(n4055), .QN(
        n8828) );
  DFF_X1 \CACHE_MEM_reg[9][77]  ( .D(n12469), .CK(N28803), .Q(n4039), .QN(
        n8844) );
  DFF_X1 \CACHE_MEM_reg[9][76]  ( .D(n12468), .CK(N28803), .Q(n4014), .QN(
        n8860) );
  DFF_X1 \CACHE_MEM_reg[9][75]  ( .D(n12467), .CK(N28803), .Q(n3998), .QN(
        n8876) );
  DFF_X1 \CACHE_MEM_reg[9][74]  ( .D(n12466), .CK(N28803), .Q(n3978), .QN(
        n8892) );
  DFF_X1 \CACHE_MEM_reg[9][73]  ( .D(n12465), .CK(N28803), .Q(n3962), .QN(
        n8908) );
  DFF_X1 \CACHE_MEM_reg[9][72]  ( .D(n12464), .CK(N28803), .Q(n3942), .QN(
        n8924) );
  DFF_X1 \CACHE_MEM_reg[9][71]  ( .D(n12463), .CK(N28803), .Q(n3926), .QN(
        n8940) );
  DFF_X1 \CACHE_MEM_reg[9][70]  ( .D(n12462), .CK(N28803), .Q(n3906), .QN(
        n8956) );
  DFF_X1 \CACHE_MEM_reg[9][69]  ( .D(n12461), .CK(N28803), .Q(n3890), .QN(
        n8972) );
  DFF_X1 \CACHE_MEM_reg[9][68]  ( .D(n12460), .CK(N28803), .Q(n3865), .QN(
        n8988) );
  DFF_X1 \CACHE_MEM_reg[9][67]  ( .D(n12459), .CK(N28803), .Q(n3849), .QN(
        n9004) );
  DFF_X1 \CACHE_MEM_reg[9][66]  ( .D(n12458), .CK(N28803), .Q(n3829), .QN(
        n9020) );
  DFF_X1 \CACHE_MEM_reg[9][65]  ( .D(n12457), .CK(N28803), .Q(n3813), .QN(
        n9036) );
  DFF_X1 \CACHE_MEM_reg[9][64]  ( .D(n12456), .CK(N28803), .Q(n3793), .QN(
        n9052) );
  DFF_X1 \CACHE_MEM_reg[9][63]  ( .D(n12455), .CK(N28803), .Q(n3785), .QN(
        n9068) );
  DFF_X1 \CACHE_MEM_reg[9][62]  ( .D(n12454), .CK(N28803), .Q(n3777), .QN(
        n9084) );
  DFF_X1 \CACHE_MEM_reg[9][61]  ( .D(n12453), .CK(N28803), .Q(n3773), .QN(
        n9100) );
  DFF_X1 \CACHE_MEM_reg[9][60]  ( .D(n12452), .CK(N28803), .Q(n3766), .QN(
        n9116) );
  DFF_X1 \CACHE_MEM_reg[9][59]  ( .D(n12451), .CK(N28803), .Q(n3756), .QN(
        n9132) );
  DFF_X1 \CACHE_MEM_reg[9][58]  ( .D(n12450), .CK(N28803), .Q(n3749), .QN(
        n9148) );
  DFF_X1 \CACHE_MEM_reg[9][57]  ( .D(n12449), .CK(N28803), .Q(n3745), .QN(
        n9164) );
  DFF_X1 \CACHE_MEM_reg[9][56]  ( .D(n12448), .CK(N28803), .Q(n3738), .QN(
        n9180) );
  DFF_X1 \CACHE_MEM_reg[9][55]  ( .D(n12447), .CK(N28803), .Q(n3732), .QN(
        n9196) );
  DFF_X1 \CACHE_MEM_reg[9][54]  ( .D(n12446), .CK(N28803), .Q(n3716), .QN(
        n9212) );
  DFF_X1 \CACHE_MEM_reg[9][53]  ( .D(n12445), .CK(N28803), .Q(n3712), .QN(
        n9228) );
  DFF_X1 \CACHE_MEM_reg[9][52]  ( .D(n12444), .CK(N28803), .Q(n3705), .QN(
        n9244) );
  DFF_X1 \CACHE_MEM_reg[9][51]  ( .D(n12443), .CK(N28803), .Q(n3699), .QN(
        n9260) );
  DFF_X1 \CACHE_MEM_reg[9][50]  ( .D(n12442), .CK(N28803), .Q(n3692), .QN(
        n9276) );
  DFF_X1 \CACHE_MEM_reg[9][49]  ( .D(n12441), .CK(N28803), .Q(n3688), .QN(
        n9292) );
  DFF_X1 \CACHE_MEM_reg[9][48]  ( .D(n12440), .CK(N28803), .Q(n3677), .QN(
        n9308) );
  DFF_X1 \CACHE_MEM_reg[9][47]  ( .D(n12439), .CK(N28803), .Q(n3671), .QN(
        n9324) );
  DFF_X1 \CACHE_MEM_reg[9][46]  ( .D(n12438), .CK(N28803), .Q(n3664), .QN(
        n9340) );
  DFF_X1 \CACHE_MEM_reg[9][45]  ( .D(n12437), .CK(N28803), .Q(n3660), .QN(
        n9356) );
  DFF_X1 \CACHE_MEM_reg[9][44]  ( .D(n12436), .CK(N28803), .Q(n3653), .QN(
        n9372) );
  DFF_X1 \CACHE_MEM_reg[9][43]  ( .D(n12435), .CK(N28803), .Q(n3643), .QN(
        n9388) );
  DFF_X1 \CACHE_MEM_reg[9][42]  ( .D(n12434), .CK(N28803), .Q(n3636), .QN(
        n9404) );
  DFF_X1 \CACHE_MEM_reg[9][41]  ( .D(n12433), .CK(N28803), .Q(n3632), .QN(
        n9420) );
  DFF_X1 \CACHE_MEM_reg[9][40]  ( .D(n12432), .CK(N28803), .Q(n3625), .QN(
        n9436) );
  DFF_X1 \CACHE_MEM_reg[9][39]  ( .D(n12431), .CK(N28803), .Q(n3619), .QN(
        n9452) );
  DFF_X1 \CACHE_MEM_reg[9][38]  ( .D(n12430), .CK(N28803), .Q(n3608), .QN(
        n9468) );
  DFF_X1 \CACHE_MEM_reg[9][37]  ( .D(n12429), .CK(N28803), .Q(n3604), .QN(
        n9484) );
  DFF_X1 \CACHE_MEM_reg[9][36]  ( .D(n12428), .CK(N28803), .Q(n3597), .QN(
        n9500) );
  DFF_X1 \CACHE_MEM_reg[9][35]  ( .D(n12427), .CK(N28803), .Q(n3591), .QN(
        n9516) );
  DFF_X1 \CACHE_MEM_reg[9][34]  ( .D(n12426), .CK(N28803), .Q(n3584), .QN(
        n9532) );
  DFF_X1 \CACHE_MEM_reg[9][33]  ( .D(n12425), .CK(N28803), .Q(n3580), .QN(
        n9548) );
  DFF_X1 \CACHE_MEM_reg[9][32]  ( .D(n12424), .CK(N28803), .Q(n3564), .QN(
        n9564) );
  DFF_X1 \CACHE_MEM_reg[9][31]  ( .D(n12423), .CK(N28803), .Q(n4817), .QN(
        n9580) );
  DFF_X1 \CACHE_MEM_reg[9][30]  ( .D(n12422), .CK(N28803), .Q(n4800), .QN(
        n9596) );
  DFF_X1 \CACHE_MEM_reg[9][29]  ( .D(n12421), .CK(N28803), .Q(n4789), .QN(
        n9612) );
  DFF_X1 \CACHE_MEM_reg[9][28]  ( .D(n12420), .CK(N28803), .Q(n4776), .QN(
        n9628) );
  DFF_X1 \CACHE_MEM_reg[9][27]  ( .D(n12419), .CK(N28803), .Q(n4756), .QN(
        n9644) );
  DFF_X1 \CACHE_MEM_reg[9][26]  ( .D(n12418), .CK(N28803), .Q(n4743), .QN(
        n9660) );
  DFF_X1 \CACHE_MEM_reg[9][25]  ( .D(n12417), .CK(N28803), .Q(n4732), .QN(
        n9676) );
  DFF_X1 \CACHE_MEM_reg[9][24]  ( .D(n12416), .CK(N28803), .Q(n4715), .QN(
        n9692) );
  DFF_X1 \CACHE_MEM_reg[9][23]  ( .D(n12415), .CK(N28803), .Q(n4704), .QN(
        n9708) );
  DFF_X1 \CACHE_MEM_reg[9][22]  ( .D(n12414), .CK(N28803), .Q(n4687), .QN(
        n9724) );
  DFF_X1 \CACHE_MEM_reg[9][21]  ( .D(n12413), .CK(N28803), .Q(n4676), .QN(
        n9740) );
  DFF_X1 \CACHE_MEM_reg[9][20]  ( .D(n12412), .CK(N28803), .Q(n4663), .QN(
        n9756) );
  DFF_X1 \CACHE_MEM_reg[9][19]  ( .D(n12411), .CK(N28803), .Q(n4648), .QN(
        n9772) );
  DFF_X1 \CACHE_MEM_reg[9][18]  ( .D(n12410), .CK(N28803), .Q(n4635), .QN(
        n9788) );
  DFF_X1 \CACHE_MEM_reg[9][17]  ( .D(n12409), .CK(N28803), .Q(n4624), .QN(
        n9804) );
  DFF_X1 \CACHE_MEM_reg[9][16]  ( .D(n12408), .CK(N28803), .Q(n4602), .QN(
        n9820) );
  DFF_X1 \CACHE_MEM_reg[9][15]  ( .D(n12407), .CK(N28803), .Q(n4591), .QN(
        n9836) );
  DFF_X1 \CACHE_MEM_reg[9][14]  ( .D(n12406), .CK(N28803), .Q(n4574), .QN(
        n9852) );
  DFF_X1 \CACHE_MEM_reg[9][13]  ( .D(n12405), .CK(N28803), .Q(n4563), .QN(
        n9868) );
  DFF_X1 \CACHE_MEM_reg[9][12]  ( .D(n12404), .CK(N28803), .Q(n4550), .QN(
        n9884) );
  DFF_X1 \CACHE_MEM_reg[9][11]  ( .D(n12403), .CK(N28803), .Q(n4535), .QN(
        n9900) );
  DFF_X1 \CACHE_MEM_reg[9][10]  ( .D(n12402), .CK(N28803), .Q(n4522), .QN(
        n9916) );
  DFF_X1 \CACHE_MEM_reg[9][9]  ( .D(n12401), .CK(N28803), .Q(n4511), .QN(n9932) );
  DFF_X1 \CACHE_MEM_reg[9][8]  ( .D(n12400), .CK(N28803), .Q(n4494), .QN(n9948) );
  DFF_X1 \CACHE_MEM_reg[9][7]  ( .D(n12399), .CK(N28803), .Q(n4483), .QN(n9964) );
  DFF_X1 \CACHE_MEM_reg[9][6]  ( .D(n12398), .CK(N28803), .Q(n4461), .QN(n9980) );
  DFF_X1 \CACHE_MEM_reg[9][5]  ( .D(n12397), .CK(N28803), .Q(n4450), .QN(n9996) );
  DFF_X1 \CACHE_MEM_reg[9][4]  ( .D(n12396), .CK(N28803), .Q(n4437), .QN(
        n10012) );
  DFF_X1 \CACHE_MEM_reg[9][3]  ( .D(n12395), .CK(N28803), .Q(n4422), .QN(
        n10028) );
  DFF_X1 \CACHE_MEM_reg[9][2]  ( .D(n12394), .CK(N28803), .Q(n4409), .QN(
        n10044) );
  DFF_X1 \CACHE_MEM_reg[9][1]  ( .D(n12393), .CK(N28803), .Q(n4398), .QN(
        n10060) );
  DFF_X1 \CACHE_MEM_reg[9][0]  ( .D(n12392), .CK(N28803), .Q(n4381), .QN(
        n10076) );
  DFF_X1 \CACHE_MEM_reg[8][255]  ( .D(n12391), .CK(N28803), .Q(n1405), .QN(
        n5992) );
  DFF_X1 \CACHE_MEM_reg[8][254]  ( .D(n12390), .CK(N28803), .Q(n1397), .QN(
        n6008) );
  DFF_X1 \CACHE_MEM_reg[8][253]  ( .D(n12389), .CK(N28803), .Q(n1390), .QN(
        n6024) );
  DFF_X1 \CACHE_MEM_reg[8][252]  ( .D(n12388), .CK(N28803), .Q(n1384), .QN(
        n6040) );
  DFF_X1 \CACHE_MEM_reg[8][251]  ( .D(n12387), .CK(N28803), .Q(n1373), .QN(
        n6056) );
  DFF_X1 \CACHE_MEM_reg[8][250]  ( .D(n12386), .CK(N28803), .Q(n1369), .QN(
        n6072) );
  DFF_X1 \CACHE_MEM_reg[8][249]  ( .D(n12385), .CK(N28803), .Q(n1362), .QN(
        n6088) );
  DFF_X1 \CACHE_MEM_reg[8][248]  ( .D(n12384), .CK(N28803), .Q(n1356), .QN(
        n6104) );
  DFF_X1 \CACHE_MEM_reg[8][247]  ( .D(n12383), .CK(N28803), .Q(n1349), .QN(
        n6120) );
  DFF_X1 \CACHE_MEM_reg[8][246]  ( .D(n12382), .CK(N28803), .Q(n1345), .QN(
        n6136) );
  DFF_X1 \CACHE_MEM_reg[8][245]  ( .D(n12381), .CK(N28803), .Q(n1329), .QN(
        n6152) );
  DFF_X1 \CACHE_MEM_reg[8][244]  ( .D(n12380), .CK(N28803), .Q(n1322), .QN(
        n6168) );
  DFF_X1 \CACHE_MEM_reg[8][243]  ( .D(n12379), .CK(N28803), .Q(n1314), .QN(
        n6184) );
  DFF_X1 \CACHE_MEM_reg[8][242]  ( .D(n12378), .CK(N28803), .Q(n1310), .QN(
        n6200) );
  DFF_X1 \CACHE_MEM_reg[8][241]  ( .D(n12377), .CK(N28803), .Q(n1302), .QN(
        n6216) );
  DFF_X1 \CACHE_MEM_reg[8][240]  ( .D(n12376), .CK(N28803), .Q(n1291), .QN(
        n6232) );
  DFF_X1 \CACHE_MEM_reg[8][239]  ( .D(n12375), .CK(N28803), .Q(n1283), .QN(
        n6248) );
  DFF_X1 \CACHE_MEM_reg[8][238]  ( .D(n12374), .CK(N28803), .Q(n1279), .QN(
        n6264) );
  DFF_X1 \CACHE_MEM_reg[8][237]  ( .D(n12373), .CK(N28803), .Q(n1271), .QN(
        n6280) );
  DFF_X1 \CACHE_MEM_reg[8][236]  ( .D(n12372), .CK(N28803), .Q(n1264), .QN(
        n6296) );
  DFF_X1 \CACHE_MEM_reg[8][235]  ( .D(n12371), .CK(N28803), .Q(n1252), .QN(
        n6312) );
  DFF_X1 \CACHE_MEM_reg[8][234]  ( .D(n12370), .CK(N28803), .Q(n1248), .QN(
        n6328) );
  DFF_X1 \CACHE_MEM_reg[8][233]  ( .D(n12369), .CK(N28803), .Q(n1240), .QN(
        n6344) );
  DFF_X1 \CACHE_MEM_reg[8][232]  ( .D(n12368), .CK(N28803), .Q(n1233), .QN(
        n6360) );
  DFF_X1 \CACHE_MEM_reg[8][231]  ( .D(n12367), .CK(N28803), .Q(n1225), .QN(
        n6376) );
  DFF_X1 \CACHE_MEM_reg[8][230]  ( .D(n12366), .CK(N28803), .Q(n1221), .QN(
        n6392) );
  DFF_X1 \CACHE_MEM_reg[8][229]  ( .D(n12365), .CK(N28803), .Q(n1209), .QN(
        n6408) );
  DFF_X1 \CACHE_MEM_reg[8][228]  ( .D(n12364), .CK(N28803), .Q(n1202), .QN(
        n6424) );
  DFF_X1 \CACHE_MEM_reg[8][227]  ( .D(n12363), .CK(N28803), .Q(n1194), .QN(
        n6440) );
  DFF_X1 \CACHE_MEM_reg[8][226]  ( .D(n12362), .CK(N28803), .Q(n1190), .QN(
        n6456) );
  DFF_X1 \CACHE_MEM_reg[8][225]  ( .D(n12361), .CK(N28803), .Q(n1182), .QN(
        n6472) );
  DFF_X1 \CACHE_MEM_reg[8][224]  ( .D(n12360), .CK(N28803), .Q(n172), .QN(
        n6488) );
  DFF_X1 \CACHE_MEM_reg[8][223]  ( .D(n12359), .CK(N28803), .Q(n2875), .QN(
        n6504) );
  DFF_X1 \CACHE_MEM_reg[8][222]  ( .D(n12358), .CK(N28803), .Q(n2860), .QN(
        n6520) );
  DFF_X1 \CACHE_MEM_reg[8][221]  ( .D(n12357), .CK(N28803), .Q(n2847), .QN(
        n6536) );
  DFF_X1 \CACHE_MEM_reg[8][220]  ( .D(n12356), .CK(N28803), .Q(n2836), .QN(
        n6552) );
  DFF_X1 \CACHE_MEM_reg[8][219]  ( .D(n12355), .CK(N28803), .Q(n2814), .QN(
        n6568) );
  DFF_X1 \CACHE_MEM_reg[8][218]  ( .D(n12354), .CK(N28803), .Q(n2803), .QN(
        n6584) );
  DFF_X1 \CACHE_MEM_reg[8][217]  ( .D(n12353), .CK(N28803), .Q(n2786), .QN(
        n6600) );
  DFF_X1 \CACHE_MEM_reg[8][216]  ( .D(n12352), .CK(N28803), .Q(n2775), .QN(
        n6616) );
  DFF_X1 \CACHE_MEM_reg[8][215]  ( .D(n12351), .CK(N28803), .Q(n2762), .QN(
        n6632) );
  DFF_X1 \CACHE_MEM_reg[8][214]  ( .D(n12350), .CK(N28803), .Q(n2747), .QN(
        n6648) );
  DFF_X1 \CACHE_MEM_reg[8][213]  ( .D(n12349), .CK(N28803), .Q(n2734), .QN(
        n6664) );
  DFF_X1 \CACHE_MEM_reg[8][212]  ( .D(n12348), .CK(N28803), .Q(n2723), .QN(
        n6680) );
  DFF_X1 \CACHE_MEM_reg[8][211]  ( .D(n12347), .CK(N28803), .Q(n2706), .QN(
        n6696) );
  DFF_X1 \CACHE_MEM_reg[8][210]  ( .D(n12346), .CK(N28803), .Q(n2695), .QN(
        n6712) );
  DFF_X1 \CACHE_MEM_reg[8][209]  ( .D(n12345), .CK(N28803), .Q(n2673), .QN(
        n6728) );
  DFF_X1 \CACHE_MEM_reg[8][208]  ( .D(n12344), .CK(N28803), .Q(n2665), .QN(
        n6744) );
  DFF_X1 \CACHE_MEM_reg[8][207]  ( .D(n12343), .CK(N28803), .Q(n2654), .QN(
        n6760) );
  DFF_X1 \CACHE_MEM_reg[8][206]  ( .D(n12342), .CK(N28803), .Q(n2637), .QN(
        n6776) );
  DFF_X1 \CACHE_MEM_reg[8][205]  ( .D(n12341), .CK(N28803), .Q(n2626), .QN(
        n6792) );
  DFF_X1 \CACHE_MEM_reg[8][204]  ( .D(n12340), .CK(N28803), .Q(n2613), .QN(
        n6808) );
  DFF_X1 \CACHE_MEM_reg[8][203]  ( .D(n12339), .CK(N28803), .Q(n2598), .QN(
        n6824) );
  DFF_X1 \CACHE_MEM_reg[8][202]  ( .D(n12338), .CK(N28803), .Q(n2585), .QN(
        n6840) );
  DFF_X1 \CACHE_MEM_reg[8][201]  ( .D(n12337), .CK(N28803), .Q(n2574), .QN(
        n6856) );
  DFF_X1 \CACHE_MEM_reg[8][200]  ( .D(n12336), .CK(N28803), .Q(n2557), .QN(
        n6872) );
  DFF_X1 \CACHE_MEM_reg[8][199]  ( .D(n12335), .CK(N28803), .Q(n2546), .QN(
        n6888) );
  DFF_X1 \CACHE_MEM_reg[8][198]  ( .D(n12334), .CK(N28803), .Q(n2524), .QN(
        n6904) );
  DFF_X1 \CACHE_MEM_reg[8][197]  ( .D(n12333), .CK(N28803), .Q(n2513), .QN(
        n6920) );
  DFF_X1 \CACHE_MEM_reg[8][196]  ( .D(n12332), .CK(N28803), .Q(n2500), .QN(
        n6936) );
  DFF_X1 \CACHE_MEM_reg[8][195]  ( .D(n12331), .CK(N28803), .Q(n2485), .QN(
        n6952) );
  DFF_X1 \CACHE_MEM_reg[8][194]  ( .D(n12330), .CK(N28803), .Q(n2472), .QN(
        n6968) );
  DFF_X1 \CACHE_MEM_reg[8][193]  ( .D(n12329), .CK(N28803), .Q(n2461), .QN(
        n6984) );
  DFF_X1 \CACHE_MEM_reg[8][192]  ( .D(n12328), .CK(N28803), .Q(n2444), .QN(
        n7000) );
  DFF_X1 \CACHE_MEM_reg[8][191]  ( .D(n12327), .CK(N28803), .Q(n3319), .QN(
        n7016) );
  DFF_X1 \CACHE_MEM_reg[8][190]  ( .D(n12326), .CK(N28803), .Q(n1398), .QN(
        n7032) );
  DFF_X1 \CACHE_MEM_reg[8][189]  ( .D(n12325), .CK(N28803), .Q(n1392), .QN(
        n7048) );
  DFF_X1 \CACHE_MEM_reg[8][188]  ( .D(n12324), .CK(N28803), .Q(n1385), .QN(
        n7064) );
  DFF_X1 \CACHE_MEM_reg[8][187]  ( .D(n12323), .CK(N28803), .Q(n1381), .QN(
        n7080) );
  DFF_X1 \CACHE_MEM_reg[8][186]  ( .D(n12322), .CK(N28803), .Q(n1370), .QN(
        n7096) );
  DFF_X1 \CACHE_MEM_reg[8][185]  ( .D(n12321), .CK(N28803), .Q(n1364), .QN(
        n7112) );
  DFF_X1 \CACHE_MEM_reg[8][184]  ( .D(n12320), .CK(N28803), .Q(n1357), .QN(
        n7128) );
  DFF_X1 \CACHE_MEM_reg[8][183]  ( .D(n12319), .CK(N28803), .Q(n1353), .QN(
        n7144) );
  DFF_X1 \CACHE_MEM_reg[8][182]  ( .D(n12318), .CK(N28803), .Q(n1346), .QN(
        n7160) );
  DFF_X1 \CACHE_MEM_reg[8][181]  ( .D(n12317), .CK(N28803), .Q(n1331), .QN(
        n7176) );
  DFF_X1 \CACHE_MEM_reg[8][180]  ( .D(n12316), .CK(N28803), .Q(n1323), .QN(
        n7192) );
  DFF_X1 \CACHE_MEM_reg[8][179]  ( .D(n12315), .CK(N28803), .Q(n1319), .QN(
        n7208) );
  DFF_X1 \CACHE_MEM_reg[8][178]  ( .D(n12314), .CK(N28803), .Q(n1311), .QN(
        n7224) );
  DFF_X1 \CACHE_MEM_reg[8][177]  ( .D(n12313), .CK(N28803), .Q(n1304), .QN(
        n7240) );
  DFF_X1 \CACHE_MEM_reg[8][176]  ( .D(n12312), .CK(N28803), .Q(n1292), .QN(
        n7256) );
  DFF_X1 \CACHE_MEM_reg[8][175]  ( .D(n12311), .CK(N28803), .Q(n1288), .QN(
        n7272) );
  DFF_X1 \CACHE_MEM_reg[8][174]  ( .D(n12310), .CK(N28803), .Q(n1280), .QN(
        n7288) );
  DFF_X1 \CACHE_MEM_reg[8][173]  ( .D(n12309), .CK(N28803), .Q(n1273), .QN(
        n7304) );
  DFF_X1 \CACHE_MEM_reg[8][172]  ( .D(n12308), .CK(N28803), .Q(n1265), .QN(
        n7320) );
  DFF_X1 \CACHE_MEM_reg[8][171]  ( .D(n12307), .CK(N28803), .Q(n1261), .QN(
        n7336) );
  DFF_X1 \CACHE_MEM_reg[8][170]  ( .D(n12306), .CK(N28803), .Q(n1249), .QN(
        n7352) );
  DFF_X1 \CACHE_MEM_reg[8][169]  ( .D(n12305), .CK(N28803), .Q(n1242), .QN(
        n7368) );
  DFF_X1 \CACHE_MEM_reg[8][168]  ( .D(n12304), .CK(N28803), .Q(n1234), .QN(
        n7384) );
  DFF_X1 \CACHE_MEM_reg[8][167]  ( .D(n12303), .CK(N28803), .Q(n1230), .QN(
        n7400) );
  DFF_X1 \CACHE_MEM_reg[8][166]  ( .D(n12302), .CK(N28803), .Q(n1222), .QN(
        n7416) );
  DFF_X1 \CACHE_MEM_reg[8][165]  ( .D(n12301), .CK(N28803), .Q(n1211), .QN(
        n7432) );
  DFF_X1 \CACHE_MEM_reg[8][164]  ( .D(n12300), .CK(N28803), .Q(n1203), .QN(
        n7448) );
  DFF_X1 \CACHE_MEM_reg[8][163]  ( .D(n12299), .CK(N28803), .Q(n1199), .QN(
        n7464) );
  DFF_X1 \CACHE_MEM_reg[8][162]  ( .D(n12298), .CK(N28803), .Q(n1191), .QN(
        n7480) );
  DFF_X1 \CACHE_MEM_reg[8][161]  ( .D(n12297), .CK(N28803), .Q(n1184), .QN(
        n7496) );
  DFF_X1 \CACHE_MEM_reg[8][160]  ( .D(n12296), .CK(N28803), .Q(n238), .QN(
        n7512) );
  DFF_X1 \CACHE_MEM_reg[8][159]  ( .D(n12295), .CK(N28803), .Q(n3322), .QN(
        n7528) );
  DFF_X1 \CACHE_MEM_reg[8][158]  ( .D(n12294), .CK(N28803), .Q(n3307), .QN(
        n7544) );
  DFF_X1 \CACHE_MEM_reg[8][157]  ( .D(n12293), .CK(N28803), .Q(n3294), .QN(
        n7560) );
  DFF_X1 \CACHE_MEM_reg[8][156]  ( .D(n12292), .CK(N28803), .Q(n3283), .QN(
        n7576) );
  DFF_X1 \CACHE_MEM_reg[8][155]  ( .D(n12291), .CK(N28803), .Q(n3261), .QN(
        n7592) );
  DFF_X1 \CACHE_MEM_reg[8][154]  ( .D(n12290), .CK(N28803), .Q(n3250), .QN(
        n7608) );
  DFF_X1 \CACHE_MEM_reg[8][153]  ( .D(n12289), .CK(N28803), .Q(n3233), .QN(
        n7624) );
  DFF_X1 \CACHE_MEM_reg[8][152]  ( .D(n12288), .CK(N28803), .Q(n3222), .QN(
        n7640) );
  DFF_X1 \CACHE_MEM_reg[8][151]  ( .D(n12287), .CK(N28803), .Q(n3209), .QN(
        n7656) );
  DFF_X1 \CACHE_MEM_reg[8][150]  ( .D(n12286), .CK(N28803), .Q(n3194), .QN(
        n7672) );
  DFF_X1 \CACHE_MEM_reg[8][149]  ( .D(n12285), .CK(N28803), .Q(n3181), .QN(
        n7688) );
  DFF_X1 \CACHE_MEM_reg[8][148]  ( .D(n12284), .CK(N28803), .Q(n3170), .QN(
        n7704) );
  DFF_X1 \CACHE_MEM_reg[8][147]  ( .D(n12283), .CK(N28803), .Q(n3153), .QN(
        n7720) );
  DFF_X1 \CACHE_MEM_reg[8][146]  ( .D(n12282), .CK(N28803), .Q(n3142), .QN(
        n7736) );
  DFF_X1 \CACHE_MEM_reg[8][145]  ( .D(n12281), .CK(N28803), .Q(n3120), .QN(
        n7752) );
  DFF_X1 \CACHE_MEM_reg[8][144]  ( .D(n12280), .CK(N28803), .Q(n3109), .QN(
        n7768) );
  DFF_X1 \CACHE_MEM_reg[8][143]  ( .D(n12279), .CK(N28803), .Q(n3096), .QN(
        n7784) );
  DFF_X1 \CACHE_MEM_reg[8][142]  ( .D(n12278), .CK(N28803), .Q(n3081), .QN(
        n7800) );
  DFF_X1 \CACHE_MEM_reg[8][141]  ( .D(n12277), .CK(N28803), .Q(n3068), .QN(
        n7816) );
  DFF_X1 \CACHE_MEM_reg[8][140]  ( .D(n12276), .CK(N28803), .Q(n3057), .QN(
        n7832) );
  DFF_X1 \CACHE_MEM_reg[8][139]  ( .D(n12275), .CK(N28803), .Q(n3040), .QN(
        n7848) );
  DFF_X1 \CACHE_MEM_reg[8][138]  ( .D(n12274), .CK(N28803), .Q(n3029), .QN(
        n7864) );
  DFF_X1 \CACHE_MEM_reg[8][137]  ( .D(n12273), .CK(N28803), .Q(n3012), .QN(
        n7880) );
  DFF_X1 \CACHE_MEM_reg[8][136]  ( .D(n12272), .CK(N28803), .Q(n3001), .QN(
        n7896) );
  DFF_X1 \CACHE_MEM_reg[8][135]  ( .D(n12271), .CK(N28803), .Q(n2988), .QN(
        n7912) );
  DFF_X1 \CACHE_MEM_reg[8][134]  ( .D(n12270), .CK(N28803), .Q(n2968), .QN(
        n7928) );
  DFF_X1 \CACHE_MEM_reg[8][133]  ( .D(n12269), .CK(N28803), .Q(n2955), .QN(
        n7944) );
  DFF_X1 \CACHE_MEM_reg[8][132]  ( .D(n12268), .CK(N28803), .Q(n2944), .QN(
        n7960) );
  DFF_X1 \CACHE_MEM_reg[8][131]  ( .D(n12267), .CK(N28803), .Q(n2927), .QN(
        n7976) );
  DFF_X1 \CACHE_MEM_reg[8][130]  ( .D(n12266), .CK(N28803), .Q(n2916), .QN(
        n7992) );
  DFF_X1 \CACHE_MEM_reg[8][129]  ( .D(n12265), .CK(N28803), .Q(n2899), .QN(
        n8008) );
  DFF_X1 \CACHE_MEM_reg[8][128]  ( .D(n12264), .CK(N28803), .Q(n2888), .QN(
        n8024) );
  DFF_X1 \CACHE_MEM_reg[8][127]  ( .D(n12263), .CK(N28803), .Q(n1400), .QN(
        n8040) );
  DFF_X1 \CACHE_MEM_reg[8][126]  ( .D(n12262), .CK(N28803), .Q(n1966), .QN(
        n8056) );
  DFF_X1 \CACHE_MEM_reg[8][125]  ( .D(n12261), .CK(N28803), .Q(n1950), .QN(
        n8072) );
  DFF_X1 \CACHE_MEM_reg[8][124]  ( .D(n12260), .CK(N28803), .Q(n1925), .QN(
        n8088) );
  DFF_X1 \CACHE_MEM_reg[8][123]  ( .D(n12259), .CK(N28803), .Q(n1909), .QN(
        n8104) );
  DFF_X1 \CACHE_MEM_reg[8][122]  ( .D(n12258), .CK(N28803), .Q(n1889), .QN(
        n8120) );
  DFF_X1 \CACHE_MEM_reg[8][121]  ( .D(n12257), .CK(N28803), .Q(n1873), .QN(
        n8136) );
  DFF_X1 \CACHE_MEM_reg[8][120]  ( .D(n12256), .CK(N28803), .Q(n1853), .QN(
        n8152) );
  DFF_X1 \CACHE_MEM_reg[8][119]  ( .D(n12255), .CK(N28803), .Q(n1837), .QN(
        n8168) );
  DFF_X1 \CACHE_MEM_reg[8][118]  ( .D(n12254), .CK(N28803), .Q(n1817), .QN(
        n8184) );
  DFF_X1 \CACHE_MEM_reg[8][117]  ( .D(n12253), .CK(N28803), .Q(n1801), .QN(
        n8200) );
  DFF_X1 \CACHE_MEM_reg[8][116]  ( .D(n12252), .CK(N28803), .Q(n1776), .QN(
        n8216) );
  DFF_X1 \CACHE_MEM_reg[8][115]  ( .D(n12251), .CK(N28803), .Q(n1760), .QN(
        n8232) );
  DFF_X1 \CACHE_MEM_reg[8][114]  ( .D(n12250), .CK(N28803), .Q(n1740), .QN(
        n8248) );
  DFF_X1 \CACHE_MEM_reg[8][113]  ( .D(n12249), .CK(N28803), .Q(n1724), .QN(
        n8264) );
  DFF_X1 \CACHE_MEM_reg[8][112]  ( .D(n12248), .CK(N28803), .Q(n1704), .QN(
        n8280) );
  DFF_X1 \CACHE_MEM_reg[8][111]  ( .D(n12247), .CK(N28803), .Q(n1688), .QN(
        n8296) );
  DFF_X1 \CACHE_MEM_reg[8][110]  ( .D(n12246), .CK(N28803), .Q(n1668), .QN(
        n8312) );
  DFF_X1 \CACHE_MEM_reg[8][109]  ( .D(n12245), .CK(N28803), .Q(n1652), .QN(
        n8328) );
  DFF_X1 \CACHE_MEM_reg[8][108]  ( .D(n12244), .CK(N28803), .Q(n1627), .QN(
        n8344) );
  DFF_X1 \CACHE_MEM_reg[8][107]  ( .D(n12243), .CK(N28803), .Q(n1611), .QN(
        n8360) );
  DFF_X1 \CACHE_MEM_reg[8][106]  ( .D(n12242), .CK(N28803), .Q(n1591), .QN(
        n8376) );
  DFF_X1 \CACHE_MEM_reg[8][105]  ( .D(n12241), .CK(N28803), .Q(n1575), .QN(
        n8392) );
  DFF_X1 \CACHE_MEM_reg[8][104]  ( .D(n12240), .CK(N28803), .Q(n1555), .QN(
        n8408) );
  DFF_X1 \CACHE_MEM_reg[8][103]  ( .D(n12239), .CK(N28803), .Q(n1539), .QN(
        n8424) );
  DFF_X1 \CACHE_MEM_reg[8][102]  ( .D(n12238), .CK(N28803), .Q(n1519), .QN(
        n8440) );
  DFF_X1 \CACHE_MEM_reg[8][101]  ( .D(n12237), .CK(N28803), .Q(n1503), .QN(
        n8456) );
  DFF_X1 \CACHE_MEM_reg[8][100]  ( .D(n12236), .CK(N28803), .Q(n1478), .QN(
        n8472) );
  DFF_X1 \CACHE_MEM_reg[8][99]  ( .D(n12235), .CK(N28803), .Q(n1462), .QN(
        n8488) );
  DFF_X1 \CACHE_MEM_reg[8][98]  ( .D(n12234), .CK(N28803), .Q(n1442), .QN(
        n8504) );
  DFF_X1 \CACHE_MEM_reg[8][97]  ( .D(n12233), .CK(N28803), .Q(n1426), .QN(
        n8520) );
  DFF_X1 \CACHE_MEM_reg[8][96]  ( .D(n12232), .CK(N28803), .Q(n1406), .QN(
        n8536) );
  DFF_X1 \CACHE_MEM_reg[8][95]  ( .D(n12231), .CK(N28803), .Q(n1986), .QN(
        n8552) );
  DFF_X1 \CACHE_MEM_reg[8][94]  ( .D(n12230), .CK(N28803), .Q(n1969), .QN(
        n8568) );
  DFF_X1 \CACHE_MEM_reg[8][93]  ( .D(n12229), .CK(N28803), .Q(n1953), .QN(
        n8584) );
  DFF_X1 \CACHE_MEM_reg[8][92]  ( .D(n12228), .CK(N28803), .Q(n1928), .QN(
        n8600) );
  DFF_X1 \CACHE_MEM_reg[8][91]  ( .D(n12227), .CK(N28803), .Q(n1912), .QN(
        n8616) );
  DFF_X1 \CACHE_MEM_reg[8][90]  ( .D(n12226), .CK(N28803), .Q(n1892), .QN(
        n8632) );
  DFF_X1 \CACHE_MEM_reg[8][89]  ( .D(n12225), .CK(N28803), .Q(n1876), .QN(
        n8648) );
  DFF_X1 \CACHE_MEM_reg[8][88]  ( .D(n12224), .CK(N28803), .Q(n1856), .QN(
        n8664) );
  DFF_X1 \CACHE_MEM_reg[8][87]  ( .D(n12223), .CK(N28803), .Q(n1840), .QN(
        n8680) );
  DFF_X1 \CACHE_MEM_reg[8][86]  ( .D(n12222), .CK(N28803), .Q(n1820), .QN(
        n8696) );
  DFF_X1 \CACHE_MEM_reg[8][85]  ( .D(n12221), .CK(N28803), .Q(n1804), .QN(
        n8712) );
  DFF_X1 \CACHE_MEM_reg[8][84]  ( .D(n12220), .CK(N28803), .Q(n1779), .QN(
        n8728) );
  DFF_X1 \CACHE_MEM_reg[8][83]  ( .D(n12219), .CK(N28803), .Q(n1763), .QN(
        n8744) );
  DFF_X1 \CACHE_MEM_reg[8][82]  ( .D(n12218), .CK(N28803), .Q(n1743), .QN(
        n8760) );
  DFF_X1 \CACHE_MEM_reg[8][81]  ( .D(n12217), .CK(N28803), .Q(n1727), .QN(
        n8776) );
  DFF_X1 \CACHE_MEM_reg[8][80]  ( .D(n12216), .CK(N28803), .Q(n1707), .QN(
        n8792) );
  DFF_X1 \CACHE_MEM_reg[8][79]  ( .D(n12215), .CK(N28803), .Q(n1691), .QN(
        n8808) );
  DFF_X1 \CACHE_MEM_reg[8][78]  ( .D(n12214), .CK(N28803), .Q(n1671), .QN(
        n8824) );
  DFF_X1 \CACHE_MEM_reg[8][77]  ( .D(n12213), .CK(N28803), .Q(n1655), .QN(
        n8840) );
  DFF_X1 \CACHE_MEM_reg[8][76]  ( .D(n12212), .CK(N28803), .Q(n1630), .QN(
        n8856) );
  DFF_X1 \CACHE_MEM_reg[8][75]  ( .D(n12211), .CK(N28803), .Q(n1614), .QN(
        n8872) );
  DFF_X1 \CACHE_MEM_reg[8][74]  ( .D(n12210), .CK(N28803), .Q(n1594), .QN(
        n8888) );
  DFF_X1 \CACHE_MEM_reg[8][73]  ( .D(n12209), .CK(N28803), .Q(n1578), .QN(
        n8904) );
  DFF_X1 \CACHE_MEM_reg[8][72]  ( .D(n12208), .CK(N28803), .Q(n1558), .QN(
        n8920) );
  DFF_X1 \CACHE_MEM_reg[8][71]  ( .D(n12207), .CK(N28803), .Q(n1542), .QN(
        n8936) );
  DFF_X1 \CACHE_MEM_reg[8][70]  ( .D(n12206), .CK(N28803), .Q(n1522), .QN(
        n8952) );
  DFF_X1 \CACHE_MEM_reg[8][69]  ( .D(n12205), .CK(N28803), .Q(n1506), .QN(
        n8968) );
  DFF_X1 \CACHE_MEM_reg[8][68]  ( .D(n12204), .CK(N28803), .Q(n1481), .QN(
        n8984) );
  DFF_X1 \CACHE_MEM_reg[8][67]  ( .D(n12203), .CK(N28803), .Q(n1465), .QN(
        n9000) );
  DFF_X1 \CACHE_MEM_reg[8][66]  ( .D(n12202), .CK(N28803), .Q(n1445), .QN(
        n9016) );
  DFF_X1 \CACHE_MEM_reg[8][65]  ( .D(n12201), .CK(N28803), .Q(n1429), .QN(
        n9032) );
  DFF_X1 \CACHE_MEM_reg[8][64]  ( .D(n12200), .CK(N28803), .Q(n1409), .QN(
        n9048) );
  DFF_X1 \CACHE_MEM_reg[8][63]  ( .D(n12199), .CK(N28803), .Q(n1401), .QN(
        n9064) );
  DFF_X1 \CACHE_MEM_reg[8][62]  ( .D(n12198), .CK(N28803), .Q(n1393), .QN(
        n9080) );
  DFF_X1 \CACHE_MEM_reg[8][61]  ( .D(n12197), .CK(N28803), .Q(n1389), .QN(
        n9096) );
  DFF_X1 \CACHE_MEM_reg[8][60]  ( .D(n12196), .CK(N28803), .Q(n1382), .QN(
        n9112) );
  DFF_X1 \CACHE_MEM_reg[8][59]  ( .D(n12195), .CK(N28803), .Q(n1372), .QN(
        n9128) );
  DFF_X1 \CACHE_MEM_reg[8][58]  ( .D(n12194), .CK(N28803), .Q(n1365), .QN(
        n9144) );
  DFF_X1 \CACHE_MEM_reg[8][57]  ( .D(n12193), .CK(N28803), .Q(n1361), .QN(
        n9160) );
  DFF_X1 \CACHE_MEM_reg[8][56]  ( .D(n12192), .CK(N28803), .Q(n1354), .QN(
        n9176) );
  DFF_X1 \CACHE_MEM_reg[8][55]  ( .D(n12191), .CK(N28803), .Q(n1348), .QN(
        n9192) );
  DFF_X1 \CACHE_MEM_reg[8][54]  ( .D(n12190), .CK(N28803), .Q(n1332), .QN(
        n9208) );
  DFF_X1 \CACHE_MEM_reg[8][53]  ( .D(n12189), .CK(N28803), .Q(n1328), .QN(
        n9224) );
  DFF_X1 \CACHE_MEM_reg[8][52]  ( .D(n12188), .CK(N28803), .Q(n1320), .QN(
        n9240) );
  DFF_X1 \CACHE_MEM_reg[8][51]  ( .D(n12187), .CK(N28803), .Q(n1313), .QN(
        n9256) );
  DFF_X1 \CACHE_MEM_reg[8][50]  ( .D(n12186), .CK(N28803), .Q(n1305), .QN(
        n9272) );
  DFF_X1 \CACHE_MEM_reg[8][49]  ( .D(n12185), .CK(N28803), .Q(n1301), .QN(
        n9288) );
  DFF_X1 \CACHE_MEM_reg[8][48]  ( .D(n12184), .CK(N28803), .Q(n1289), .QN(
        n9304) );
  DFF_X1 \CACHE_MEM_reg[8][47]  ( .D(n12183), .CK(N28803), .Q(n1282), .QN(
        n9320) );
  DFF_X1 \CACHE_MEM_reg[8][46]  ( .D(n12182), .CK(N28803), .Q(n1274), .QN(
        n9336) );
  DFF_X1 \CACHE_MEM_reg[8][45]  ( .D(n12181), .CK(N28803), .Q(n1270), .QN(
        n9352) );
  DFF_X1 \CACHE_MEM_reg[8][44]  ( .D(n12180), .CK(N28803), .Q(n1262), .QN(
        n9368) );
  DFF_X1 \CACHE_MEM_reg[8][43]  ( .D(n12179), .CK(N28803), .Q(n1251), .QN(
        n9384) );
  DFF_X1 \CACHE_MEM_reg[8][42]  ( .D(n12178), .CK(N28803), .Q(n1243), .QN(
        n9400) );
  DFF_X1 \CACHE_MEM_reg[8][41]  ( .D(n12177), .CK(N28803), .Q(n1239), .QN(
        n9416) );
  DFF_X1 \CACHE_MEM_reg[8][40]  ( .D(n12176), .CK(N28803), .Q(n1231), .QN(
        n9432) );
  DFF_X1 \CACHE_MEM_reg[8][39]  ( .D(n12175), .CK(N28803), .Q(n1224), .QN(
        n9448) );
  DFF_X1 \CACHE_MEM_reg[8][38]  ( .D(n12174), .CK(N28803), .Q(n1212), .QN(
        n9464) );
  DFF_X1 \CACHE_MEM_reg[8][37]  ( .D(n12173), .CK(N28803), .Q(n1208), .QN(
        n9480) );
  DFF_X1 \CACHE_MEM_reg[8][36]  ( .D(n12172), .CK(N28803), .Q(n1200), .QN(
        n9496) );
  DFF_X1 \CACHE_MEM_reg[8][35]  ( .D(n12171), .CK(N28803), .Q(n1193), .QN(
        n9512) );
  DFF_X1 \CACHE_MEM_reg[8][34]  ( .D(n12170), .CK(N28803), .Q(n1185), .QN(
        n9528) );
  DFF_X1 \CACHE_MEM_reg[8][33]  ( .D(n12169), .CK(N28803), .Q(n1181), .QN(
        n9544) );
  DFF_X1 \CACHE_MEM_reg[8][32]  ( .D(n12168), .CK(N28803), .Q(n170), .QN(n9560) );
  DFF_X1 \CACHE_MEM_reg[8][31]  ( .D(n12167), .CK(N28803), .Q(n2433), .QN(
        n9576) );
  DFF_X1 \CACHE_MEM_reg[8][30]  ( .D(n12166), .CK(N28803), .Q(n2416), .QN(
        n9592) );
  DFF_X1 \CACHE_MEM_reg[8][29]  ( .D(n12165), .CK(N28803), .Q(n2405), .QN(
        n9608) );
  DFF_X1 \CACHE_MEM_reg[8][28]  ( .D(n12164), .CK(N28803), .Q(n2392), .QN(
        n9624) );
  DFF_X1 \CACHE_MEM_reg[8][27]  ( .D(n12163), .CK(N28803), .Q(n2372), .QN(
        n9640) );
  DFF_X1 \CACHE_MEM_reg[8][26]  ( .D(n12162), .CK(N28803), .Q(n2359), .QN(
        n9656) );
  DFF_X1 \CACHE_MEM_reg[8][25]  ( .D(n12161), .CK(N28803), .Q(n2348), .QN(
        n9672) );
  DFF_X1 \CACHE_MEM_reg[8][24]  ( .D(n12160), .CK(N28803), .Q(n2331), .QN(
        n9688) );
  DFF_X1 \CACHE_MEM_reg[8][23]  ( .D(n12159), .CK(N28803), .Q(n2320), .QN(
        n9704) );
  DFF_X1 \CACHE_MEM_reg[8][22]  ( .D(n12158), .CK(N28803), .Q(n2303), .QN(
        n9720) );
  DFF_X1 \CACHE_MEM_reg[8][21]  ( .D(n12157), .CK(N28803), .Q(n2292), .QN(
        n9736) );
  DFF_X1 \CACHE_MEM_reg[8][20]  ( .D(n12156), .CK(N28803), .Q(n2279), .QN(
        n9752) );
  DFF_X1 \CACHE_MEM_reg[8][19]  ( .D(n12155), .CK(N28803), .Q(n2264), .QN(
        n9768) );
  DFF_X1 \CACHE_MEM_reg[8][18]  ( .D(n12154), .CK(N28803), .Q(n2251), .QN(
        n9784) );
  DFF_X1 \CACHE_MEM_reg[8][17]  ( .D(n12153), .CK(N28803), .Q(n2240), .QN(
        n9800) );
  DFF_X1 \CACHE_MEM_reg[8][16]  ( .D(n12152), .CK(N28803), .Q(n2218), .QN(
        n9816) );
  DFF_X1 \CACHE_MEM_reg[8][15]  ( .D(n12151), .CK(N28803), .Q(n2207), .QN(
        n9832) );
  DFF_X1 \CACHE_MEM_reg[8][14]  ( .D(n12150), .CK(N28803), .Q(n2190), .QN(
        n9848) );
  DFF_X1 \CACHE_MEM_reg[8][13]  ( .D(n12149), .CK(N28803), .Q(n2179), .QN(
        n9864) );
  DFF_X1 \CACHE_MEM_reg[8][12]  ( .D(n12148), .CK(N28803), .Q(n2166), .QN(
        n9880) );
  DFF_X1 \CACHE_MEM_reg[8][11]  ( .D(n12147), .CK(N28803), .Q(n2151), .QN(
        n9896) );
  DFF_X1 \CACHE_MEM_reg[8][10]  ( .D(n12146), .CK(N28803), .Q(n2138), .QN(
        n9912) );
  DFF_X1 \CACHE_MEM_reg[8][9]  ( .D(n12145), .CK(N28803), .Q(n2127), .QN(n9928) );
  DFF_X1 \CACHE_MEM_reg[8][8]  ( .D(n12144), .CK(N28803), .Q(n2110), .QN(n9944) );
  DFF_X1 \CACHE_MEM_reg[8][7]  ( .D(n12143), .CK(N28803), .Q(n2099), .QN(n9960) );
  DFF_X1 \CACHE_MEM_reg[8][6]  ( .D(n12142), .CK(N28803), .Q(n2077), .QN(n9976) );
  DFF_X1 \CACHE_MEM_reg[8][5]  ( .D(n12141), .CK(N28803), .Q(n2066), .QN(n9992) );
  DFF_X1 \CACHE_MEM_reg[8][4]  ( .D(n12140), .CK(N28803), .Q(n2053), .QN(
        n10008) );
  DFF_X1 \CACHE_MEM_reg[8][3]  ( .D(n12139), .CK(N28803), .Q(n2038), .QN(
        n10024) );
  DFF_X1 \CACHE_MEM_reg[8][2]  ( .D(n12138), .CK(N28803), .Q(n2025), .QN(
        n10040) );
  DFF_X1 \CACHE_MEM_reg[8][1]  ( .D(n12137), .CK(N28803), .Q(n2014), .QN(
        n10056) );
  DFF_X1 \CACHE_MEM_reg[8][0]  ( .D(n12136), .CK(N28803), .Q(n1997), .QN(
        n10072) );
  DFF_X1 \CACHE_MEM_reg[7][255]  ( .D(n12135), .CK(N28803), .QN(n6007) );
  DFF_X1 \CACHE_MEM_reg[7][254]  ( .D(n12134), .CK(N28803), .QN(n6023) );
  DFF_X1 \CACHE_MEM_reg[7][253]  ( .D(n12133), .CK(N28803), .QN(n6039) );
  DFF_X1 \CACHE_MEM_reg[7][252]  ( .D(n12132), .CK(N28803), .QN(n6055) );
  DFF_X1 \CACHE_MEM_reg[7][251]  ( .D(n12131), .CK(N28803), .QN(n6071) );
  DFF_X1 \CACHE_MEM_reg[7][250]  ( .D(n12130), .CK(N28803), .QN(n6087) );
  DFF_X1 \CACHE_MEM_reg[7][249]  ( .D(n12129), .CK(N28803), .QN(n6103) );
  DFF_X1 \CACHE_MEM_reg[7][248]  ( .D(n12128), .CK(N28803), .QN(n6119) );
  DFF_X1 \CACHE_MEM_reg[7][247]  ( .D(n12127), .CK(N28803), .QN(n6135) );
  DFF_X1 \CACHE_MEM_reg[7][246]  ( .D(n12126), .CK(N28803), .QN(n6151) );
  DFF_X1 \CACHE_MEM_reg[7][245]  ( .D(n12125), .CK(N28803), .QN(n6167) );
  DFF_X1 \CACHE_MEM_reg[7][244]  ( .D(n12124), .CK(N28803), .QN(n6183) );
  DFF_X1 \CACHE_MEM_reg[7][243]  ( .D(n12123), .CK(N28803), .QN(n6199) );
  DFF_X1 \CACHE_MEM_reg[7][242]  ( .D(n12122), .CK(N28803), .QN(n6215) );
  DFF_X1 \CACHE_MEM_reg[7][241]  ( .D(n12121), .CK(N28803), .QN(n6231) );
  DFF_X1 \CACHE_MEM_reg[7][240]  ( .D(n12120), .CK(N28803), .QN(n6247) );
  DFF_X1 \CACHE_MEM_reg[7][239]  ( .D(n12119), .CK(N28803), .QN(n6263) );
  DFF_X1 \CACHE_MEM_reg[7][238]  ( .D(n12118), .CK(N28803), .QN(n6279) );
  DFF_X1 \CACHE_MEM_reg[7][237]  ( .D(n12117), .CK(N28803), .QN(n6295) );
  DFF_X1 \CACHE_MEM_reg[7][236]  ( .D(n12116), .CK(N28803), .QN(n6311) );
  DFF_X1 \CACHE_MEM_reg[7][235]  ( .D(n12115), .CK(N28803), .QN(n6327) );
  DFF_X1 \CACHE_MEM_reg[7][234]  ( .D(n12114), .CK(N28803), .QN(n6343) );
  DFF_X1 \CACHE_MEM_reg[7][233]  ( .D(n12113), .CK(N28803), .QN(n6359) );
  DFF_X1 \CACHE_MEM_reg[7][232]  ( .D(n12112), .CK(N28803), .QN(n6375) );
  DFF_X1 \CACHE_MEM_reg[7][231]  ( .D(n12111), .CK(N28803), .QN(n6391) );
  DFF_X1 \CACHE_MEM_reg[7][230]  ( .D(n12110), .CK(N28803), .QN(n6407) );
  DFF_X1 \CACHE_MEM_reg[7][229]  ( .D(n12109), .CK(N28803), .QN(n6423) );
  DFF_X1 \CACHE_MEM_reg[7][228]  ( .D(n12108), .CK(N28803), .QN(n6439) );
  DFF_X1 \CACHE_MEM_reg[7][227]  ( .D(n12107), .CK(N28803), .QN(n6455) );
  DFF_X1 \CACHE_MEM_reg[7][226]  ( .D(n12106), .CK(N28803), .QN(n6471) );
  DFF_X1 \CACHE_MEM_reg[7][225]  ( .D(n12105), .CK(N28803), .QN(n6487) );
  DFF_X1 \CACHE_MEM_reg[7][224]  ( .D(n12104), .CK(N28803), .QN(n6503) );
  DFF_X1 \CACHE_MEM_reg[7][223]  ( .D(n12103), .CK(N28803), .QN(n6519) );
  DFF_X1 \CACHE_MEM_reg[7][222]  ( .D(n12102), .CK(N28803), .QN(n6535) );
  DFF_X1 \CACHE_MEM_reg[7][221]  ( .D(n12101), .CK(N28803), .QN(n6551) );
  DFF_X1 \CACHE_MEM_reg[7][220]  ( .D(n12100), .CK(N28803), .QN(n6567) );
  DFF_X1 \CACHE_MEM_reg[7][219]  ( .D(n12099), .CK(N28803), .QN(n6583) );
  DFF_X1 \CACHE_MEM_reg[7][218]  ( .D(n12098), .CK(N28803), .QN(n6599) );
  DFF_X1 \CACHE_MEM_reg[7][217]  ( .D(n12097), .CK(N28803), .QN(n6615) );
  DFF_X1 \CACHE_MEM_reg[7][216]  ( .D(n12096), .CK(N28803), .QN(n6631) );
  DFF_X1 \CACHE_MEM_reg[7][215]  ( .D(n12095), .CK(N28803), .QN(n6647) );
  DFF_X1 \CACHE_MEM_reg[7][214]  ( .D(n12094), .CK(N28803), .QN(n6663) );
  DFF_X1 \CACHE_MEM_reg[7][213]  ( .D(n12093), .CK(N28803), .QN(n6679) );
  DFF_X1 \CACHE_MEM_reg[7][212]  ( .D(n12092), .CK(N28803), .QN(n6695) );
  DFF_X1 \CACHE_MEM_reg[7][211]  ( .D(n12091), .CK(N28803), .QN(n6711) );
  DFF_X1 \CACHE_MEM_reg[7][210]  ( .D(n12090), .CK(N28803), .QN(n6727) );
  DFF_X1 \CACHE_MEM_reg[7][209]  ( .D(n12089), .CK(N28803), .QN(n6743) );
  DFF_X1 \CACHE_MEM_reg[7][208]  ( .D(n12088), .CK(N28803), .QN(n6759) );
  DFF_X1 \CACHE_MEM_reg[7][207]  ( .D(n12087), .CK(N28803), .QN(n6775) );
  DFF_X1 \CACHE_MEM_reg[7][206]  ( .D(n12086), .CK(N28803), .QN(n6791) );
  DFF_X1 \CACHE_MEM_reg[7][205]  ( .D(n12085), .CK(N28803), .QN(n6807) );
  DFF_X1 \CACHE_MEM_reg[7][204]  ( .D(n12084), .CK(N28803), .QN(n6823) );
  DFF_X1 \CACHE_MEM_reg[7][203]  ( .D(n12083), .CK(N28803), .QN(n6839) );
  DFF_X1 \CACHE_MEM_reg[7][202]  ( .D(n12082), .CK(N28803), .QN(n6855) );
  DFF_X1 \CACHE_MEM_reg[7][201]  ( .D(n12081), .CK(N28803), .QN(n6871) );
  DFF_X1 \CACHE_MEM_reg[7][200]  ( .D(n12080), .CK(N28803), .QN(n6887) );
  DFF_X1 \CACHE_MEM_reg[7][199]  ( .D(n12079), .CK(N28803), .QN(n6903) );
  DFF_X1 \CACHE_MEM_reg[7][198]  ( .D(n12078), .CK(N28803), .QN(n6919) );
  DFF_X1 \CACHE_MEM_reg[7][197]  ( .D(n12077), .CK(N28803), .QN(n6935) );
  DFF_X1 \CACHE_MEM_reg[7][196]  ( .D(n12076), .CK(N28803), .QN(n6951) );
  DFF_X1 \CACHE_MEM_reg[7][195]  ( .D(n12075), .CK(N28803), .QN(n6967) );
  DFF_X1 \CACHE_MEM_reg[7][194]  ( .D(n12074), .CK(N28803), .QN(n6983) );
  DFF_X1 \CACHE_MEM_reg[7][193]  ( .D(n12073), .CK(N28803), .QN(n6999) );
  DFF_X1 \CACHE_MEM_reg[7][192]  ( .D(n12072), .CK(N28803), .QN(n7015) );
  DFF_X1 \CACHE_MEM_reg[7][191]  ( .D(n12071), .CK(N28803), .QN(n7031) );
  DFF_X1 \CACHE_MEM_reg[7][190]  ( .D(n12070), .CK(N28803), .QN(n7047) );
  DFF_X1 \CACHE_MEM_reg[7][189]  ( .D(n12069), .CK(N28803), .QN(n7063) );
  DFF_X1 \CACHE_MEM_reg[7][188]  ( .D(n12068), .CK(N28803), .QN(n7079) );
  DFF_X1 \CACHE_MEM_reg[7][187]  ( .D(n12067), .CK(N28803), .QN(n7095) );
  DFF_X1 \CACHE_MEM_reg[7][186]  ( .D(n12066), .CK(N28803), .QN(n7111) );
  DFF_X1 \CACHE_MEM_reg[7][185]  ( .D(n12065), .CK(N28803), .QN(n7127) );
  DFF_X1 \CACHE_MEM_reg[7][184]  ( .D(n12064), .CK(N28803), .QN(n7143) );
  DFF_X1 \CACHE_MEM_reg[7][183]  ( .D(n12063), .CK(N28803), .QN(n7159) );
  DFF_X1 \CACHE_MEM_reg[7][182]  ( .D(n12062), .CK(N28803), .QN(n7175) );
  DFF_X1 \CACHE_MEM_reg[7][181]  ( .D(n12061), .CK(N28803), .QN(n7191) );
  DFF_X1 \CACHE_MEM_reg[7][180]  ( .D(n12060), .CK(N28803), .QN(n7207) );
  DFF_X1 \CACHE_MEM_reg[7][179]  ( .D(n12059), .CK(N28803), .QN(n7223) );
  DFF_X1 \CACHE_MEM_reg[7][178]  ( .D(n12058), .CK(N28803), .QN(n7239) );
  DFF_X1 \CACHE_MEM_reg[7][177]  ( .D(n12057), .CK(N28803), .QN(n7255) );
  DFF_X1 \CACHE_MEM_reg[7][176]  ( .D(n12056), .CK(N28803), .QN(n7271) );
  DFF_X1 \CACHE_MEM_reg[7][175]  ( .D(n12055), .CK(N28803), .QN(n7287) );
  DFF_X1 \CACHE_MEM_reg[7][174]  ( .D(n12054), .CK(N28803), .QN(n7303) );
  DFF_X1 \CACHE_MEM_reg[7][173]  ( .D(n12053), .CK(N28803), .QN(n7319) );
  DFF_X1 \CACHE_MEM_reg[7][172]  ( .D(n12052), .CK(N28803), .QN(n7335) );
  DFF_X1 \CACHE_MEM_reg[7][171]  ( .D(n12051), .CK(N28803), .QN(n7351) );
  DFF_X1 \CACHE_MEM_reg[7][170]  ( .D(n12050), .CK(N28803), .QN(n7367) );
  DFF_X1 \CACHE_MEM_reg[7][169]  ( .D(n12049), .CK(N28803), .QN(n7383) );
  DFF_X1 \CACHE_MEM_reg[7][168]  ( .D(n12048), .CK(N28803), .QN(n7399) );
  DFF_X1 \CACHE_MEM_reg[7][167]  ( .D(n12047), .CK(N28803), .QN(n7415) );
  DFF_X1 \CACHE_MEM_reg[7][166]  ( .D(n12046), .CK(N28803), .QN(n7431) );
  DFF_X1 \CACHE_MEM_reg[7][165]  ( .D(n12045), .CK(N28803), .QN(n7447) );
  DFF_X1 \CACHE_MEM_reg[7][164]  ( .D(n12044), .CK(N28803), .QN(n7463) );
  DFF_X1 \CACHE_MEM_reg[7][163]  ( .D(n12043), .CK(N28803), .QN(n7479) );
  DFF_X1 \CACHE_MEM_reg[7][162]  ( .D(n12042), .CK(N28803), .QN(n7495) );
  DFF_X1 \CACHE_MEM_reg[7][161]  ( .D(n12041), .CK(N28803), .QN(n7511) );
  DFF_X1 \CACHE_MEM_reg[7][160]  ( .D(n12040), .CK(N28803), .QN(n7527) );
  DFF_X1 \CACHE_MEM_reg[7][159]  ( .D(n12039), .CK(N28803), .QN(n7543) );
  DFF_X1 \CACHE_MEM_reg[7][158]  ( .D(n12038), .CK(N28803), .QN(n7559) );
  DFF_X1 \CACHE_MEM_reg[7][157]  ( .D(n12037), .CK(N28803), .QN(n7575) );
  DFF_X1 \CACHE_MEM_reg[7][156]  ( .D(n12036), .CK(N28803), .QN(n7591) );
  DFF_X1 \CACHE_MEM_reg[7][155]  ( .D(n12035), .CK(N28803), .QN(n7607) );
  DFF_X1 \CACHE_MEM_reg[7][154]  ( .D(n12034), .CK(N28803), .QN(n7623) );
  DFF_X1 \CACHE_MEM_reg[7][153]  ( .D(n12033), .CK(N28803), .QN(n7639) );
  DFF_X1 \CACHE_MEM_reg[7][152]  ( .D(n12032), .CK(N28803), .QN(n7655) );
  DFF_X1 \CACHE_MEM_reg[7][151]  ( .D(n12031), .CK(N28803), .QN(n7671) );
  DFF_X1 \CACHE_MEM_reg[7][150]  ( .D(n12030), .CK(N28803), .QN(n7687) );
  DFF_X1 \CACHE_MEM_reg[7][149]  ( .D(n12029), .CK(N28803), .QN(n7703) );
  DFF_X1 \CACHE_MEM_reg[7][148]  ( .D(n12028), .CK(N28803), .QN(n7719) );
  DFF_X1 \CACHE_MEM_reg[7][147]  ( .D(n12027), .CK(N28803), .QN(n7735) );
  DFF_X1 \CACHE_MEM_reg[7][146]  ( .D(n12026), .CK(N28803), .QN(n7751) );
  DFF_X1 \CACHE_MEM_reg[7][145]  ( .D(n12025), .CK(N28803), .QN(n7767) );
  DFF_X1 \CACHE_MEM_reg[7][144]  ( .D(n12024), .CK(N28803), .QN(n7783) );
  DFF_X1 \CACHE_MEM_reg[7][143]  ( .D(n12023), .CK(N28803), .QN(n7799) );
  DFF_X1 \CACHE_MEM_reg[7][142]  ( .D(n12022), .CK(N28803), .QN(n7815) );
  DFF_X1 \CACHE_MEM_reg[7][141]  ( .D(n12021), .CK(N28803), .QN(n7831) );
  DFF_X1 \CACHE_MEM_reg[7][140]  ( .D(n12020), .CK(N28803), .QN(n7847) );
  DFF_X1 \CACHE_MEM_reg[7][139]  ( .D(n12019), .CK(N28803), .QN(n7863) );
  DFF_X1 \CACHE_MEM_reg[7][138]  ( .D(n12018), .CK(N28803), .QN(n7879) );
  DFF_X1 \CACHE_MEM_reg[7][137]  ( .D(n12017), .CK(N28803), .QN(n7895) );
  DFF_X1 \CACHE_MEM_reg[7][136]  ( .D(n12016), .CK(N28803), .QN(n7911) );
  DFF_X1 \CACHE_MEM_reg[7][135]  ( .D(n12015), .CK(N28803), .QN(n7927) );
  DFF_X1 \CACHE_MEM_reg[7][134]  ( .D(n12014), .CK(N28803), .QN(n7943) );
  DFF_X1 \CACHE_MEM_reg[7][133]  ( .D(n12013), .CK(N28803), .QN(n7959) );
  DFF_X1 \CACHE_MEM_reg[7][132]  ( .D(n12012), .CK(N28803), .QN(n7975) );
  DFF_X1 \CACHE_MEM_reg[7][131]  ( .D(n12011), .CK(N28803), .QN(n7991) );
  DFF_X1 \CACHE_MEM_reg[7][130]  ( .D(n12010), .CK(N28803), .QN(n8007) );
  DFF_X1 \CACHE_MEM_reg[7][129]  ( .D(n12009), .CK(N28803), .QN(n8023) );
  DFF_X1 \CACHE_MEM_reg[7][128]  ( .D(n12008), .CK(N28803), .QN(n8039) );
  DFF_X1 \CACHE_MEM_reg[7][127]  ( .D(n12007), .CK(N28803), .QN(n8055) );
  DFF_X1 \CACHE_MEM_reg[7][126]  ( .D(n12006), .CK(N28803), .QN(n8071) );
  DFF_X1 \CACHE_MEM_reg[7][125]  ( .D(n12005), .CK(N28803), .QN(n8087) );
  DFF_X1 \CACHE_MEM_reg[7][124]  ( .D(n12004), .CK(N28803), .QN(n8103) );
  DFF_X1 \CACHE_MEM_reg[7][123]  ( .D(n12003), .CK(N28803), .QN(n8119) );
  DFF_X1 \CACHE_MEM_reg[7][122]  ( .D(n12002), .CK(N28803), .QN(n8135) );
  DFF_X1 \CACHE_MEM_reg[7][121]  ( .D(n12001), .CK(N28803), .QN(n8151) );
  DFF_X1 \CACHE_MEM_reg[7][120]  ( .D(n12000), .CK(N28803), .QN(n8167) );
  DFF_X1 \CACHE_MEM_reg[7][119]  ( .D(n11999), .CK(N28803), .QN(n8183) );
  DFF_X1 \CACHE_MEM_reg[7][118]  ( .D(n11998), .CK(N28803), .QN(n8199) );
  DFF_X1 \CACHE_MEM_reg[7][117]  ( .D(n11997), .CK(N28803), .QN(n8215) );
  DFF_X1 \CACHE_MEM_reg[7][116]  ( .D(n11996), .CK(N28803), .QN(n8231) );
  DFF_X1 \CACHE_MEM_reg[7][115]  ( .D(n11995), .CK(N28803), .QN(n8247) );
  DFF_X1 \CACHE_MEM_reg[7][114]  ( .D(n11994), .CK(N28803), .QN(n8263) );
  DFF_X1 \CACHE_MEM_reg[7][113]  ( .D(n11993), .CK(N28803), .QN(n8279) );
  DFF_X1 \CACHE_MEM_reg[7][112]  ( .D(n11992), .CK(N28803), .QN(n8295) );
  DFF_X1 \CACHE_MEM_reg[7][111]  ( .D(n11991), .CK(N28803), .QN(n8311) );
  DFF_X1 \CACHE_MEM_reg[7][110]  ( .D(n11990), .CK(N28803), .QN(n8327) );
  DFF_X1 \CACHE_MEM_reg[7][109]  ( .D(n11989), .CK(N28803), .QN(n8343) );
  DFF_X1 \CACHE_MEM_reg[7][108]  ( .D(n11988), .CK(N28803), .QN(n8359) );
  DFF_X1 \CACHE_MEM_reg[7][107]  ( .D(n11987), .CK(N28803), .QN(n8375) );
  DFF_X1 \CACHE_MEM_reg[7][106]  ( .D(n11986), .CK(N28803), .QN(n8391) );
  DFF_X1 \CACHE_MEM_reg[7][105]  ( .D(n11985), .CK(N28803), .QN(n8407) );
  DFF_X1 \CACHE_MEM_reg[7][104]  ( .D(n11984), .CK(N28803), .QN(n8423) );
  DFF_X1 \CACHE_MEM_reg[7][103]  ( .D(n11983), .CK(N28803), .QN(n8439) );
  DFF_X1 \CACHE_MEM_reg[7][102]  ( .D(n11982), .CK(N28803), .QN(n8455) );
  DFF_X1 \CACHE_MEM_reg[7][101]  ( .D(n11981), .CK(N28803), .QN(n8471) );
  DFF_X1 \CACHE_MEM_reg[7][100]  ( .D(n11980), .CK(N28803), .QN(n8487) );
  DFF_X1 \CACHE_MEM_reg[7][99]  ( .D(n11979), .CK(N28803), .QN(n8503) );
  DFF_X1 \CACHE_MEM_reg[7][98]  ( .D(n11978), .CK(N28803), .QN(n8519) );
  DFF_X1 \CACHE_MEM_reg[7][97]  ( .D(n11977), .CK(N28803), .QN(n8535) );
  DFF_X1 \CACHE_MEM_reg[7][96]  ( .D(n11976), .CK(N28803), .QN(n8551) );
  DFF_X1 \CACHE_MEM_reg[7][95]  ( .D(n11975), .CK(N28803), .QN(n8567) );
  DFF_X1 \CACHE_MEM_reg[7][94]  ( .D(n11974), .CK(N28803), .QN(n8583) );
  DFF_X1 \CACHE_MEM_reg[7][93]  ( .D(n11973), .CK(N28803), .QN(n8599) );
  DFF_X1 \CACHE_MEM_reg[7][92]  ( .D(n11972), .CK(N28803), .QN(n8615) );
  DFF_X1 \CACHE_MEM_reg[7][91]  ( .D(n11971), .CK(N28803), .QN(n8631) );
  DFF_X1 \CACHE_MEM_reg[7][90]  ( .D(n11970), .CK(N28803), .QN(n8647) );
  DFF_X1 \CACHE_MEM_reg[7][89]  ( .D(n11969), .CK(N28803), .QN(n8663) );
  DFF_X1 \CACHE_MEM_reg[7][88]  ( .D(n11968), .CK(N28803), .QN(n8679) );
  DFF_X1 \CACHE_MEM_reg[7][87]  ( .D(n11967), .CK(N28803), .QN(n8695) );
  DFF_X1 \CACHE_MEM_reg[7][86]  ( .D(n11966), .CK(N28803), .QN(n8711) );
  DFF_X1 \CACHE_MEM_reg[7][85]  ( .D(n11965), .CK(N28803), .QN(n8727) );
  DFF_X1 \CACHE_MEM_reg[7][84]  ( .D(n11964), .CK(N28803), .QN(n8743) );
  DFF_X1 \CACHE_MEM_reg[7][83]  ( .D(n11963), .CK(N28803), .QN(n8759) );
  DFF_X1 \CACHE_MEM_reg[7][82]  ( .D(n11962), .CK(N28803), .QN(n8775) );
  DFF_X1 \CACHE_MEM_reg[7][81]  ( .D(n11961), .CK(N28803), .QN(n8791) );
  DFF_X1 \CACHE_MEM_reg[7][80]  ( .D(n11960), .CK(N28803), .QN(n8807) );
  DFF_X1 \CACHE_MEM_reg[7][79]  ( .D(n11959), .CK(N28803), .QN(n8823) );
  DFF_X1 \CACHE_MEM_reg[7][78]  ( .D(n11958), .CK(N28803), .QN(n8839) );
  DFF_X1 \CACHE_MEM_reg[7][77]  ( .D(n11957), .CK(N28803), .QN(n8855) );
  DFF_X1 \CACHE_MEM_reg[7][76]  ( .D(n11956), .CK(N28803), .QN(n8871) );
  DFF_X1 \CACHE_MEM_reg[7][75]  ( .D(n11955), .CK(N28803), .QN(n8887) );
  DFF_X1 \CACHE_MEM_reg[7][74]  ( .D(n11954), .CK(N28803), .QN(n8903) );
  DFF_X1 \CACHE_MEM_reg[7][73]  ( .D(n11953), .CK(N28803), .QN(n8919) );
  DFF_X1 \CACHE_MEM_reg[7][72]  ( .D(n11952), .CK(N28803), .QN(n8935) );
  DFF_X1 \CACHE_MEM_reg[7][71]  ( .D(n11951), .CK(N28803), .QN(n8951) );
  DFF_X1 \CACHE_MEM_reg[7][70]  ( .D(n11950), .CK(N28803), .QN(n8967) );
  DFF_X1 \CACHE_MEM_reg[7][69]  ( .D(n11949), .CK(N28803), .QN(n8983) );
  DFF_X1 \CACHE_MEM_reg[7][68]  ( .D(n11948), .CK(N28803), .QN(n8999) );
  DFF_X1 \CACHE_MEM_reg[7][67]  ( .D(n11947), .CK(N28803), .QN(n9015) );
  DFF_X1 \CACHE_MEM_reg[7][66]  ( .D(n11946), .CK(N28803), .QN(n9031) );
  DFF_X1 \CACHE_MEM_reg[7][65]  ( .D(n11945), .CK(N28803), .QN(n9047) );
  DFF_X1 \CACHE_MEM_reg[7][64]  ( .D(n11944), .CK(N28803), .QN(n9063) );
  DFF_X1 \CACHE_MEM_reg[7][63]  ( .D(n11943), .CK(N28803), .QN(n9079) );
  DFF_X1 \CACHE_MEM_reg[7][62]  ( .D(n11942), .CK(N28803), .QN(n9095) );
  DFF_X1 \CACHE_MEM_reg[7][61]  ( .D(n11941), .CK(N28803), .QN(n9111) );
  DFF_X1 \CACHE_MEM_reg[7][60]  ( .D(n11940), .CK(N28803), .QN(n9127) );
  DFF_X1 \CACHE_MEM_reg[7][59]  ( .D(n11939), .CK(N28803), .QN(n9143) );
  DFF_X1 \CACHE_MEM_reg[7][58]  ( .D(n11938), .CK(N28803), .QN(n9159) );
  DFF_X1 \CACHE_MEM_reg[7][57]  ( .D(n11937), .CK(N28803), .QN(n9175) );
  DFF_X1 \CACHE_MEM_reg[7][56]  ( .D(n11936), .CK(N28803), .QN(n9191) );
  DFF_X1 \CACHE_MEM_reg[7][55]  ( .D(n11935), .CK(N28803), .QN(n9207) );
  DFF_X1 \CACHE_MEM_reg[7][54]  ( .D(n11934), .CK(N28803), .QN(n9223) );
  DFF_X1 \CACHE_MEM_reg[7][53]  ( .D(n11933), .CK(N28803), .QN(n9239) );
  DFF_X1 \CACHE_MEM_reg[7][52]  ( .D(n11932), .CK(N28803), .QN(n9255) );
  DFF_X1 \CACHE_MEM_reg[7][51]  ( .D(n11931), .CK(N28803), .QN(n9271) );
  DFF_X1 \CACHE_MEM_reg[7][50]  ( .D(n11930), .CK(N28803), .QN(n9287) );
  DFF_X1 \CACHE_MEM_reg[7][49]  ( .D(n11929), .CK(N28803), .QN(n9303) );
  DFF_X1 \CACHE_MEM_reg[7][48]  ( .D(n11928), .CK(N28803), .QN(n9319) );
  DFF_X1 \CACHE_MEM_reg[7][47]  ( .D(n11927), .CK(N28803), .QN(n9335) );
  DFF_X1 \CACHE_MEM_reg[7][46]  ( .D(n11926), .CK(N28803), .QN(n9351) );
  DFF_X1 \CACHE_MEM_reg[7][45]  ( .D(n11925), .CK(N28803), .QN(n9367) );
  DFF_X1 \CACHE_MEM_reg[7][44]  ( .D(n11924), .CK(N28803), .QN(n9383) );
  DFF_X1 \CACHE_MEM_reg[7][43]  ( .D(n11923), .CK(N28803), .QN(n9399) );
  DFF_X1 \CACHE_MEM_reg[7][42]  ( .D(n11922), .CK(N28803), .QN(n9415) );
  DFF_X1 \CACHE_MEM_reg[7][41]  ( .D(n11921), .CK(N28803), .QN(n9431) );
  DFF_X1 \CACHE_MEM_reg[7][40]  ( .D(n11920), .CK(N28803), .QN(n9447) );
  DFF_X1 \CACHE_MEM_reg[7][39]  ( .D(n11919), .CK(N28803), .QN(n9463) );
  DFF_X1 \CACHE_MEM_reg[7][38]  ( .D(n11918), .CK(N28803), .QN(n9479) );
  DFF_X1 \CACHE_MEM_reg[7][37]  ( .D(n11917), .CK(N28803), .QN(n9495) );
  DFF_X1 \CACHE_MEM_reg[7][36]  ( .D(n11916), .CK(N28803), .QN(n9511) );
  DFF_X1 \CACHE_MEM_reg[7][35]  ( .D(n11915), .CK(N28803), .QN(n9527) );
  DFF_X1 \CACHE_MEM_reg[7][34]  ( .D(n11914), .CK(N28803), .QN(n9543) );
  DFF_X1 \CACHE_MEM_reg[7][33]  ( .D(n11913), .CK(N28803), .QN(n9559) );
  DFF_X1 \CACHE_MEM_reg[7][32]  ( .D(n11912), .CK(N28803), .QN(n9575) );
  DFF_X1 \CACHE_MEM_reg[7][31]  ( .D(n11911), .CK(N28803), .QN(n9591) );
  DFF_X1 \CACHE_MEM_reg[7][30]  ( .D(n11910), .CK(N28803), .QN(n9607) );
  DFF_X1 \CACHE_MEM_reg[7][29]  ( .D(n11909), .CK(N28803), .QN(n9623) );
  DFF_X1 \CACHE_MEM_reg[7][28]  ( .D(n11908), .CK(N28803), .QN(n9639) );
  DFF_X1 \CACHE_MEM_reg[7][27]  ( .D(n11907), .CK(N28803), .QN(n9655) );
  DFF_X1 \CACHE_MEM_reg[7][26]  ( .D(n11906), .CK(N28803), .QN(n9671) );
  DFF_X1 \CACHE_MEM_reg[7][25]  ( .D(n11905), .CK(N28803), .QN(n9687) );
  DFF_X1 \CACHE_MEM_reg[7][24]  ( .D(n11904), .CK(N28803), .QN(n9703) );
  DFF_X1 \CACHE_MEM_reg[7][23]  ( .D(n11903), .CK(N28803), .QN(n9719) );
  DFF_X1 \CACHE_MEM_reg[7][22]  ( .D(n11902), .CK(N28803), .QN(n9735) );
  DFF_X1 \CACHE_MEM_reg[7][21]  ( .D(n11901), .CK(N28803), .QN(n9751) );
  DFF_X1 \CACHE_MEM_reg[7][20]  ( .D(n11900), .CK(N28803), .QN(n9767) );
  DFF_X1 \CACHE_MEM_reg[7][19]  ( .D(n11899), .CK(N28803), .QN(n9783) );
  DFF_X1 \CACHE_MEM_reg[7][18]  ( .D(n11898), .CK(N28803), .QN(n9799) );
  DFF_X1 \CACHE_MEM_reg[7][17]  ( .D(n11897), .CK(N28803), .QN(n9815) );
  DFF_X1 \CACHE_MEM_reg[7][16]  ( .D(n11896), .CK(N28803), .QN(n9831) );
  DFF_X1 \CACHE_MEM_reg[7][15]  ( .D(n11895), .CK(N28803), .QN(n9847) );
  DFF_X1 \CACHE_MEM_reg[7][14]  ( .D(n11894), .CK(N28803), .QN(n9863) );
  DFF_X1 \CACHE_MEM_reg[7][13]  ( .D(n11893), .CK(N28803), .QN(n9879) );
  DFF_X1 \CACHE_MEM_reg[7][12]  ( .D(n11892), .CK(N28803), .QN(n9895) );
  DFF_X1 \CACHE_MEM_reg[7][11]  ( .D(n11891), .CK(N28803), .QN(n9911) );
  DFF_X1 \CACHE_MEM_reg[7][10]  ( .D(n11890), .CK(N28803), .QN(n9927) );
  DFF_X1 \CACHE_MEM_reg[7][9]  ( .D(n11889), .CK(N28803), .QN(n9943) );
  DFF_X1 \CACHE_MEM_reg[7][8]  ( .D(n11888), .CK(N28803), .QN(n9959) );
  DFF_X1 \CACHE_MEM_reg[7][7]  ( .D(n11887), .CK(N28803), .QN(n9975) );
  DFF_X1 \CACHE_MEM_reg[7][6]  ( .D(n11886), .CK(N28803), .QN(n9991) );
  DFF_X1 \CACHE_MEM_reg[7][5]  ( .D(n11885), .CK(N28803), .QN(n10007) );
  DFF_X1 \CACHE_MEM_reg[7][4]  ( .D(n11884), .CK(N28803), .QN(n10023) );
  DFF_X1 \CACHE_MEM_reg[7][3]  ( .D(n11883), .CK(N28803), .QN(n10039) );
  DFF_X1 \CACHE_MEM_reg[7][2]  ( .D(n11882), .CK(N28803), .QN(n10055) );
  DFF_X1 \CACHE_MEM_reg[7][1]  ( .D(n11881), .CK(N28803), .QN(n10071) );
  DFF_X1 \CACHE_MEM_reg[7][0]  ( .D(n11880), .CK(N28803), .QN(n10087) );
  DFF_X1 \CACHE_MEM_reg[6][255]  ( .D(n11879), .CK(N28803), .QN(n6003) );
  DFF_X1 \CACHE_MEM_reg[6][254]  ( .D(n11878), .CK(N28803), .QN(n6019) );
  DFF_X1 \CACHE_MEM_reg[6][253]  ( .D(n11877), .CK(N28803), .QN(n6035) );
  DFF_X1 \CACHE_MEM_reg[6][252]  ( .D(n11876), .CK(N28803), .QN(n6051) );
  DFF_X1 \CACHE_MEM_reg[6][251]  ( .D(n11875), .CK(N28803), .QN(n6067) );
  DFF_X1 \CACHE_MEM_reg[6][250]  ( .D(n11874), .CK(N28803), .QN(n6083) );
  DFF_X1 \CACHE_MEM_reg[6][249]  ( .D(n11873), .CK(N28803), .QN(n6099) );
  DFF_X1 \CACHE_MEM_reg[6][248]  ( .D(n11872), .CK(N28803), .QN(n6115) );
  DFF_X1 \CACHE_MEM_reg[6][247]  ( .D(n11871), .CK(N28803), .QN(n6131) );
  DFF_X1 \CACHE_MEM_reg[6][246]  ( .D(n11870), .CK(N28803), .QN(n6147) );
  DFF_X1 \CACHE_MEM_reg[6][245]  ( .D(n11869), .CK(N28803), .QN(n6163) );
  DFF_X1 \CACHE_MEM_reg[6][244]  ( .D(n11868), .CK(N28803), .QN(n6179) );
  DFF_X1 \CACHE_MEM_reg[6][243]  ( .D(n11867), .CK(N28803), .QN(n6195) );
  DFF_X1 \CACHE_MEM_reg[6][242]  ( .D(n11866), .CK(N28803), .QN(n6211) );
  DFF_X1 \CACHE_MEM_reg[6][241]  ( .D(n11865), .CK(N28803), .QN(n6227) );
  DFF_X1 \CACHE_MEM_reg[6][240]  ( .D(n11864), .CK(N28803), .QN(n6243) );
  DFF_X1 \CACHE_MEM_reg[6][239]  ( .D(n11863), .CK(N28803), .QN(n6259) );
  DFF_X1 \CACHE_MEM_reg[6][238]  ( .D(n11862), .CK(N28803), .QN(n6275) );
  DFF_X1 \CACHE_MEM_reg[6][237]  ( .D(n11861), .CK(N28803), .QN(n6291) );
  DFF_X1 \CACHE_MEM_reg[6][236]  ( .D(n11860), .CK(N28803), .QN(n6307) );
  DFF_X1 \CACHE_MEM_reg[6][235]  ( .D(n11859), .CK(N28803), .QN(n6323) );
  DFF_X1 \CACHE_MEM_reg[6][234]  ( .D(n11858), .CK(N28803), .QN(n6339) );
  DFF_X1 \CACHE_MEM_reg[6][233]  ( .D(n11857), .CK(N28803), .QN(n6355) );
  DFF_X1 \CACHE_MEM_reg[6][232]  ( .D(n11856), .CK(N28803), .QN(n6371) );
  DFF_X1 \CACHE_MEM_reg[6][231]  ( .D(n11855), .CK(N28803), .QN(n6387) );
  DFF_X1 \CACHE_MEM_reg[6][230]  ( .D(n11854), .CK(N28803), .QN(n6403) );
  DFF_X1 \CACHE_MEM_reg[6][229]  ( .D(n11853), .CK(N28803), .QN(n6419) );
  DFF_X1 \CACHE_MEM_reg[6][228]  ( .D(n11852), .CK(N28803), .QN(n6435) );
  DFF_X1 \CACHE_MEM_reg[6][227]  ( .D(n11851), .CK(N28803), .QN(n6451) );
  DFF_X1 \CACHE_MEM_reg[6][226]  ( .D(n11850), .CK(N28803), .QN(n6467) );
  DFF_X1 \CACHE_MEM_reg[6][225]  ( .D(n11849), .CK(N28803), .QN(n6483) );
  DFF_X1 \CACHE_MEM_reg[6][224]  ( .D(n11848), .CK(N28803), .QN(n6499) );
  DFF_X1 \CACHE_MEM_reg[6][223]  ( .D(n11847), .CK(N28803), .QN(n6515) );
  DFF_X1 \CACHE_MEM_reg[6][222]  ( .D(n11846), .CK(N28803), .QN(n6531) );
  DFF_X1 \CACHE_MEM_reg[6][221]  ( .D(n11845), .CK(N28803), .QN(n6547) );
  DFF_X1 \CACHE_MEM_reg[6][220]  ( .D(n11844), .CK(N28803), .QN(n6563) );
  DFF_X1 \CACHE_MEM_reg[6][219]  ( .D(n11843), .CK(N28803), .QN(n6579) );
  DFF_X1 \CACHE_MEM_reg[6][218]  ( .D(n11842), .CK(N28803), .QN(n6595) );
  DFF_X1 \CACHE_MEM_reg[6][217]  ( .D(n11841), .CK(N28803), .QN(n6611) );
  DFF_X1 \CACHE_MEM_reg[6][216]  ( .D(n11840), .CK(N28803), .QN(n6627) );
  DFF_X1 \CACHE_MEM_reg[6][215]  ( .D(n11839), .CK(N28803), .QN(n6643) );
  DFF_X1 \CACHE_MEM_reg[6][214]  ( .D(n11838), .CK(N28803), .QN(n6659) );
  DFF_X1 \CACHE_MEM_reg[6][213]  ( .D(n11837), .CK(N28803), .QN(n6675) );
  DFF_X1 \CACHE_MEM_reg[6][212]  ( .D(n11836), .CK(N28803), .QN(n6691) );
  DFF_X1 \CACHE_MEM_reg[6][211]  ( .D(n11835), .CK(N28803), .QN(n6707) );
  DFF_X1 \CACHE_MEM_reg[6][210]  ( .D(n11834), .CK(N28803), .QN(n6723) );
  DFF_X1 \CACHE_MEM_reg[6][209]  ( .D(n11833), .CK(N28803), .QN(n6739) );
  DFF_X1 \CACHE_MEM_reg[6][208]  ( .D(n11832), .CK(N28803), .QN(n6755) );
  DFF_X1 \CACHE_MEM_reg[6][207]  ( .D(n11831), .CK(N28803), .QN(n6771) );
  DFF_X1 \CACHE_MEM_reg[6][206]  ( .D(n11830), .CK(N28803), .QN(n6787) );
  DFF_X1 \CACHE_MEM_reg[6][205]  ( .D(n11829), .CK(N28803), .QN(n6803) );
  DFF_X1 \CACHE_MEM_reg[6][204]  ( .D(n11828), .CK(N28803), .QN(n6819) );
  DFF_X1 \CACHE_MEM_reg[6][203]  ( .D(n11827), .CK(N28803), .QN(n6835) );
  DFF_X1 \CACHE_MEM_reg[6][202]  ( .D(n11826), .CK(N28803), .QN(n6851) );
  DFF_X1 \CACHE_MEM_reg[6][201]  ( .D(n11825), .CK(N28803), .QN(n6867) );
  DFF_X1 \CACHE_MEM_reg[6][200]  ( .D(n11824), .CK(N28803), .QN(n6883) );
  DFF_X1 \CACHE_MEM_reg[6][199]  ( .D(n11823), .CK(N28803), .QN(n6899) );
  DFF_X1 \CACHE_MEM_reg[6][198]  ( .D(n11822), .CK(N28803), .QN(n6915) );
  DFF_X1 \CACHE_MEM_reg[6][197]  ( .D(n11821), .CK(N28803), .QN(n6931) );
  DFF_X1 \CACHE_MEM_reg[6][196]  ( .D(n11820), .CK(N28803), .QN(n6947) );
  DFF_X1 \CACHE_MEM_reg[6][195]  ( .D(n11819), .CK(N28803), .QN(n6963) );
  DFF_X1 \CACHE_MEM_reg[6][194]  ( .D(n11818), .CK(N28803), .QN(n6979) );
  DFF_X1 \CACHE_MEM_reg[6][193]  ( .D(n11817), .CK(N28803), .QN(n6995) );
  DFF_X1 \CACHE_MEM_reg[6][192]  ( .D(n11816), .CK(N28803), .QN(n7011) );
  DFF_X1 \CACHE_MEM_reg[6][191]  ( .D(n11815), .CK(N28803), .QN(n7027) );
  DFF_X1 \CACHE_MEM_reg[6][190]  ( .D(n11814), .CK(N28803), .QN(n7043) );
  DFF_X1 \CACHE_MEM_reg[6][189]  ( .D(n11813), .CK(N28803), .QN(n7059) );
  DFF_X1 \CACHE_MEM_reg[6][188]  ( .D(n11812), .CK(N28803), .QN(n7075) );
  DFF_X1 \CACHE_MEM_reg[6][187]  ( .D(n11811), .CK(N28803), .QN(n7091) );
  DFF_X1 \CACHE_MEM_reg[6][186]  ( .D(n11810), .CK(N28803), .QN(n7107) );
  DFF_X1 \CACHE_MEM_reg[6][185]  ( .D(n11809), .CK(N28803), .QN(n7123) );
  DFF_X1 \CACHE_MEM_reg[6][184]  ( .D(n11808), .CK(N28803), .QN(n7139) );
  DFF_X1 \CACHE_MEM_reg[6][183]  ( .D(n11807), .CK(N28803), .QN(n7155) );
  DFF_X1 \CACHE_MEM_reg[6][182]  ( .D(n11806), .CK(N28803), .QN(n7171) );
  DFF_X1 \CACHE_MEM_reg[6][181]  ( .D(n11805), .CK(N28803), .QN(n7187) );
  DFF_X1 \CACHE_MEM_reg[6][180]  ( .D(n11804), .CK(N28803), .QN(n7203) );
  DFF_X1 \CACHE_MEM_reg[6][179]  ( .D(n11803), .CK(N28803), .QN(n7219) );
  DFF_X1 \CACHE_MEM_reg[6][178]  ( .D(n11802), .CK(N28803), .QN(n7235) );
  DFF_X1 \CACHE_MEM_reg[6][177]  ( .D(n11801), .CK(N28803), .QN(n7251) );
  DFF_X1 \CACHE_MEM_reg[6][176]  ( .D(n11800), .CK(N28803), .QN(n7267) );
  DFF_X1 \CACHE_MEM_reg[6][175]  ( .D(n11799), .CK(N28803), .QN(n7283) );
  DFF_X1 \CACHE_MEM_reg[6][174]  ( .D(n11798), .CK(N28803), .QN(n7299) );
  DFF_X1 \CACHE_MEM_reg[6][173]  ( .D(n11797), .CK(N28803), .QN(n7315) );
  DFF_X1 \CACHE_MEM_reg[6][172]  ( .D(n11796), .CK(N28803), .QN(n7331) );
  DFF_X1 \CACHE_MEM_reg[6][171]  ( .D(n11795), .CK(N28803), .QN(n7347) );
  DFF_X1 \CACHE_MEM_reg[6][170]  ( .D(n11794), .CK(N28803), .QN(n7363) );
  DFF_X1 \CACHE_MEM_reg[6][169]  ( .D(n11793), .CK(N28803), .QN(n7379) );
  DFF_X1 \CACHE_MEM_reg[6][168]  ( .D(n11792), .CK(N28803), .QN(n7395) );
  DFF_X1 \CACHE_MEM_reg[6][167]  ( .D(n11791), .CK(N28803), .QN(n7411) );
  DFF_X1 \CACHE_MEM_reg[6][166]  ( .D(n11790), .CK(N28803), .QN(n7427) );
  DFF_X1 \CACHE_MEM_reg[6][165]  ( .D(n11789), .CK(N28803), .QN(n7443) );
  DFF_X1 \CACHE_MEM_reg[6][164]  ( .D(n11788), .CK(N28803), .QN(n7459) );
  DFF_X1 \CACHE_MEM_reg[6][163]  ( .D(n11787), .CK(N28803), .QN(n7475) );
  DFF_X1 \CACHE_MEM_reg[6][162]  ( .D(n11786), .CK(N28803), .QN(n7491) );
  DFF_X1 \CACHE_MEM_reg[6][161]  ( .D(n11785), .CK(N28803), .QN(n7507) );
  DFF_X1 \CACHE_MEM_reg[6][160]  ( .D(n11784), .CK(N28803), .QN(n7523) );
  DFF_X1 \CACHE_MEM_reg[6][159]  ( .D(n11783), .CK(N28803), .QN(n7539) );
  DFF_X1 \CACHE_MEM_reg[6][158]  ( .D(n11782), .CK(N28803), .QN(n7555) );
  DFF_X1 \CACHE_MEM_reg[6][157]  ( .D(n11781), .CK(N28803), .QN(n7571) );
  DFF_X1 \CACHE_MEM_reg[6][156]  ( .D(n11780), .CK(N28803), .QN(n7587) );
  DFF_X1 \CACHE_MEM_reg[6][155]  ( .D(n11779), .CK(N28803), .QN(n7603) );
  DFF_X1 \CACHE_MEM_reg[6][154]  ( .D(n11778), .CK(N28803), .QN(n7619) );
  DFF_X1 \CACHE_MEM_reg[6][153]  ( .D(n11777), .CK(N28803), .QN(n7635) );
  DFF_X1 \CACHE_MEM_reg[6][152]  ( .D(n11776), .CK(N28803), .QN(n7651) );
  DFF_X1 \CACHE_MEM_reg[6][151]  ( .D(n11775), .CK(N28803), .QN(n7667) );
  DFF_X1 \CACHE_MEM_reg[6][150]  ( .D(n11774), .CK(N28803), .QN(n7683) );
  DFF_X1 \CACHE_MEM_reg[6][149]  ( .D(n11773), .CK(N28803), .QN(n7699) );
  DFF_X1 \CACHE_MEM_reg[6][148]  ( .D(n11772), .CK(N28803), .QN(n7715) );
  DFF_X1 \CACHE_MEM_reg[6][147]  ( .D(n11771), .CK(N28803), .QN(n7731) );
  DFF_X1 \CACHE_MEM_reg[6][146]  ( .D(n11770), .CK(N28803), .QN(n7747) );
  DFF_X1 \CACHE_MEM_reg[6][145]  ( .D(n11769), .CK(N28803), .QN(n7763) );
  DFF_X1 \CACHE_MEM_reg[6][144]  ( .D(n11768), .CK(N28803), .QN(n7779) );
  DFF_X1 \CACHE_MEM_reg[6][143]  ( .D(n11767), .CK(N28803), .QN(n7795) );
  DFF_X1 \CACHE_MEM_reg[6][142]  ( .D(n11766), .CK(N28803), .QN(n7811) );
  DFF_X1 \CACHE_MEM_reg[6][141]  ( .D(n11765), .CK(N28803), .QN(n7827) );
  DFF_X1 \CACHE_MEM_reg[6][140]  ( .D(n11764), .CK(N28803), .QN(n7843) );
  DFF_X1 \CACHE_MEM_reg[6][139]  ( .D(n11763), .CK(N28803), .QN(n7859) );
  DFF_X1 \CACHE_MEM_reg[6][138]  ( .D(n11762), .CK(N28803), .QN(n7875) );
  DFF_X1 \CACHE_MEM_reg[6][137]  ( .D(n11761), .CK(N28803), .QN(n7891) );
  DFF_X1 \CACHE_MEM_reg[6][136]  ( .D(n11760), .CK(N28803), .QN(n7907) );
  DFF_X1 \CACHE_MEM_reg[6][135]  ( .D(n11759), .CK(N28803), .QN(n7923) );
  DFF_X1 \CACHE_MEM_reg[6][134]  ( .D(n11758), .CK(N28803), .QN(n7939) );
  DFF_X1 \CACHE_MEM_reg[6][133]  ( .D(n11757), .CK(N28803), .QN(n7955) );
  DFF_X1 \CACHE_MEM_reg[6][132]  ( .D(n11756), .CK(N28803), .QN(n7971) );
  DFF_X1 \CACHE_MEM_reg[6][131]  ( .D(n11755), .CK(N28803), .QN(n7987) );
  DFF_X1 \CACHE_MEM_reg[6][130]  ( .D(n11754), .CK(N28803), .QN(n8003) );
  DFF_X1 \CACHE_MEM_reg[6][129]  ( .D(n11753), .CK(N28803), .QN(n8019) );
  DFF_X1 \CACHE_MEM_reg[6][128]  ( .D(n11752), .CK(N28803), .QN(n8035) );
  DFF_X1 \CACHE_MEM_reg[6][127]  ( .D(n11751), .CK(N28803), .QN(n8051) );
  DFF_X1 \CACHE_MEM_reg[6][126]  ( .D(n11750), .CK(N28803), .QN(n8067) );
  DFF_X1 \CACHE_MEM_reg[6][125]  ( .D(n11749), .CK(N28803), .QN(n8083) );
  DFF_X1 \CACHE_MEM_reg[6][124]  ( .D(n11748), .CK(N28803), .QN(n8099) );
  DFF_X1 \CACHE_MEM_reg[6][123]  ( .D(n11747), .CK(N28803), .QN(n8115) );
  DFF_X1 \CACHE_MEM_reg[6][122]  ( .D(n11746), .CK(N28803), .QN(n8131) );
  DFF_X1 \CACHE_MEM_reg[6][121]  ( .D(n11745), .CK(N28803), .QN(n8147) );
  DFF_X1 \CACHE_MEM_reg[6][120]  ( .D(n11744), .CK(N28803), .QN(n8163) );
  DFF_X1 \CACHE_MEM_reg[6][119]  ( .D(n11743), .CK(N28803), .QN(n8179) );
  DFF_X1 \CACHE_MEM_reg[6][118]  ( .D(n11742), .CK(N28803), .QN(n8195) );
  DFF_X1 \CACHE_MEM_reg[6][117]  ( .D(n11741), .CK(N28803), .QN(n8211) );
  DFF_X1 \CACHE_MEM_reg[6][116]  ( .D(n11740), .CK(N28803), .QN(n8227) );
  DFF_X1 \CACHE_MEM_reg[6][115]  ( .D(n11739), .CK(N28803), .QN(n8243) );
  DFF_X1 \CACHE_MEM_reg[6][114]  ( .D(n11738), .CK(N28803), .QN(n8259) );
  DFF_X1 \CACHE_MEM_reg[6][113]  ( .D(n11737), .CK(N28803), .QN(n8275) );
  DFF_X1 \CACHE_MEM_reg[6][112]  ( .D(n11736), .CK(N28803), .QN(n8291) );
  DFF_X1 \CACHE_MEM_reg[6][111]  ( .D(n11735), .CK(N28803), .QN(n8307) );
  DFF_X1 \CACHE_MEM_reg[6][110]  ( .D(n11734), .CK(N28803), .QN(n8323) );
  DFF_X1 \CACHE_MEM_reg[6][109]  ( .D(n11733), .CK(N28803), .QN(n8339) );
  DFF_X1 \CACHE_MEM_reg[6][108]  ( .D(n11732), .CK(N28803), .QN(n8355) );
  DFF_X1 \CACHE_MEM_reg[6][107]  ( .D(n11731), .CK(N28803), .QN(n8371) );
  DFF_X1 \CACHE_MEM_reg[6][106]  ( .D(n11730), .CK(N28803), .QN(n8387) );
  DFF_X1 \CACHE_MEM_reg[6][105]  ( .D(n11729), .CK(N28803), .QN(n8403) );
  DFF_X1 \CACHE_MEM_reg[6][104]  ( .D(n11728), .CK(N28803), .QN(n8419) );
  DFF_X1 \CACHE_MEM_reg[6][103]  ( .D(n11727), .CK(N28803), .QN(n8435) );
  DFF_X1 \CACHE_MEM_reg[6][102]  ( .D(n11726), .CK(N28803), .QN(n8451) );
  DFF_X1 \CACHE_MEM_reg[6][101]  ( .D(n11725), .CK(N28803), .QN(n8467) );
  DFF_X1 \CACHE_MEM_reg[6][100]  ( .D(n11724), .CK(N28803), .QN(n8483) );
  DFF_X1 \CACHE_MEM_reg[6][99]  ( .D(n11723), .CK(N28803), .QN(n8499) );
  DFF_X1 \CACHE_MEM_reg[6][98]  ( .D(n11722), .CK(N28803), .QN(n8515) );
  DFF_X1 \CACHE_MEM_reg[6][97]  ( .D(n11721), .CK(N28803), .QN(n8531) );
  DFF_X1 \CACHE_MEM_reg[6][96]  ( .D(n11720), .CK(N28803), .QN(n8547) );
  DFF_X1 \CACHE_MEM_reg[6][95]  ( .D(n11719), .CK(N28803), .QN(n8563) );
  DFF_X1 \CACHE_MEM_reg[6][94]  ( .D(n11718), .CK(N28803), .QN(n8579) );
  DFF_X1 \CACHE_MEM_reg[6][93]  ( .D(n11717), .CK(N28803), .QN(n8595) );
  DFF_X1 \CACHE_MEM_reg[6][92]  ( .D(n11716), .CK(N28803), .QN(n8611) );
  DFF_X1 \CACHE_MEM_reg[6][91]  ( .D(n11715), .CK(N28803), .QN(n8627) );
  DFF_X1 \CACHE_MEM_reg[6][90]  ( .D(n11714), .CK(N28803), .QN(n8643) );
  DFF_X1 \CACHE_MEM_reg[6][89]  ( .D(n11713), .CK(N28803), .QN(n8659) );
  DFF_X1 \CACHE_MEM_reg[6][88]  ( .D(n11712), .CK(N28803), .QN(n8675) );
  DFF_X1 \CACHE_MEM_reg[6][87]  ( .D(n11711), .CK(N28803), .QN(n8691) );
  DFF_X1 \CACHE_MEM_reg[6][86]  ( .D(n11710), .CK(N28803), .QN(n8707) );
  DFF_X1 \CACHE_MEM_reg[6][85]  ( .D(n11709), .CK(N28803), .QN(n8723) );
  DFF_X1 \CACHE_MEM_reg[6][84]  ( .D(n11708), .CK(N28803), .QN(n8739) );
  DFF_X1 \CACHE_MEM_reg[6][83]  ( .D(n11707), .CK(N28803), .QN(n8755) );
  DFF_X1 \CACHE_MEM_reg[6][82]  ( .D(n11706), .CK(N28803), .QN(n8771) );
  DFF_X1 \CACHE_MEM_reg[6][81]  ( .D(n11705), .CK(N28803), .QN(n8787) );
  DFF_X1 \CACHE_MEM_reg[6][80]  ( .D(n11704), .CK(N28803), .QN(n8803) );
  DFF_X1 \CACHE_MEM_reg[6][79]  ( .D(n11703), .CK(N28803), .QN(n8819) );
  DFF_X1 \CACHE_MEM_reg[6][78]  ( .D(n11702), .CK(N28803), .QN(n8835) );
  DFF_X1 \CACHE_MEM_reg[6][77]  ( .D(n11701), .CK(N28803), .QN(n8851) );
  DFF_X1 \CACHE_MEM_reg[6][76]  ( .D(n11700), .CK(N28803), .QN(n8867) );
  DFF_X1 \CACHE_MEM_reg[6][75]  ( .D(n11699), .CK(N28803), .QN(n8883) );
  DFF_X1 \CACHE_MEM_reg[6][74]  ( .D(n11698), .CK(N28803), .QN(n8899) );
  DFF_X1 \CACHE_MEM_reg[6][73]  ( .D(n11697), .CK(N28803), .QN(n8915) );
  DFF_X1 \CACHE_MEM_reg[6][72]  ( .D(n11696), .CK(N28803), .QN(n8931) );
  DFF_X1 \CACHE_MEM_reg[6][71]  ( .D(n11695), .CK(N28803), .QN(n8947) );
  DFF_X1 \CACHE_MEM_reg[6][70]  ( .D(n11694), .CK(N28803), .QN(n8963) );
  DFF_X1 \CACHE_MEM_reg[6][69]  ( .D(n11693), .CK(N28803), .QN(n8979) );
  DFF_X1 \CACHE_MEM_reg[6][68]  ( .D(n11692), .CK(N28803), .QN(n8995) );
  DFF_X1 \CACHE_MEM_reg[6][67]  ( .D(n11691), .CK(N28803), .QN(n9011) );
  DFF_X1 \CACHE_MEM_reg[6][66]  ( .D(n11690), .CK(N28803), .QN(n9027) );
  DFF_X1 \CACHE_MEM_reg[6][65]  ( .D(n11689), .CK(N28803), .QN(n9043) );
  DFF_X1 \CACHE_MEM_reg[6][64]  ( .D(n11688), .CK(N28803), .QN(n9059) );
  DFF_X1 \CACHE_MEM_reg[6][63]  ( .D(n11687), .CK(N28803), .QN(n9075) );
  DFF_X1 \CACHE_MEM_reg[6][62]  ( .D(n11686), .CK(N28803), .QN(n9091) );
  DFF_X1 \CACHE_MEM_reg[6][61]  ( .D(n11685), .CK(N28803), .QN(n9107) );
  DFF_X1 \CACHE_MEM_reg[6][60]  ( .D(n11684), .CK(N28803), .QN(n9123) );
  DFF_X1 \CACHE_MEM_reg[6][59]  ( .D(n11683), .CK(N28803), .QN(n9139) );
  DFF_X1 \CACHE_MEM_reg[6][58]  ( .D(n11682), .CK(N28803), .QN(n9155) );
  DFF_X1 \CACHE_MEM_reg[6][57]  ( .D(n11681), .CK(N28803), .QN(n9171) );
  DFF_X1 \CACHE_MEM_reg[6][56]  ( .D(n11680), .CK(N28803), .QN(n9187) );
  DFF_X1 \CACHE_MEM_reg[6][55]  ( .D(n11679), .CK(N28803), .QN(n9203) );
  DFF_X1 \CACHE_MEM_reg[6][54]  ( .D(n11678), .CK(N28803), .QN(n9219) );
  DFF_X1 \CACHE_MEM_reg[6][53]  ( .D(n11677), .CK(N28803), .QN(n9235) );
  DFF_X1 \CACHE_MEM_reg[6][52]  ( .D(n11676), .CK(N28803), .QN(n9251) );
  DFF_X1 \CACHE_MEM_reg[6][51]  ( .D(n11675), .CK(N28803), .QN(n9267) );
  DFF_X1 \CACHE_MEM_reg[6][50]  ( .D(n11674), .CK(N28803), .QN(n9283) );
  DFF_X1 \CACHE_MEM_reg[6][49]  ( .D(n11673), .CK(N28803), .QN(n9299) );
  DFF_X1 \CACHE_MEM_reg[6][48]  ( .D(n11672), .CK(N28803), .QN(n9315) );
  DFF_X1 \CACHE_MEM_reg[6][47]  ( .D(n11671), .CK(N28803), .QN(n9331) );
  DFF_X1 \CACHE_MEM_reg[6][46]  ( .D(n11670), .CK(N28803), .QN(n9347) );
  DFF_X1 \CACHE_MEM_reg[6][45]  ( .D(n11669), .CK(N28803), .QN(n9363) );
  DFF_X1 \CACHE_MEM_reg[6][44]  ( .D(n11668), .CK(N28803), .QN(n9379) );
  DFF_X1 \CACHE_MEM_reg[6][43]  ( .D(n11667), .CK(N28803), .QN(n9395) );
  DFF_X1 \CACHE_MEM_reg[6][42]  ( .D(n11666), .CK(N28803), .QN(n9411) );
  DFF_X1 \CACHE_MEM_reg[6][41]  ( .D(n11665), .CK(N28803), .QN(n9427) );
  DFF_X1 \CACHE_MEM_reg[6][40]  ( .D(n11664), .CK(N28803), .QN(n9443) );
  DFF_X1 \CACHE_MEM_reg[6][39]  ( .D(n11663), .CK(N28803), .QN(n9459) );
  DFF_X1 \CACHE_MEM_reg[6][38]  ( .D(n11662), .CK(N28803), .QN(n9475) );
  DFF_X1 \CACHE_MEM_reg[6][37]  ( .D(n11661), .CK(N28803), .QN(n9491) );
  DFF_X1 \CACHE_MEM_reg[6][36]  ( .D(n11660), .CK(N28803), .QN(n9507) );
  DFF_X1 \CACHE_MEM_reg[6][35]  ( .D(n11659), .CK(N28803), .QN(n9523) );
  DFF_X1 \CACHE_MEM_reg[6][34]  ( .D(n11658), .CK(N28803), .QN(n9539) );
  DFF_X1 \CACHE_MEM_reg[6][33]  ( .D(n11657), .CK(N28803), .QN(n9555) );
  DFF_X1 \CACHE_MEM_reg[6][32]  ( .D(n11656), .CK(N28803), .QN(n9571) );
  DFF_X1 \CACHE_MEM_reg[6][31]  ( .D(n11655), .CK(N28803), .QN(n9587) );
  DFF_X1 \CACHE_MEM_reg[6][30]  ( .D(n11654), .CK(N28803), .QN(n9603) );
  DFF_X1 \CACHE_MEM_reg[6][29]  ( .D(n11653), .CK(N28803), .QN(n9619) );
  DFF_X1 \CACHE_MEM_reg[6][28]  ( .D(n11652), .CK(N28803), .QN(n9635) );
  DFF_X1 \CACHE_MEM_reg[6][27]  ( .D(n11651), .CK(N28803), .QN(n9651) );
  DFF_X1 \CACHE_MEM_reg[6][26]  ( .D(n11650), .CK(N28803), .QN(n9667) );
  DFF_X1 \CACHE_MEM_reg[6][25]  ( .D(n11649), .CK(N28803), .QN(n9683) );
  DFF_X1 \CACHE_MEM_reg[6][24]  ( .D(n11648), .CK(N28803), .QN(n9699) );
  DFF_X1 \CACHE_MEM_reg[6][23]  ( .D(n11647), .CK(N28803), .QN(n9715) );
  DFF_X1 \CACHE_MEM_reg[6][22]  ( .D(n11646), .CK(N28803), .QN(n9731) );
  DFF_X1 \CACHE_MEM_reg[6][21]  ( .D(n11645), .CK(N28803), .QN(n9747) );
  DFF_X1 \CACHE_MEM_reg[6][20]  ( .D(n11644), .CK(N28803), .QN(n9763) );
  DFF_X1 \CACHE_MEM_reg[6][19]  ( .D(n11643), .CK(N28803), .QN(n9779) );
  DFF_X1 \CACHE_MEM_reg[6][18]  ( .D(n11642), .CK(N28803), .QN(n9795) );
  DFF_X1 \CACHE_MEM_reg[6][17]  ( .D(n11641), .CK(N28803), .QN(n9811) );
  DFF_X1 \CACHE_MEM_reg[6][16]  ( .D(n11640), .CK(N28803), .QN(n9827) );
  DFF_X1 \CACHE_MEM_reg[6][15]  ( .D(n11639), .CK(N28803), .QN(n9843) );
  DFF_X1 \CACHE_MEM_reg[6][14]  ( .D(n11638), .CK(N28803), .QN(n9859) );
  DFF_X1 \CACHE_MEM_reg[6][13]  ( .D(n11637), .CK(N28803), .QN(n9875) );
  DFF_X1 \CACHE_MEM_reg[6][12]  ( .D(n11636), .CK(N28803), .QN(n9891) );
  DFF_X1 \CACHE_MEM_reg[6][11]  ( .D(n11635), .CK(N28803), .QN(n9907) );
  DFF_X1 \CACHE_MEM_reg[6][10]  ( .D(n11634), .CK(N28803), .QN(n9923) );
  DFF_X1 \CACHE_MEM_reg[6][9]  ( .D(n11633), .CK(N28803), .QN(n9939) );
  DFF_X1 \CACHE_MEM_reg[6][8]  ( .D(n11632), .CK(N28803), .QN(n9955) );
  DFF_X1 \CACHE_MEM_reg[6][7]  ( .D(n11631), .CK(N28803), .QN(n9971) );
  DFF_X1 \CACHE_MEM_reg[6][6]  ( .D(n11630), .CK(N28803), .QN(n9987) );
  DFF_X1 \CACHE_MEM_reg[6][5]  ( .D(n11629), .CK(N28803), .QN(n10003) );
  DFF_X1 \CACHE_MEM_reg[6][4]  ( .D(n11628), .CK(N28803), .QN(n10019) );
  DFF_X1 \CACHE_MEM_reg[6][3]  ( .D(n11627), .CK(N28803), .QN(n10035) );
  DFF_X1 \CACHE_MEM_reg[6][2]  ( .D(n11626), .CK(N28803), .QN(n10051) );
  DFF_X1 \CACHE_MEM_reg[6][1]  ( .D(n11625), .CK(N28803), .QN(n10067) );
  DFF_X1 \CACHE_MEM_reg[6][0]  ( .D(n11624), .CK(N28803), .QN(n10083) );
  DFF_X1 \CACHE_MEM_reg[5][255]  ( .D(n11623), .CK(N28803), .QN(n5999) );
  DFF_X1 \CACHE_MEM_reg[5][254]  ( .D(n11622), .CK(N28803), .QN(n6015) );
  DFF_X1 \CACHE_MEM_reg[5][253]  ( .D(n11621), .CK(N28803), .QN(n6031) );
  DFF_X1 \CACHE_MEM_reg[5][252]  ( .D(n11620), .CK(N28803), .QN(n6047) );
  DFF_X1 \CACHE_MEM_reg[5][251]  ( .D(n11619), .CK(N28803), .QN(n6063) );
  DFF_X1 \CACHE_MEM_reg[5][250]  ( .D(n11618), .CK(N28803), .QN(n6079) );
  DFF_X1 \CACHE_MEM_reg[5][249]  ( .D(n11617), .CK(N28803), .QN(n6095) );
  DFF_X1 \CACHE_MEM_reg[5][248]  ( .D(n11616), .CK(N28803), .QN(n6111) );
  DFF_X1 \CACHE_MEM_reg[5][247]  ( .D(n11615), .CK(N28803), .QN(n6127) );
  DFF_X1 \CACHE_MEM_reg[5][246]  ( .D(n11614), .CK(N28803), .QN(n6143) );
  DFF_X1 \CACHE_MEM_reg[5][245]  ( .D(n11613), .CK(N28803), .QN(n6159) );
  DFF_X1 \CACHE_MEM_reg[5][244]  ( .D(n11612), .CK(N28803), .QN(n6175) );
  DFF_X1 \CACHE_MEM_reg[5][243]  ( .D(n11611), .CK(N28803), .QN(n6191) );
  DFF_X1 \CACHE_MEM_reg[5][242]  ( .D(n11610), .CK(N28803), .QN(n6207) );
  DFF_X1 \CACHE_MEM_reg[5][241]  ( .D(n11609), .CK(N28803), .QN(n6223) );
  DFF_X1 \CACHE_MEM_reg[5][240]  ( .D(n11608), .CK(N28803), .QN(n6239) );
  DFF_X1 \CACHE_MEM_reg[5][239]  ( .D(n11607), .CK(N28803), .QN(n6255) );
  DFF_X1 \CACHE_MEM_reg[5][238]  ( .D(n11606), .CK(N28803), .QN(n6271) );
  DFF_X1 \CACHE_MEM_reg[5][237]  ( .D(n11605), .CK(N28803), .QN(n6287) );
  DFF_X1 \CACHE_MEM_reg[5][236]  ( .D(n11604), .CK(N28803), .QN(n6303) );
  DFF_X1 \CACHE_MEM_reg[5][235]  ( .D(n11603), .CK(N28803), .QN(n6319) );
  DFF_X1 \CACHE_MEM_reg[5][234]  ( .D(n11602), .CK(N28803), .QN(n6335) );
  DFF_X1 \CACHE_MEM_reg[5][233]  ( .D(n11601), .CK(N28803), .QN(n6351) );
  DFF_X1 \CACHE_MEM_reg[5][232]  ( .D(n11600), .CK(N28803), .QN(n6367) );
  DFF_X1 \CACHE_MEM_reg[5][231]  ( .D(n11599), .CK(N28803), .QN(n6383) );
  DFF_X1 \CACHE_MEM_reg[5][230]  ( .D(n11598), .CK(N28803), .QN(n6399) );
  DFF_X1 \CACHE_MEM_reg[5][229]  ( .D(n11597), .CK(N28803), .QN(n6415) );
  DFF_X1 \CACHE_MEM_reg[5][228]  ( .D(n11596), .CK(N28803), .QN(n6431) );
  DFF_X1 \CACHE_MEM_reg[5][227]  ( .D(n11595), .CK(N28803), .QN(n6447) );
  DFF_X1 \CACHE_MEM_reg[5][226]  ( .D(n11594), .CK(N28803), .QN(n6463) );
  DFF_X1 \CACHE_MEM_reg[5][225]  ( .D(n11593), .CK(N28803), .QN(n6479) );
  DFF_X1 \CACHE_MEM_reg[5][224]  ( .D(n11592), .CK(N28803), .QN(n6495) );
  DFF_X1 \CACHE_MEM_reg[5][223]  ( .D(n11591), .CK(N28803), .QN(n6511) );
  DFF_X1 \CACHE_MEM_reg[5][222]  ( .D(n11590), .CK(N28803), .QN(n6527) );
  DFF_X1 \CACHE_MEM_reg[5][221]  ( .D(n11589), .CK(N28803), .QN(n6543) );
  DFF_X1 \CACHE_MEM_reg[5][220]  ( .D(n11588), .CK(N28803), .QN(n6559) );
  DFF_X1 \CACHE_MEM_reg[5][219]  ( .D(n11587), .CK(N28803), .QN(n6575) );
  DFF_X1 \CACHE_MEM_reg[5][218]  ( .D(n11586), .CK(N28803), .QN(n6591) );
  DFF_X1 \CACHE_MEM_reg[5][217]  ( .D(n11585), .CK(N28803), .QN(n6607) );
  DFF_X1 \CACHE_MEM_reg[5][216]  ( .D(n11584), .CK(N28803), .QN(n6623) );
  DFF_X1 \CACHE_MEM_reg[5][215]  ( .D(n11583), .CK(N28803), .QN(n6639) );
  DFF_X1 \CACHE_MEM_reg[5][214]  ( .D(n11582), .CK(N28803), .QN(n6655) );
  DFF_X1 \CACHE_MEM_reg[5][213]  ( .D(n11581), .CK(N28803), .QN(n6671) );
  DFF_X1 \CACHE_MEM_reg[5][212]  ( .D(n11580), .CK(N28803), .QN(n6687) );
  DFF_X1 \CACHE_MEM_reg[5][211]  ( .D(n11579), .CK(N28803), .QN(n6703) );
  DFF_X1 \CACHE_MEM_reg[5][210]  ( .D(n11578), .CK(N28803), .QN(n6719) );
  DFF_X1 \CACHE_MEM_reg[5][209]  ( .D(n11577), .CK(N28803), .QN(n6735) );
  DFF_X1 \CACHE_MEM_reg[5][208]  ( .D(n11576), .CK(N28803), .QN(n6751) );
  DFF_X1 \CACHE_MEM_reg[5][207]  ( .D(n11575), .CK(N28803), .QN(n6767) );
  DFF_X1 \CACHE_MEM_reg[5][206]  ( .D(n11574), .CK(N28803), .QN(n6783) );
  DFF_X1 \CACHE_MEM_reg[5][205]  ( .D(n11573), .CK(N28803), .QN(n6799) );
  DFF_X1 \CACHE_MEM_reg[5][204]  ( .D(n11572), .CK(N28803), .QN(n6815) );
  DFF_X1 \CACHE_MEM_reg[5][203]  ( .D(n11571), .CK(N28803), .QN(n6831) );
  DFF_X1 \CACHE_MEM_reg[5][202]  ( .D(n11570), .CK(N28803), .QN(n6847) );
  DFF_X1 \CACHE_MEM_reg[5][201]  ( .D(n11569), .CK(N28803), .QN(n6863) );
  DFF_X1 \CACHE_MEM_reg[5][200]  ( .D(n11568), .CK(N28803), .QN(n6879) );
  DFF_X1 \CACHE_MEM_reg[5][199]  ( .D(n11567), .CK(N28803), .QN(n6895) );
  DFF_X1 \CACHE_MEM_reg[5][198]  ( .D(n11566), .CK(N28803), .QN(n6911) );
  DFF_X1 \CACHE_MEM_reg[5][197]  ( .D(n11565), .CK(N28803), .QN(n6927) );
  DFF_X1 \CACHE_MEM_reg[5][196]  ( .D(n11564), .CK(N28803), .QN(n6943) );
  DFF_X1 \CACHE_MEM_reg[5][195]  ( .D(n11563), .CK(N28803), .QN(n6959) );
  DFF_X1 \CACHE_MEM_reg[5][194]  ( .D(n11562), .CK(N28803), .QN(n6975) );
  DFF_X1 \CACHE_MEM_reg[5][193]  ( .D(n11561), .CK(N28803), .QN(n6991) );
  DFF_X1 \CACHE_MEM_reg[5][192]  ( .D(n11560), .CK(N28803), .QN(n7007) );
  DFF_X1 \CACHE_MEM_reg[5][191]  ( .D(n11559), .CK(N28803), .QN(n7023) );
  DFF_X1 \CACHE_MEM_reg[5][190]  ( .D(n11558), .CK(N28803), .QN(n7039) );
  DFF_X1 \CACHE_MEM_reg[5][189]  ( .D(n11557), .CK(N28803), .QN(n7055) );
  DFF_X1 \CACHE_MEM_reg[5][188]  ( .D(n11556), .CK(N28803), .QN(n7071) );
  DFF_X1 \CACHE_MEM_reg[5][187]  ( .D(n11555), .CK(N28803), .QN(n7087) );
  DFF_X1 \CACHE_MEM_reg[5][186]  ( .D(n11554), .CK(N28803), .QN(n7103) );
  DFF_X1 \CACHE_MEM_reg[5][185]  ( .D(n11553), .CK(N28803), .QN(n7119) );
  DFF_X1 \CACHE_MEM_reg[5][184]  ( .D(n11552), .CK(N28803), .QN(n7135) );
  DFF_X1 \CACHE_MEM_reg[5][183]  ( .D(n11551), .CK(N28803), .QN(n7151) );
  DFF_X1 \CACHE_MEM_reg[5][182]  ( .D(n11550), .CK(N28803), .QN(n7167) );
  DFF_X1 \CACHE_MEM_reg[5][181]  ( .D(n11549), .CK(N28803), .QN(n7183) );
  DFF_X1 \CACHE_MEM_reg[5][180]  ( .D(n11548), .CK(N28803), .QN(n7199) );
  DFF_X1 \CACHE_MEM_reg[5][179]  ( .D(n11547), .CK(N28803), .QN(n7215) );
  DFF_X1 \CACHE_MEM_reg[5][178]  ( .D(n11546), .CK(N28803), .QN(n7231) );
  DFF_X1 \CACHE_MEM_reg[5][177]  ( .D(n11545), .CK(N28803), .QN(n7247) );
  DFF_X1 \CACHE_MEM_reg[5][176]  ( .D(n11544), .CK(N28803), .QN(n7263) );
  DFF_X1 \CACHE_MEM_reg[5][175]  ( .D(n11543), .CK(N28803), .QN(n7279) );
  DFF_X1 \CACHE_MEM_reg[5][174]  ( .D(n11542), .CK(N28803), .QN(n7295) );
  DFF_X1 \CACHE_MEM_reg[5][173]  ( .D(n11541), .CK(N28803), .QN(n7311) );
  DFF_X1 \CACHE_MEM_reg[5][172]  ( .D(n11540), .CK(N28803), .QN(n7327) );
  DFF_X1 \CACHE_MEM_reg[5][171]  ( .D(n11539), .CK(N28803), .QN(n7343) );
  DFF_X1 \CACHE_MEM_reg[5][170]  ( .D(n11538), .CK(N28803), .QN(n7359) );
  DFF_X1 \CACHE_MEM_reg[5][169]  ( .D(n11537), .CK(N28803), .QN(n7375) );
  DFF_X1 \CACHE_MEM_reg[5][168]  ( .D(n11536), .CK(N28803), .QN(n7391) );
  DFF_X1 \CACHE_MEM_reg[5][167]  ( .D(n11535), .CK(N28803), .QN(n7407) );
  DFF_X1 \CACHE_MEM_reg[5][166]  ( .D(n11534), .CK(N28803), .QN(n7423) );
  DFF_X1 \CACHE_MEM_reg[5][165]  ( .D(n11533), .CK(N28803), .QN(n7439) );
  DFF_X1 \CACHE_MEM_reg[5][164]  ( .D(n11532), .CK(N28803), .QN(n7455) );
  DFF_X1 \CACHE_MEM_reg[5][163]  ( .D(n11531), .CK(N28803), .QN(n7471) );
  DFF_X1 \CACHE_MEM_reg[5][162]  ( .D(n11530), .CK(N28803), .QN(n7487) );
  DFF_X1 \CACHE_MEM_reg[5][161]  ( .D(n11529), .CK(N28803), .QN(n7503) );
  DFF_X1 \CACHE_MEM_reg[5][160]  ( .D(n11528), .CK(N28803), .QN(n7519) );
  DFF_X1 \CACHE_MEM_reg[5][159]  ( .D(n11527), .CK(N28803), .QN(n7535) );
  DFF_X1 \CACHE_MEM_reg[5][158]  ( .D(n11526), .CK(N28803), .QN(n7551) );
  DFF_X1 \CACHE_MEM_reg[5][157]  ( .D(n11525), .CK(N28803), .QN(n7567) );
  DFF_X1 \CACHE_MEM_reg[5][156]  ( .D(n11524), .CK(N28803), .QN(n7583) );
  DFF_X1 \CACHE_MEM_reg[5][155]  ( .D(n11523), .CK(N28803), .QN(n7599) );
  DFF_X1 \CACHE_MEM_reg[5][154]  ( .D(n11522), .CK(N28803), .QN(n7615) );
  DFF_X1 \CACHE_MEM_reg[5][153]  ( .D(n11521), .CK(N28803), .QN(n7631) );
  DFF_X1 \CACHE_MEM_reg[5][152]  ( .D(n11520), .CK(N28803), .QN(n7647) );
  DFF_X1 \CACHE_MEM_reg[5][151]  ( .D(n11519), .CK(N28803), .QN(n7663) );
  DFF_X1 \CACHE_MEM_reg[5][150]  ( .D(n11518), .CK(N28803), .QN(n7679) );
  DFF_X1 \CACHE_MEM_reg[5][149]  ( .D(n11517), .CK(N28803), .QN(n7695) );
  DFF_X1 \CACHE_MEM_reg[5][148]  ( .D(n11516), .CK(N28803), .QN(n7711) );
  DFF_X1 \CACHE_MEM_reg[5][147]  ( .D(n11515), .CK(N28803), .QN(n7727) );
  DFF_X1 \CACHE_MEM_reg[5][146]  ( .D(n11514), .CK(N28803), .QN(n7743) );
  DFF_X1 \CACHE_MEM_reg[5][145]  ( .D(n11513), .CK(N28803), .QN(n7759) );
  DFF_X1 \CACHE_MEM_reg[5][144]  ( .D(n11512), .CK(N28803), .QN(n7775) );
  DFF_X1 \CACHE_MEM_reg[5][143]  ( .D(n11511), .CK(N28803), .QN(n7791) );
  DFF_X1 \CACHE_MEM_reg[5][142]  ( .D(n11510), .CK(N28803), .QN(n7807) );
  DFF_X1 \CACHE_MEM_reg[5][141]  ( .D(n11509), .CK(N28803), .QN(n7823) );
  DFF_X1 \CACHE_MEM_reg[5][140]  ( .D(n11508), .CK(N28803), .QN(n7839) );
  DFF_X1 \CACHE_MEM_reg[5][139]  ( .D(n11507), .CK(N28803), .QN(n7855) );
  DFF_X1 \CACHE_MEM_reg[5][138]  ( .D(n11506), .CK(N28803), .QN(n7871) );
  DFF_X1 \CACHE_MEM_reg[5][137]  ( .D(n11505), .CK(N28803), .QN(n7887) );
  DFF_X1 \CACHE_MEM_reg[5][136]  ( .D(n11504), .CK(N28803), .QN(n7903) );
  DFF_X1 \CACHE_MEM_reg[5][135]  ( .D(n11503), .CK(N28803), .QN(n7919) );
  DFF_X1 \CACHE_MEM_reg[5][134]  ( .D(n11502), .CK(N28803), .QN(n7935) );
  DFF_X1 \CACHE_MEM_reg[5][133]  ( .D(n11501), .CK(N28803), .QN(n7951) );
  DFF_X1 \CACHE_MEM_reg[5][132]  ( .D(n11500), .CK(N28803), .QN(n7967) );
  DFF_X1 \CACHE_MEM_reg[5][131]  ( .D(n11499), .CK(N28803), .QN(n7983) );
  DFF_X1 \CACHE_MEM_reg[5][130]  ( .D(n11498), .CK(N28803), .QN(n7999) );
  DFF_X1 \CACHE_MEM_reg[5][129]  ( .D(n11497), .CK(N28803), .QN(n8015) );
  DFF_X1 \CACHE_MEM_reg[5][128]  ( .D(n11496), .CK(N28803), .QN(n8031) );
  DFF_X1 \CACHE_MEM_reg[5][127]  ( .D(n11495), .CK(N28803), .QN(n8047) );
  DFF_X1 \CACHE_MEM_reg[5][126]  ( .D(n11494), .CK(N28803), .QN(n8063) );
  DFF_X1 \CACHE_MEM_reg[5][125]  ( .D(n11493), .CK(N28803), .QN(n8079) );
  DFF_X1 \CACHE_MEM_reg[5][124]  ( .D(n11492), .CK(N28803), .QN(n8095) );
  DFF_X1 \CACHE_MEM_reg[5][123]  ( .D(n11491), .CK(N28803), .QN(n8111) );
  DFF_X1 \CACHE_MEM_reg[5][122]  ( .D(n11490), .CK(N28803), .QN(n8127) );
  DFF_X1 \CACHE_MEM_reg[5][121]  ( .D(n11489), .CK(N28803), .QN(n8143) );
  DFF_X1 \CACHE_MEM_reg[5][120]  ( .D(n11488), .CK(N28803), .QN(n8159) );
  DFF_X1 \CACHE_MEM_reg[5][119]  ( .D(n11487), .CK(N28803), .QN(n8175) );
  DFF_X1 \CACHE_MEM_reg[5][118]  ( .D(n11486), .CK(N28803), .QN(n8191) );
  DFF_X1 \CACHE_MEM_reg[5][117]  ( .D(n11485), .CK(N28803), .QN(n8207) );
  DFF_X1 \CACHE_MEM_reg[5][116]  ( .D(n11484), .CK(N28803), .QN(n8223) );
  DFF_X1 \CACHE_MEM_reg[5][115]  ( .D(n11483), .CK(N28803), .QN(n8239) );
  DFF_X1 \CACHE_MEM_reg[5][114]  ( .D(n11482), .CK(N28803), .QN(n8255) );
  DFF_X1 \CACHE_MEM_reg[5][113]  ( .D(n11481), .CK(N28803), .QN(n8271) );
  DFF_X1 \CACHE_MEM_reg[5][112]  ( .D(n11480), .CK(N28803), .QN(n8287) );
  DFF_X1 \CACHE_MEM_reg[5][111]  ( .D(n11479), .CK(N28803), .QN(n8303) );
  DFF_X1 \CACHE_MEM_reg[5][110]  ( .D(n11478), .CK(N28803), .QN(n8319) );
  DFF_X1 \CACHE_MEM_reg[5][109]  ( .D(n11477), .CK(N28803), .QN(n8335) );
  DFF_X1 \CACHE_MEM_reg[5][108]  ( .D(n11476), .CK(N28803), .QN(n8351) );
  DFF_X1 \CACHE_MEM_reg[5][107]  ( .D(n11475), .CK(N28803), .QN(n8367) );
  DFF_X1 \CACHE_MEM_reg[5][106]  ( .D(n11474), .CK(N28803), .QN(n8383) );
  DFF_X1 \CACHE_MEM_reg[5][105]  ( .D(n11473), .CK(N28803), .QN(n8399) );
  DFF_X1 \CACHE_MEM_reg[5][104]  ( .D(n11472), .CK(N28803), .QN(n8415) );
  DFF_X1 \CACHE_MEM_reg[5][103]  ( .D(n11471), .CK(N28803), .QN(n8431) );
  DFF_X1 \CACHE_MEM_reg[5][102]  ( .D(n11470), .CK(N28803), .QN(n8447) );
  DFF_X1 \CACHE_MEM_reg[5][101]  ( .D(n11469), .CK(N28803), .QN(n8463) );
  DFF_X1 \CACHE_MEM_reg[5][100]  ( .D(n11468), .CK(N28803), .QN(n8479) );
  DFF_X1 \CACHE_MEM_reg[5][99]  ( .D(n11467), .CK(N28803), .QN(n8495) );
  DFF_X1 \CACHE_MEM_reg[5][98]  ( .D(n11466), .CK(N28803), .QN(n8511) );
  DFF_X1 \CACHE_MEM_reg[5][97]  ( .D(n11465), .CK(N28803), .QN(n8527) );
  DFF_X1 \CACHE_MEM_reg[5][96]  ( .D(n11464), .CK(N28803), .QN(n8543) );
  DFF_X1 \CACHE_MEM_reg[5][95]  ( .D(n11463), .CK(N28803), .QN(n8559) );
  DFF_X1 \CACHE_MEM_reg[5][94]  ( .D(n11462), .CK(N28803), .QN(n8575) );
  DFF_X1 \CACHE_MEM_reg[5][93]  ( .D(n11461), .CK(N28803), .QN(n8591) );
  DFF_X1 \CACHE_MEM_reg[5][92]  ( .D(n11460), .CK(N28803), .QN(n8607) );
  DFF_X1 \CACHE_MEM_reg[5][91]  ( .D(n11459), .CK(N28803), .QN(n8623) );
  DFF_X1 \CACHE_MEM_reg[5][90]  ( .D(n11458), .CK(N28803), .QN(n8639) );
  DFF_X1 \CACHE_MEM_reg[5][89]  ( .D(n11457), .CK(N28803), .QN(n8655) );
  DFF_X1 \CACHE_MEM_reg[5][88]  ( .D(n11456), .CK(N28803), .QN(n8671) );
  DFF_X1 \CACHE_MEM_reg[5][87]  ( .D(n11455), .CK(N28803), .QN(n8687) );
  DFF_X1 \CACHE_MEM_reg[5][86]  ( .D(n11454), .CK(N28803), .QN(n8703) );
  DFF_X1 \CACHE_MEM_reg[5][85]  ( .D(n11453), .CK(N28803), .QN(n8719) );
  DFF_X1 \CACHE_MEM_reg[5][84]  ( .D(n11452), .CK(N28803), .QN(n8735) );
  DFF_X1 \CACHE_MEM_reg[5][83]  ( .D(n11451), .CK(N28803), .QN(n8751) );
  DFF_X1 \CACHE_MEM_reg[5][82]  ( .D(n11450), .CK(N28803), .QN(n8767) );
  DFF_X1 \CACHE_MEM_reg[5][81]  ( .D(n11449), .CK(N28803), .QN(n8783) );
  DFF_X1 \CACHE_MEM_reg[5][80]  ( .D(n11448), .CK(N28803), .QN(n8799) );
  DFF_X1 \CACHE_MEM_reg[5][79]  ( .D(n11447), .CK(N28803), .QN(n8815) );
  DFF_X1 \CACHE_MEM_reg[5][78]  ( .D(n11446), .CK(N28803), .QN(n8831) );
  DFF_X1 \CACHE_MEM_reg[5][77]  ( .D(n11445), .CK(N28803), .QN(n8847) );
  DFF_X1 \CACHE_MEM_reg[5][76]  ( .D(n11444), .CK(N28803), .QN(n8863) );
  DFF_X1 \CACHE_MEM_reg[5][75]  ( .D(n11443), .CK(N28803), .QN(n8879) );
  DFF_X1 \CACHE_MEM_reg[5][74]  ( .D(n11442), .CK(N28803), .QN(n8895) );
  DFF_X1 \CACHE_MEM_reg[5][73]  ( .D(n11441), .CK(N28803), .QN(n8911) );
  DFF_X1 \CACHE_MEM_reg[5][72]  ( .D(n11440), .CK(N28803), .QN(n8927) );
  DFF_X1 \CACHE_MEM_reg[5][71]  ( .D(n11439), .CK(N28803), .QN(n8943) );
  DFF_X1 \CACHE_MEM_reg[5][70]  ( .D(n11438), .CK(N28803), .QN(n8959) );
  DFF_X1 \CACHE_MEM_reg[5][69]  ( .D(n11437), .CK(N28803), .QN(n8975) );
  DFF_X1 \CACHE_MEM_reg[5][68]  ( .D(n11436), .CK(N28803), .QN(n8991) );
  DFF_X1 \CACHE_MEM_reg[5][67]  ( .D(n11435), .CK(N28803), .QN(n9007) );
  DFF_X1 \CACHE_MEM_reg[5][66]  ( .D(n11434), .CK(N28803), .QN(n9023) );
  DFF_X1 \CACHE_MEM_reg[5][65]  ( .D(n11433), .CK(N28803), .QN(n9039) );
  DFF_X1 \CACHE_MEM_reg[5][64]  ( .D(n11432), .CK(N28803), .QN(n9055) );
  DFF_X1 \CACHE_MEM_reg[5][63]  ( .D(n11431), .CK(N28803), .QN(n9071) );
  DFF_X1 \CACHE_MEM_reg[5][62]  ( .D(n11430), .CK(N28803), .QN(n9087) );
  DFF_X1 \CACHE_MEM_reg[5][61]  ( .D(n11429), .CK(N28803), .QN(n9103) );
  DFF_X1 \CACHE_MEM_reg[5][60]  ( .D(n11428), .CK(N28803), .QN(n9119) );
  DFF_X1 \CACHE_MEM_reg[5][59]  ( .D(n11427), .CK(N28803), .QN(n9135) );
  DFF_X1 \CACHE_MEM_reg[5][58]  ( .D(n11426), .CK(N28803), .QN(n9151) );
  DFF_X1 \CACHE_MEM_reg[5][57]  ( .D(n11425), .CK(N28803), .QN(n9167) );
  DFF_X1 \CACHE_MEM_reg[5][56]  ( .D(n11424), .CK(N28803), .QN(n9183) );
  DFF_X1 \CACHE_MEM_reg[5][55]  ( .D(n11423), .CK(N28803), .QN(n9199) );
  DFF_X1 \CACHE_MEM_reg[5][54]  ( .D(n11422), .CK(N28803), .QN(n9215) );
  DFF_X1 \CACHE_MEM_reg[5][53]  ( .D(n11421), .CK(N28803), .QN(n9231) );
  DFF_X1 \CACHE_MEM_reg[5][52]  ( .D(n11420), .CK(N28803), .QN(n9247) );
  DFF_X1 \CACHE_MEM_reg[5][51]  ( .D(n11419), .CK(N28803), .QN(n9263) );
  DFF_X1 \CACHE_MEM_reg[5][50]  ( .D(n11418), .CK(N28803), .QN(n9279) );
  DFF_X1 \CACHE_MEM_reg[5][49]  ( .D(n11417), .CK(N28803), .QN(n9295) );
  DFF_X1 \CACHE_MEM_reg[5][48]  ( .D(n11416), .CK(N28803), .QN(n9311) );
  DFF_X1 \CACHE_MEM_reg[5][47]  ( .D(n11415), .CK(N28803), .QN(n9327) );
  DFF_X1 \CACHE_MEM_reg[5][46]  ( .D(n11414), .CK(N28803), .QN(n9343) );
  DFF_X1 \CACHE_MEM_reg[5][45]  ( .D(n11413), .CK(N28803), .QN(n9359) );
  DFF_X1 \CACHE_MEM_reg[5][44]  ( .D(n11412), .CK(N28803), .QN(n9375) );
  DFF_X1 \CACHE_MEM_reg[5][43]  ( .D(n11411), .CK(N28803), .QN(n9391) );
  DFF_X1 \CACHE_MEM_reg[5][42]  ( .D(n11410), .CK(N28803), .QN(n9407) );
  DFF_X1 \CACHE_MEM_reg[5][41]  ( .D(n11409), .CK(N28803), .QN(n9423) );
  DFF_X1 \CACHE_MEM_reg[5][40]  ( .D(n11408), .CK(N28803), .QN(n9439) );
  DFF_X1 \CACHE_MEM_reg[5][39]  ( .D(n11407), .CK(N28803), .QN(n9455) );
  DFF_X1 \CACHE_MEM_reg[5][38]  ( .D(n11406), .CK(N28803), .QN(n9471) );
  DFF_X1 \CACHE_MEM_reg[5][37]  ( .D(n11405), .CK(N28803), .QN(n9487) );
  DFF_X1 \CACHE_MEM_reg[5][36]  ( .D(n11404), .CK(N28803), .QN(n9503) );
  DFF_X1 \CACHE_MEM_reg[5][35]  ( .D(n11403), .CK(N28803), .QN(n9519) );
  DFF_X1 \CACHE_MEM_reg[5][34]  ( .D(n11402), .CK(N28803), .QN(n9535) );
  DFF_X1 \CACHE_MEM_reg[5][33]  ( .D(n11401), .CK(N28803), .QN(n9551) );
  DFF_X1 \CACHE_MEM_reg[5][32]  ( .D(n11400), .CK(N28803), .QN(n9567) );
  DFF_X1 \CACHE_MEM_reg[5][31]  ( .D(n11399), .CK(N28803), .QN(n9583) );
  DFF_X1 \CACHE_MEM_reg[5][30]  ( .D(n11398), .CK(N28803), .QN(n9599) );
  DFF_X1 \CACHE_MEM_reg[5][29]  ( .D(n11397), .CK(N28803), .QN(n9615) );
  DFF_X1 \CACHE_MEM_reg[5][28]  ( .D(n11396), .CK(N28803), .QN(n9631) );
  DFF_X1 \CACHE_MEM_reg[5][27]  ( .D(n11395), .CK(N28803), .QN(n9647) );
  DFF_X1 \CACHE_MEM_reg[5][26]  ( .D(n11394), .CK(N28803), .QN(n9663) );
  DFF_X1 \CACHE_MEM_reg[5][25]  ( .D(n11393), .CK(N28803), .QN(n9679) );
  DFF_X1 \CACHE_MEM_reg[5][24]  ( .D(n11392), .CK(N28803), .QN(n9695) );
  DFF_X1 \CACHE_MEM_reg[5][23]  ( .D(n11391), .CK(N28803), .QN(n9711) );
  DFF_X1 \CACHE_MEM_reg[5][22]  ( .D(n11390), .CK(N28803), .QN(n9727) );
  DFF_X1 \CACHE_MEM_reg[5][21]  ( .D(n11389), .CK(N28803), .QN(n9743) );
  DFF_X1 \CACHE_MEM_reg[5][20]  ( .D(n11388), .CK(N28803), .QN(n9759) );
  DFF_X1 \CACHE_MEM_reg[5][19]  ( .D(n11387), .CK(N28803), .QN(n9775) );
  DFF_X1 \CACHE_MEM_reg[5][18]  ( .D(n11386), .CK(N28803), .QN(n9791) );
  DFF_X1 \CACHE_MEM_reg[5][17]  ( .D(n11385), .CK(N28803), .QN(n9807) );
  DFF_X1 \CACHE_MEM_reg[5][16]  ( .D(n11384), .CK(N28803), .QN(n9823) );
  DFF_X1 \CACHE_MEM_reg[5][15]  ( .D(n11383), .CK(N28803), .QN(n9839) );
  DFF_X1 \CACHE_MEM_reg[5][14]  ( .D(n11382), .CK(N28803), .QN(n9855) );
  DFF_X1 \CACHE_MEM_reg[5][13]  ( .D(n11381), .CK(N28803), .QN(n9871) );
  DFF_X1 \CACHE_MEM_reg[5][12]  ( .D(n11380), .CK(N28803), .QN(n9887) );
  DFF_X1 \CACHE_MEM_reg[5][11]  ( .D(n11379), .CK(N28803), .QN(n9903) );
  DFF_X1 \CACHE_MEM_reg[5][10]  ( .D(n11378), .CK(N28803), .QN(n9919) );
  DFF_X1 \CACHE_MEM_reg[5][9]  ( .D(n11377), .CK(N28803), .QN(n9935) );
  DFF_X1 \CACHE_MEM_reg[5][8]  ( .D(n11376), .CK(N28803), .QN(n9951) );
  DFF_X1 \CACHE_MEM_reg[5][7]  ( .D(n11375), .CK(N28803), .QN(n9967) );
  DFF_X1 \CACHE_MEM_reg[5][6]  ( .D(n11374), .CK(N28803), .QN(n9983) );
  DFF_X1 \CACHE_MEM_reg[5][5]  ( .D(n11373), .CK(N28803), .QN(n9999) );
  DFF_X1 \CACHE_MEM_reg[5][4]  ( .D(n11372), .CK(N28803), .QN(n10015) );
  DFF_X1 \CACHE_MEM_reg[5][3]  ( .D(n11371), .CK(N28803), .QN(n10031) );
  DFF_X1 \CACHE_MEM_reg[5][2]  ( .D(n11370), .CK(N28803), .QN(n10047) );
  DFF_X1 \CACHE_MEM_reg[5][1]  ( .D(n11369), .CK(N28803), .QN(n10063) );
  DFF_X1 \CACHE_MEM_reg[5][0]  ( .D(n11368), .CK(N28803), .QN(n10079) );
  DFF_X1 \CACHE_MEM_reg[4][255]  ( .D(n11367), .CK(N28803), .QN(n5995) );
  DFF_X1 \CACHE_MEM_reg[4][254]  ( .D(n11366), .CK(N28803), .QN(n6011) );
  DFF_X1 \CACHE_MEM_reg[4][253]  ( .D(n11365), .CK(N28803), .QN(n6027) );
  DFF_X1 \CACHE_MEM_reg[4][252]  ( .D(n11364), .CK(N28803), .QN(n6043) );
  DFF_X1 \CACHE_MEM_reg[4][251]  ( .D(n11363), .CK(N28803), .QN(n6059) );
  DFF_X1 \CACHE_MEM_reg[4][250]  ( .D(n11362), .CK(N28803), .QN(n6075) );
  DFF_X1 \CACHE_MEM_reg[4][249]  ( .D(n11361), .CK(N28803), .QN(n6091) );
  DFF_X1 \CACHE_MEM_reg[4][248]  ( .D(n11360), .CK(N28803), .QN(n6107) );
  DFF_X1 \CACHE_MEM_reg[4][247]  ( .D(n11359), .CK(N28803), .QN(n6123) );
  DFF_X1 \CACHE_MEM_reg[4][246]  ( .D(n11358), .CK(N28803), .QN(n6139) );
  DFF_X1 \CACHE_MEM_reg[4][245]  ( .D(n11357), .CK(N28803), .QN(n6155) );
  DFF_X1 \CACHE_MEM_reg[4][244]  ( .D(n11356), .CK(N28803), .QN(n6171) );
  DFF_X1 \CACHE_MEM_reg[4][243]  ( .D(n11355), .CK(N28803), .QN(n6187) );
  DFF_X1 \CACHE_MEM_reg[4][242]  ( .D(n11354), .CK(N28803), .QN(n6203) );
  DFF_X1 \CACHE_MEM_reg[4][241]  ( .D(n11353), .CK(N28803), .QN(n6219) );
  DFF_X1 \CACHE_MEM_reg[4][240]  ( .D(n11352), .CK(N28803), .QN(n6235) );
  DFF_X1 \CACHE_MEM_reg[4][239]  ( .D(n11351), .CK(N28803), .QN(n6251) );
  DFF_X1 \CACHE_MEM_reg[4][238]  ( .D(n11350), .CK(N28803), .QN(n6267) );
  DFF_X1 \CACHE_MEM_reg[4][237]  ( .D(n11349), .CK(N28803), .QN(n6283) );
  DFF_X1 \CACHE_MEM_reg[4][236]  ( .D(n11348), .CK(N28803), .QN(n6299) );
  DFF_X1 \CACHE_MEM_reg[4][235]  ( .D(n11347), .CK(N28803), .QN(n6315) );
  DFF_X1 \CACHE_MEM_reg[4][234]  ( .D(n11346), .CK(N28803), .QN(n6331) );
  DFF_X1 \CACHE_MEM_reg[4][233]  ( .D(n11345), .CK(N28803), .QN(n6347) );
  DFF_X1 \CACHE_MEM_reg[4][232]  ( .D(n11344), .CK(N28803), .QN(n6363) );
  DFF_X1 \CACHE_MEM_reg[4][231]  ( .D(n11343), .CK(N28803), .QN(n6379) );
  DFF_X1 \CACHE_MEM_reg[4][230]  ( .D(n11342), .CK(N28803), .QN(n6395) );
  DFF_X1 \CACHE_MEM_reg[4][229]  ( .D(n11341), .CK(N28803), .QN(n6411) );
  DFF_X1 \CACHE_MEM_reg[4][228]  ( .D(n11340), .CK(N28803), .QN(n6427) );
  DFF_X1 \CACHE_MEM_reg[4][227]  ( .D(n11339), .CK(N28803), .QN(n6443) );
  DFF_X1 \CACHE_MEM_reg[4][226]  ( .D(n11338), .CK(N28803), .QN(n6459) );
  DFF_X1 \CACHE_MEM_reg[4][225]  ( .D(n11337), .CK(N28803), .QN(n6475) );
  DFF_X1 \CACHE_MEM_reg[4][224]  ( .D(n11336), .CK(N28803), .QN(n6491) );
  DFF_X1 \CACHE_MEM_reg[4][223]  ( .D(n11335), .CK(N28803), .QN(n6507) );
  DFF_X1 \CACHE_MEM_reg[4][222]  ( .D(n11334), .CK(N28803), .QN(n6523) );
  DFF_X1 \CACHE_MEM_reg[4][221]  ( .D(n11333), .CK(N28803), .QN(n6539) );
  DFF_X1 \CACHE_MEM_reg[4][220]  ( .D(n11332), .CK(N28803), .QN(n6555) );
  DFF_X1 \CACHE_MEM_reg[4][219]  ( .D(n11331), .CK(N28803), .QN(n6571) );
  DFF_X1 \CACHE_MEM_reg[4][218]  ( .D(n11330), .CK(N28803), .QN(n6587) );
  DFF_X1 \CACHE_MEM_reg[4][217]  ( .D(n11329), .CK(N28803), .QN(n6603) );
  DFF_X1 \CACHE_MEM_reg[4][216]  ( .D(n11328), .CK(N28803), .QN(n6619) );
  DFF_X1 \CACHE_MEM_reg[4][215]  ( .D(n11327), .CK(N28803), .QN(n6635) );
  DFF_X1 \CACHE_MEM_reg[4][214]  ( .D(n11326), .CK(N28803), .QN(n6651) );
  DFF_X1 \CACHE_MEM_reg[4][213]  ( .D(n11325), .CK(N28803), .QN(n6667) );
  DFF_X1 \CACHE_MEM_reg[4][212]  ( .D(n11324), .CK(N28803), .QN(n6683) );
  DFF_X1 \CACHE_MEM_reg[4][211]  ( .D(n11323), .CK(N28803), .QN(n6699) );
  DFF_X1 \CACHE_MEM_reg[4][210]  ( .D(n11322), .CK(N28803), .QN(n6715) );
  DFF_X1 \CACHE_MEM_reg[4][209]  ( .D(n11321), .CK(N28803), .QN(n6731) );
  DFF_X1 \CACHE_MEM_reg[4][208]  ( .D(n11320), .CK(N28803), .QN(n6747) );
  DFF_X1 \CACHE_MEM_reg[4][207]  ( .D(n11319), .CK(N28803), .QN(n6763) );
  DFF_X1 \CACHE_MEM_reg[4][206]  ( .D(n11318), .CK(N28803), .QN(n6779) );
  DFF_X1 \CACHE_MEM_reg[4][205]  ( .D(n11317), .CK(N28803), .QN(n6795) );
  DFF_X1 \CACHE_MEM_reg[4][204]  ( .D(n11316), .CK(N28803), .QN(n6811) );
  DFF_X1 \CACHE_MEM_reg[4][203]  ( .D(n11315), .CK(N28803), .QN(n6827) );
  DFF_X1 \CACHE_MEM_reg[4][202]  ( .D(n11314), .CK(N28803), .QN(n6843) );
  DFF_X1 \CACHE_MEM_reg[4][201]  ( .D(n11313), .CK(N28803), .QN(n6859) );
  DFF_X1 \CACHE_MEM_reg[4][200]  ( .D(n11312), .CK(N28803), .QN(n6875) );
  DFF_X1 \CACHE_MEM_reg[4][199]  ( .D(n11311), .CK(N28803), .QN(n6891) );
  DFF_X1 \CACHE_MEM_reg[4][198]  ( .D(n11310), .CK(N28803), .QN(n6907) );
  DFF_X1 \CACHE_MEM_reg[4][197]  ( .D(n11309), .CK(N28803), .QN(n6923) );
  DFF_X1 \CACHE_MEM_reg[4][196]  ( .D(n11308), .CK(N28803), .QN(n6939) );
  DFF_X1 \CACHE_MEM_reg[4][195]  ( .D(n11307), .CK(N28803), .QN(n6955) );
  DFF_X1 \CACHE_MEM_reg[4][194]  ( .D(n11306), .CK(N28803), .QN(n6971) );
  DFF_X1 \CACHE_MEM_reg[4][193]  ( .D(n11305), .CK(N28803), .QN(n6987) );
  DFF_X1 \CACHE_MEM_reg[4][192]  ( .D(n11304), .CK(N28803), .QN(n7003) );
  DFF_X1 \CACHE_MEM_reg[4][191]  ( .D(n11303), .CK(N28803), .QN(n7019) );
  DFF_X1 \CACHE_MEM_reg[4][190]  ( .D(n11302), .CK(N28803), .QN(n7035) );
  DFF_X1 \CACHE_MEM_reg[4][189]  ( .D(n11301), .CK(N28803), .QN(n7051) );
  DFF_X1 \CACHE_MEM_reg[4][188]  ( .D(n11300), .CK(N28803), .QN(n7067) );
  DFF_X1 \CACHE_MEM_reg[4][187]  ( .D(n11299), .CK(N28803), .QN(n7083) );
  DFF_X1 \CACHE_MEM_reg[4][186]  ( .D(n11298), .CK(N28803), .QN(n7099) );
  DFF_X1 \CACHE_MEM_reg[4][185]  ( .D(n11297), .CK(N28803), .QN(n7115) );
  DFF_X1 \CACHE_MEM_reg[4][184]  ( .D(n11296), .CK(N28803), .QN(n7131) );
  DFF_X1 \CACHE_MEM_reg[4][183]  ( .D(n11295), .CK(N28803), .QN(n7147) );
  DFF_X1 \CACHE_MEM_reg[4][182]  ( .D(n11294), .CK(N28803), .QN(n7163) );
  DFF_X1 \CACHE_MEM_reg[4][181]  ( .D(n11293), .CK(N28803), .QN(n7179) );
  DFF_X1 \CACHE_MEM_reg[4][180]  ( .D(n11292), .CK(N28803), .QN(n7195) );
  DFF_X1 \CACHE_MEM_reg[4][179]  ( .D(n11291), .CK(N28803), .QN(n7211) );
  DFF_X1 \CACHE_MEM_reg[4][178]  ( .D(n11290), .CK(N28803), .QN(n7227) );
  DFF_X1 \CACHE_MEM_reg[4][177]  ( .D(n11289), .CK(N28803), .QN(n7243) );
  DFF_X1 \CACHE_MEM_reg[4][176]  ( .D(n11288), .CK(N28803), .QN(n7259) );
  DFF_X1 \CACHE_MEM_reg[4][175]  ( .D(n11287), .CK(N28803), .QN(n7275) );
  DFF_X1 \CACHE_MEM_reg[4][174]  ( .D(n11286), .CK(N28803), .QN(n7291) );
  DFF_X1 \CACHE_MEM_reg[4][173]  ( .D(n11285), .CK(N28803), .QN(n7307) );
  DFF_X1 \CACHE_MEM_reg[4][172]  ( .D(n11284), .CK(N28803), .QN(n7323) );
  DFF_X1 \CACHE_MEM_reg[4][171]  ( .D(n11283), .CK(N28803), .QN(n7339) );
  DFF_X1 \CACHE_MEM_reg[4][170]  ( .D(n11282), .CK(N28803), .QN(n7355) );
  DFF_X1 \CACHE_MEM_reg[4][169]  ( .D(n11281), .CK(N28803), .QN(n7371) );
  DFF_X1 \CACHE_MEM_reg[4][168]  ( .D(n11280), .CK(N28803), .QN(n7387) );
  DFF_X1 \CACHE_MEM_reg[4][167]  ( .D(n11279), .CK(N28803), .QN(n7403) );
  DFF_X1 \CACHE_MEM_reg[4][166]  ( .D(n11278), .CK(N28803), .QN(n7419) );
  DFF_X1 \CACHE_MEM_reg[4][165]  ( .D(n11277), .CK(N28803), .QN(n7435) );
  DFF_X1 \CACHE_MEM_reg[4][164]  ( .D(n11276), .CK(N28803), .QN(n7451) );
  DFF_X1 \CACHE_MEM_reg[4][163]  ( .D(n11275), .CK(N28803), .QN(n7467) );
  DFF_X1 \CACHE_MEM_reg[4][162]  ( .D(n11274), .CK(N28803), .QN(n7483) );
  DFF_X1 \CACHE_MEM_reg[4][161]  ( .D(n11273), .CK(N28803), .QN(n7499) );
  DFF_X1 \CACHE_MEM_reg[4][160]  ( .D(n11272), .CK(N28803), .QN(n7515) );
  DFF_X1 \CACHE_MEM_reg[4][159]  ( .D(n11271), .CK(N28803), .QN(n7531) );
  DFF_X1 \CACHE_MEM_reg[4][158]  ( .D(n11270), .CK(N28803), .QN(n7547) );
  DFF_X1 \CACHE_MEM_reg[4][157]  ( .D(n11269), .CK(N28803), .QN(n7563) );
  DFF_X1 \CACHE_MEM_reg[4][156]  ( .D(n11268), .CK(N28803), .QN(n7579) );
  DFF_X1 \CACHE_MEM_reg[4][155]  ( .D(n11267), .CK(N28803), .QN(n7595) );
  DFF_X1 \CACHE_MEM_reg[4][154]  ( .D(n11266), .CK(N28803), .QN(n7611) );
  DFF_X1 \CACHE_MEM_reg[4][153]  ( .D(n11265), .CK(N28803), .QN(n7627) );
  DFF_X1 \CACHE_MEM_reg[4][152]  ( .D(n11264), .CK(N28803), .QN(n7643) );
  DFF_X1 \CACHE_MEM_reg[4][151]  ( .D(n11263), .CK(N28803), .QN(n7659) );
  DFF_X1 \CACHE_MEM_reg[4][150]  ( .D(n11262), .CK(N28803), .QN(n7675) );
  DFF_X1 \CACHE_MEM_reg[4][149]  ( .D(n11261), .CK(N28803), .QN(n7691) );
  DFF_X1 \CACHE_MEM_reg[4][148]  ( .D(n11260), .CK(N28803), .QN(n7707) );
  DFF_X1 \CACHE_MEM_reg[4][147]  ( .D(n11259), .CK(N28803), .QN(n7723) );
  DFF_X1 \CACHE_MEM_reg[4][146]  ( .D(n11258), .CK(N28803), .QN(n7739) );
  DFF_X1 \CACHE_MEM_reg[4][145]  ( .D(n11257), .CK(N28803), .QN(n7755) );
  DFF_X1 \CACHE_MEM_reg[4][144]  ( .D(n11256), .CK(N28803), .QN(n7771) );
  DFF_X1 \CACHE_MEM_reg[4][143]  ( .D(n11255), .CK(N28803), .QN(n7787) );
  DFF_X1 \CACHE_MEM_reg[4][142]  ( .D(n11254), .CK(N28803), .QN(n7803) );
  DFF_X1 \CACHE_MEM_reg[4][141]  ( .D(n11253), .CK(N28803), .QN(n7819) );
  DFF_X1 \CACHE_MEM_reg[4][140]  ( .D(n11252), .CK(N28803), .QN(n7835) );
  DFF_X1 \CACHE_MEM_reg[4][139]  ( .D(n11251), .CK(N28803), .QN(n7851) );
  DFF_X1 \CACHE_MEM_reg[4][138]  ( .D(n11250), .CK(N28803), .QN(n7867) );
  DFF_X1 \CACHE_MEM_reg[4][137]  ( .D(n11249), .CK(N28803), .QN(n7883) );
  DFF_X1 \CACHE_MEM_reg[4][136]  ( .D(n11248), .CK(N28803), .QN(n7899) );
  DFF_X1 \CACHE_MEM_reg[4][135]  ( .D(n11247), .CK(N28803), .QN(n7915) );
  DFF_X1 \CACHE_MEM_reg[4][134]  ( .D(n11246), .CK(N28803), .QN(n7931) );
  DFF_X1 \CACHE_MEM_reg[4][133]  ( .D(n11245), .CK(N28803), .QN(n7947) );
  DFF_X1 \CACHE_MEM_reg[4][132]  ( .D(n11244), .CK(N28803), .QN(n7963) );
  DFF_X1 \CACHE_MEM_reg[4][131]  ( .D(n11243), .CK(N28803), .QN(n7979) );
  DFF_X1 \CACHE_MEM_reg[4][130]  ( .D(n11242), .CK(N28803), .QN(n7995) );
  DFF_X1 \CACHE_MEM_reg[4][129]  ( .D(n11241), .CK(N28803), .QN(n8011) );
  DFF_X1 \CACHE_MEM_reg[4][128]  ( .D(n11240), .CK(N28803), .QN(n8027) );
  DFF_X1 \CACHE_MEM_reg[4][127]  ( .D(n11239), .CK(N28803), .QN(n8043) );
  DFF_X1 \CACHE_MEM_reg[4][126]  ( .D(n11238), .CK(N28803), .QN(n8059) );
  DFF_X1 \CACHE_MEM_reg[4][125]  ( .D(n11237), .CK(N28803), .QN(n8075) );
  DFF_X1 \CACHE_MEM_reg[4][124]  ( .D(n11236), .CK(N28803), .QN(n8091) );
  DFF_X1 \CACHE_MEM_reg[4][123]  ( .D(n11235), .CK(N28803), .QN(n8107) );
  DFF_X1 \CACHE_MEM_reg[4][122]  ( .D(n11234), .CK(N28803), .QN(n8123) );
  DFF_X1 \CACHE_MEM_reg[4][121]  ( .D(n11233), .CK(N28803), .QN(n8139) );
  DFF_X1 \CACHE_MEM_reg[4][120]  ( .D(n11232), .CK(N28803), .QN(n8155) );
  DFF_X1 \CACHE_MEM_reg[4][119]  ( .D(n11231), .CK(N28803), .QN(n8171) );
  DFF_X1 \CACHE_MEM_reg[4][118]  ( .D(n11230), .CK(N28803), .QN(n8187) );
  DFF_X1 \CACHE_MEM_reg[4][117]  ( .D(n11229), .CK(N28803), .QN(n8203) );
  DFF_X1 \CACHE_MEM_reg[4][116]  ( .D(n11228), .CK(N28803), .QN(n8219) );
  DFF_X1 \CACHE_MEM_reg[4][115]  ( .D(n11227), .CK(N28803), .QN(n8235) );
  DFF_X1 \CACHE_MEM_reg[4][114]  ( .D(n11226), .CK(N28803), .QN(n8251) );
  DFF_X1 \CACHE_MEM_reg[4][113]  ( .D(n11225), .CK(N28803), .QN(n8267) );
  DFF_X1 \CACHE_MEM_reg[4][112]  ( .D(n11224), .CK(N28803), .QN(n8283) );
  DFF_X1 \CACHE_MEM_reg[4][111]  ( .D(n11223), .CK(N28803), .QN(n8299) );
  DFF_X1 \CACHE_MEM_reg[4][110]  ( .D(n11222), .CK(N28803), .QN(n8315) );
  DFF_X1 \CACHE_MEM_reg[4][109]  ( .D(n11221), .CK(N28803), .QN(n8331) );
  DFF_X1 \CACHE_MEM_reg[4][108]  ( .D(n11220), .CK(N28803), .QN(n8347) );
  DFF_X1 \CACHE_MEM_reg[4][107]  ( .D(n11219), .CK(N28803), .QN(n8363) );
  DFF_X1 \CACHE_MEM_reg[4][106]  ( .D(n11218), .CK(N28803), .QN(n8379) );
  DFF_X1 \CACHE_MEM_reg[4][105]  ( .D(n11217), .CK(N28803), .QN(n8395) );
  DFF_X1 \CACHE_MEM_reg[4][104]  ( .D(n11216), .CK(N28803), .QN(n8411) );
  DFF_X1 \CACHE_MEM_reg[4][103]  ( .D(n11215), .CK(N28803), .QN(n8427) );
  DFF_X1 \CACHE_MEM_reg[4][102]  ( .D(n11214), .CK(N28803), .QN(n8443) );
  DFF_X1 \CACHE_MEM_reg[4][101]  ( .D(n11213), .CK(N28803), .QN(n8459) );
  DFF_X1 \CACHE_MEM_reg[4][100]  ( .D(n11212), .CK(N28803), .QN(n8475) );
  DFF_X1 \CACHE_MEM_reg[4][99]  ( .D(n11211), .CK(N28803), .QN(n8491) );
  DFF_X1 \CACHE_MEM_reg[4][98]  ( .D(n11210), .CK(N28803), .QN(n8507) );
  DFF_X1 \CACHE_MEM_reg[4][97]  ( .D(n11209), .CK(N28803), .QN(n8523) );
  DFF_X1 \CACHE_MEM_reg[4][96]  ( .D(n11208), .CK(N28803), .QN(n8539) );
  DFF_X1 \CACHE_MEM_reg[4][95]  ( .D(n11207), .CK(N28803), .QN(n8555) );
  DFF_X1 \CACHE_MEM_reg[4][94]  ( .D(n11206), .CK(N28803), .QN(n8571) );
  DFF_X1 \CACHE_MEM_reg[4][93]  ( .D(n11205), .CK(N28803), .QN(n8587) );
  DFF_X1 \CACHE_MEM_reg[4][92]  ( .D(n11204), .CK(N28803), .QN(n8603) );
  DFF_X1 \CACHE_MEM_reg[4][91]  ( .D(n11203), .CK(N28803), .QN(n8619) );
  DFF_X1 \CACHE_MEM_reg[4][90]  ( .D(n11202), .CK(N28803), .QN(n8635) );
  DFF_X1 \CACHE_MEM_reg[4][89]  ( .D(n11201), .CK(N28803), .QN(n8651) );
  DFF_X1 \CACHE_MEM_reg[4][88]  ( .D(n11200), .CK(N28803), .QN(n8667) );
  DFF_X1 \CACHE_MEM_reg[4][87]  ( .D(n11199), .CK(N28803), .QN(n8683) );
  DFF_X1 \CACHE_MEM_reg[4][86]  ( .D(n11198), .CK(N28803), .QN(n8699) );
  DFF_X1 \CACHE_MEM_reg[4][85]  ( .D(n11197), .CK(N28803), .QN(n8715) );
  DFF_X1 \CACHE_MEM_reg[4][84]  ( .D(n11196), .CK(N28803), .QN(n8731) );
  DFF_X1 \CACHE_MEM_reg[4][83]  ( .D(n11195), .CK(N28803), .QN(n8747) );
  DFF_X1 \CACHE_MEM_reg[4][82]  ( .D(n11194), .CK(N28803), .QN(n8763) );
  DFF_X1 \CACHE_MEM_reg[4][81]  ( .D(n11193), .CK(N28803), .QN(n8779) );
  DFF_X1 \CACHE_MEM_reg[4][80]  ( .D(n11192), .CK(N28803), .QN(n8795) );
  DFF_X1 \CACHE_MEM_reg[4][79]  ( .D(n11191), .CK(N28803), .QN(n8811) );
  DFF_X1 \CACHE_MEM_reg[4][78]  ( .D(n11190), .CK(N28803), .QN(n8827) );
  DFF_X1 \CACHE_MEM_reg[4][77]  ( .D(n11189), .CK(N28803), .QN(n8843) );
  DFF_X1 \CACHE_MEM_reg[4][76]  ( .D(n11188), .CK(N28803), .QN(n8859) );
  DFF_X1 \CACHE_MEM_reg[4][75]  ( .D(n11187), .CK(N28803), .QN(n8875) );
  DFF_X1 \CACHE_MEM_reg[4][74]  ( .D(n11186), .CK(N28803), .QN(n8891) );
  DFF_X1 \CACHE_MEM_reg[4][73]  ( .D(n11185), .CK(N28803), .QN(n8907) );
  DFF_X1 \CACHE_MEM_reg[4][72]  ( .D(n11184), .CK(N28803), .QN(n8923) );
  DFF_X1 \CACHE_MEM_reg[4][71]  ( .D(n11183), .CK(N28803), .QN(n8939) );
  DFF_X1 \CACHE_MEM_reg[4][70]  ( .D(n11182), .CK(N28803), .QN(n8955) );
  DFF_X1 \CACHE_MEM_reg[4][69]  ( .D(n11181), .CK(N28803), .QN(n8971) );
  DFF_X1 \CACHE_MEM_reg[4][68]  ( .D(n11180), .CK(N28803), .QN(n8987) );
  DFF_X1 \CACHE_MEM_reg[4][67]  ( .D(n11179), .CK(N28803), .QN(n9003) );
  DFF_X1 \CACHE_MEM_reg[4][66]  ( .D(n11178), .CK(N28803), .QN(n9019) );
  DFF_X1 \CACHE_MEM_reg[4][65]  ( .D(n11177), .CK(N28803), .QN(n9035) );
  DFF_X1 \CACHE_MEM_reg[4][64]  ( .D(n11176), .CK(N28803), .QN(n9051) );
  DFF_X1 \CACHE_MEM_reg[4][63]  ( .D(n11175), .CK(N28803), .QN(n9067) );
  DFF_X1 \CACHE_MEM_reg[4][62]  ( .D(n11174), .CK(N28803), .QN(n9083) );
  DFF_X1 \CACHE_MEM_reg[4][61]  ( .D(n11173), .CK(N28803), .QN(n9099) );
  DFF_X1 \CACHE_MEM_reg[4][60]  ( .D(n11172), .CK(N28803), .QN(n9115) );
  DFF_X1 \CACHE_MEM_reg[4][59]  ( .D(n11171), .CK(N28803), .QN(n9131) );
  DFF_X1 \CACHE_MEM_reg[4][58]  ( .D(n11170), .CK(N28803), .QN(n9147) );
  DFF_X1 \CACHE_MEM_reg[4][57]  ( .D(n11169), .CK(N28803), .QN(n9163) );
  DFF_X1 \CACHE_MEM_reg[4][56]  ( .D(n11168), .CK(N28803), .QN(n9179) );
  DFF_X1 \CACHE_MEM_reg[4][55]  ( .D(n11167), .CK(N28803), .QN(n9195) );
  DFF_X1 \CACHE_MEM_reg[4][54]  ( .D(n11166), .CK(N28803), .QN(n9211) );
  DFF_X1 \CACHE_MEM_reg[4][53]  ( .D(n11165), .CK(N28803), .QN(n9227) );
  DFF_X1 \CACHE_MEM_reg[4][52]  ( .D(n11164), .CK(N28803), .QN(n9243) );
  DFF_X1 \CACHE_MEM_reg[4][51]  ( .D(n11163), .CK(N28803), .QN(n9259) );
  DFF_X1 \CACHE_MEM_reg[4][50]  ( .D(n11162), .CK(N28803), .QN(n9275) );
  DFF_X1 \CACHE_MEM_reg[4][49]  ( .D(n11161), .CK(N28803), .QN(n9291) );
  DFF_X1 \CACHE_MEM_reg[4][48]  ( .D(n11160), .CK(N28803), .QN(n9307) );
  DFF_X1 \CACHE_MEM_reg[4][47]  ( .D(n11159), .CK(N28803), .QN(n9323) );
  DFF_X1 \CACHE_MEM_reg[4][46]  ( .D(n11158), .CK(N28803), .QN(n9339) );
  DFF_X1 \CACHE_MEM_reg[4][45]  ( .D(n11157), .CK(N28803), .QN(n9355) );
  DFF_X1 \CACHE_MEM_reg[4][44]  ( .D(n11156), .CK(N28803), .QN(n9371) );
  DFF_X1 \CACHE_MEM_reg[4][43]  ( .D(n11155), .CK(N28803), .QN(n9387) );
  DFF_X1 \CACHE_MEM_reg[4][42]  ( .D(n11154), .CK(N28803), .QN(n9403) );
  DFF_X1 \CACHE_MEM_reg[4][41]  ( .D(n11153), .CK(N28803), .QN(n9419) );
  DFF_X1 \CACHE_MEM_reg[4][40]  ( .D(n11152), .CK(N28803), .QN(n9435) );
  DFF_X1 \CACHE_MEM_reg[4][39]  ( .D(n11151), .CK(N28803), .QN(n9451) );
  DFF_X1 \CACHE_MEM_reg[4][38]  ( .D(n11150), .CK(N28803), .QN(n9467) );
  DFF_X1 \CACHE_MEM_reg[4][37]  ( .D(n11149), .CK(N28803), .QN(n9483) );
  DFF_X1 \CACHE_MEM_reg[4][36]  ( .D(n11148), .CK(N28803), .QN(n9499) );
  DFF_X1 \CACHE_MEM_reg[4][35]  ( .D(n11147), .CK(N28803), .QN(n9515) );
  DFF_X1 \CACHE_MEM_reg[4][34]  ( .D(n11146), .CK(N28803), .QN(n9531) );
  DFF_X1 \CACHE_MEM_reg[4][33]  ( .D(n11145), .CK(N28803), .QN(n9547) );
  DFF_X1 \CACHE_MEM_reg[4][32]  ( .D(n11144), .CK(N28803), .QN(n9563) );
  DFF_X1 \CACHE_MEM_reg[4][31]  ( .D(n11143), .CK(N28803), .QN(n9579) );
  DFF_X1 \CACHE_MEM_reg[4][30]  ( .D(n11142), .CK(N28803), .QN(n9595) );
  DFF_X1 \CACHE_MEM_reg[4][29]  ( .D(n11141), .CK(N28803), .QN(n9611) );
  DFF_X1 \CACHE_MEM_reg[4][28]  ( .D(n11140), .CK(N28803), .QN(n9627) );
  DFF_X1 \CACHE_MEM_reg[4][27]  ( .D(n11139), .CK(N28803), .QN(n9643) );
  DFF_X1 \CACHE_MEM_reg[4][26]  ( .D(n11138), .CK(N28803), .QN(n9659) );
  DFF_X1 \CACHE_MEM_reg[4][25]  ( .D(n11137), .CK(N28803), .QN(n9675) );
  DFF_X1 \CACHE_MEM_reg[4][24]  ( .D(n11136), .CK(N28803), .QN(n9691) );
  DFF_X1 \CACHE_MEM_reg[4][23]  ( .D(n11135), .CK(N28803), .QN(n9707) );
  DFF_X1 \CACHE_MEM_reg[4][22]  ( .D(n11134), .CK(N28803), .QN(n9723) );
  DFF_X1 \CACHE_MEM_reg[4][21]  ( .D(n11133), .CK(N28803), .QN(n9739) );
  DFF_X1 \CACHE_MEM_reg[4][20]  ( .D(n11132), .CK(N28803), .QN(n9755) );
  DFF_X1 \CACHE_MEM_reg[4][19]  ( .D(n11131), .CK(N28803), .QN(n9771) );
  DFF_X1 \CACHE_MEM_reg[4][18]  ( .D(n11130), .CK(N28803), .QN(n9787) );
  DFF_X1 \CACHE_MEM_reg[4][17]  ( .D(n11129), .CK(N28803), .QN(n9803) );
  DFF_X1 \CACHE_MEM_reg[4][16]  ( .D(n11128), .CK(N28803), .QN(n9819) );
  DFF_X1 \CACHE_MEM_reg[4][15]  ( .D(n11127), .CK(N28803), .QN(n9835) );
  DFF_X1 \CACHE_MEM_reg[4][14]  ( .D(n11126), .CK(N28803), .QN(n9851) );
  DFF_X1 \CACHE_MEM_reg[4][13]  ( .D(n11125), .CK(N28803), .QN(n9867) );
  DFF_X1 \CACHE_MEM_reg[4][12]  ( .D(n11124), .CK(N28803), .QN(n9883) );
  DFF_X1 \CACHE_MEM_reg[4][11]  ( .D(n11123), .CK(N28803), .QN(n9899) );
  DFF_X1 \CACHE_MEM_reg[4][10]  ( .D(n11122), .CK(N28803), .QN(n9915) );
  DFF_X1 \CACHE_MEM_reg[4][9]  ( .D(n11121), .CK(N28803), .QN(n9931) );
  DFF_X1 \CACHE_MEM_reg[4][8]  ( .D(n11120), .CK(N28803), .QN(n9947) );
  DFF_X1 \CACHE_MEM_reg[4][7]  ( .D(n11119), .CK(N28803), .QN(n9963) );
  DFF_X1 \CACHE_MEM_reg[4][6]  ( .D(n11118), .CK(N28803), .QN(n9979) );
  DFF_X1 \CACHE_MEM_reg[4][5]  ( .D(n11117), .CK(N28803), .QN(n9995) );
  DFF_X1 \CACHE_MEM_reg[4][4]  ( .D(n11116), .CK(N28803), .QN(n10011) );
  DFF_X1 \CACHE_MEM_reg[4][3]  ( .D(n11115), .CK(N28803), .QN(n10027) );
  DFF_X1 \CACHE_MEM_reg[4][2]  ( .D(n11114), .CK(N28803), .QN(n10043) );
  DFF_X1 \CACHE_MEM_reg[4][1]  ( .D(n11113), .CK(N28803), .QN(n10059) );
  DFF_X1 \CACHE_MEM_reg[4][0]  ( .D(n11112), .CK(N28803), .QN(n10075) );
  DFF_X1 \CACHE_MEM_reg[3][255]  ( .D(n11111), .CK(N28803), .Q(n2882), .QN(
        n6005) );
  DFF_X1 \CACHE_MEM_reg[3][254]  ( .D(n11110), .CK(N28803), .Q(n2871), .QN(
        n6021) );
  DFF_X1 \CACHE_MEM_reg[3][253]  ( .D(n11109), .CK(N28803), .Q(n2854), .QN(
        n6037) );
  DFF_X1 \CACHE_MEM_reg[3][252]  ( .D(n11108), .CK(N28803), .Q(n2843), .QN(
        n6053) );
  DFF_X1 \CACHE_MEM_reg[3][251]  ( .D(n11107), .CK(N28803), .Q(n2821), .QN(
        n6069) );
  DFF_X1 \CACHE_MEM_reg[3][250]  ( .D(n11106), .CK(N28803), .Q(n2810), .QN(
        n6085) );
  DFF_X1 \CACHE_MEM_reg[3][249]  ( .D(n11105), .CK(N28803), .Q(n2797), .QN(
        n6101) );
  DFF_X1 \CACHE_MEM_reg[3][248]  ( .D(n11104), .CK(N28803), .Q(n2782), .QN(
        n6117) );
  DFF_X1 \CACHE_MEM_reg[3][247]  ( .D(n11103), .CK(N28803), .Q(n2769), .QN(
        n6133) );
  DFF_X1 \CACHE_MEM_reg[3][246]  ( .D(n11102), .CK(N28803), .Q(n2758), .QN(
        n6149) );
  DFF_X1 \CACHE_MEM_reg[3][245]  ( .D(n11101), .CK(N28803), .Q(n2741), .QN(
        n6165) );
  DFF_X1 \CACHE_MEM_reg[3][244]  ( .D(n11100), .CK(N28803), .Q(n2730), .QN(
        n6181) );
  DFF_X1 \CACHE_MEM_reg[3][243]  ( .D(n11099), .CK(N28803), .Q(n2713), .QN(
        n6197) );
  DFF_X1 \CACHE_MEM_reg[3][242]  ( .D(n11098), .CK(N28803), .Q(n2702), .QN(
        n6213) );
  DFF_X1 \CACHE_MEM_reg[3][241]  ( .D(n11097), .CK(N28803), .Q(n2689), .QN(
        n6229) );
  DFF_X1 \CACHE_MEM_reg[3][240]  ( .D(n11096), .CK(N28803), .Q(n3337), .QN(
        n6245) );
  DFF_X1 \CACHE_MEM_reg[3][239]  ( .D(n11095), .CK(N28803), .Q(n2661), .QN(
        n6261) );
  DFF_X1 \CACHE_MEM_reg[3][238]  ( .D(n11094), .CK(N28803), .Q(n2648), .QN(
        n6277) );
  DFF_X1 \CACHE_MEM_reg[3][237]  ( .D(n11093), .CK(N28803), .Q(n2633), .QN(
        n6293) );
  DFF_X1 \CACHE_MEM_reg[3][236]  ( .D(n11092), .CK(N28803), .Q(n2620), .QN(
        n6309) );
  DFF_X1 \CACHE_MEM_reg[3][235]  ( .D(n11091), .CK(N28803), .Q(n2609), .QN(
        n6325) );
  DFF_X1 \CACHE_MEM_reg[3][234]  ( .D(n11090), .CK(N28803), .Q(n2592), .QN(
        n6341) );
  DFF_X1 \CACHE_MEM_reg[3][233]  ( .D(n11089), .CK(N28803), .Q(n2581), .QN(
        n6357) );
  DFF_X1 \CACHE_MEM_reg[3][232]  ( .D(n11088), .CK(N28803), .Q(n2564), .QN(
        n6373) );
  DFF_X1 \CACHE_MEM_reg[3][231]  ( .D(n11087), .CK(N28803), .Q(n2553), .QN(
        n6389) );
  DFF_X1 \CACHE_MEM_reg[3][230]  ( .D(n11086), .CK(N28803), .Q(n2540), .QN(
        n6405) );
  DFF_X1 \CACHE_MEM_reg[3][229]  ( .D(n11085), .CK(N28803), .Q(n2520), .QN(
        n6421) );
  DFF_X1 \CACHE_MEM_reg[3][228]  ( .D(n11084), .CK(N28803), .Q(n2507), .QN(
        n6437) );
  DFF_X1 \CACHE_MEM_reg[3][227]  ( .D(n11083), .CK(N28803), .Q(n2496), .QN(
        n6453) );
  DFF_X1 \CACHE_MEM_reg[3][226]  ( .D(n11082), .CK(N28803), .Q(n2479), .QN(
        n6469) );
  DFF_X1 \CACHE_MEM_reg[3][225]  ( .D(n11081), .CK(N28803), .Q(n2468), .QN(
        n6485) );
  DFF_X1 \CACHE_MEM_reg[3][224]  ( .D(n11080), .CK(N28803), .Q(n2451), .QN(
        n6501) );
  DFF_X1 \CACHE_MEM_reg[3][223]  ( .D(n11079), .CK(N28803), .Q(n2887), .QN(
        n6517) );
  DFF_X1 \CACHE_MEM_reg[3][222]  ( .D(n11078), .CK(N28803), .Q(n2874), .QN(
        n6533) );
  DFF_X1 \CACHE_MEM_reg[3][221]  ( .D(n11077), .CK(N28803), .Q(n2859), .QN(
        n6549) );
  DFF_X1 \CACHE_MEM_reg[3][220]  ( .D(n11076), .CK(N28803), .Q(n2846), .QN(
        n6565) );
  DFF_X1 \CACHE_MEM_reg[3][219]  ( .D(n11075), .CK(N28803), .Q(n2835), .QN(
        n6581) );
  DFF_X1 \CACHE_MEM_reg[3][218]  ( .D(n11074), .CK(N28803), .Q(n2813), .QN(
        n6597) );
  DFF_X1 \CACHE_MEM_reg[3][217]  ( .D(n11073), .CK(N28803), .Q(n2802), .QN(
        n6613) );
  DFF_X1 \CACHE_MEM_reg[3][216]  ( .D(n11072), .CK(N28803), .Q(n2785), .QN(
        n6629) );
  DFF_X1 \CACHE_MEM_reg[3][215]  ( .D(n11071), .CK(N28803), .Q(n2774), .QN(
        n6645) );
  DFF_X1 \CACHE_MEM_reg[3][214]  ( .D(n11070), .CK(N28803), .Q(n2761), .QN(
        n6661) );
  DFF_X1 \CACHE_MEM_reg[3][213]  ( .D(n11069), .CK(N28803), .Q(n2746), .QN(
        n6677) );
  DFF_X1 \CACHE_MEM_reg[3][212]  ( .D(n11068), .CK(N28803), .Q(n2733), .QN(
        n6693) );
  DFF_X1 \CACHE_MEM_reg[3][211]  ( .D(n11067), .CK(N28803), .Q(n2722), .QN(
        n6709) );
  DFF_X1 \CACHE_MEM_reg[3][210]  ( .D(n11066), .CK(N28803), .Q(n2705), .QN(
        n6725) );
  DFF_X1 \CACHE_MEM_reg[3][209]  ( .D(n11065), .CK(N28803), .Q(n2694), .QN(
        n6741) );
  DFF_X1 \CACHE_MEM_reg[3][208]  ( .D(n11064), .CK(N28803), .Q(n2672), .QN(
        n6757) );
  DFF_X1 \CACHE_MEM_reg[3][207]  ( .D(n11063), .CK(N28803), .Q(n2664), .QN(
        n6773) );
  DFF_X1 \CACHE_MEM_reg[3][206]  ( .D(n11062), .CK(N28803), .Q(n2653), .QN(
        n6789) );
  DFF_X1 \CACHE_MEM_reg[3][205]  ( .D(n11061), .CK(N28803), .Q(n2636), .QN(
        n6805) );
  DFF_X1 \CACHE_MEM_reg[3][204]  ( .D(n11060), .CK(N28803), .Q(n2625), .QN(
        n6821) );
  DFF_X1 \CACHE_MEM_reg[3][203]  ( .D(n11059), .CK(N28803), .Q(n2612), .QN(
        n6837) );
  DFF_X1 \CACHE_MEM_reg[3][202]  ( .D(n11058), .CK(N28803), .Q(n2597), .QN(
        n6853) );
  DFF_X1 \CACHE_MEM_reg[3][201]  ( .D(n11057), .CK(N28803), .Q(n2584), .QN(
        n6869) );
  DFF_X1 \CACHE_MEM_reg[3][200]  ( .D(n11056), .CK(N28803), .Q(n2573), .QN(
        n6885) );
  DFF_X1 \CACHE_MEM_reg[3][199]  ( .D(n11055), .CK(N28803), .Q(n2556), .QN(
        n6901) );
  DFF_X1 \CACHE_MEM_reg[3][198]  ( .D(n11054), .CK(N28803), .Q(n2545), .QN(
        n6917) );
  DFF_X1 \CACHE_MEM_reg[3][197]  ( .D(n11053), .CK(N28803), .Q(n2523), .QN(
        n6933) );
  DFF_X1 \CACHE_MEM_reg[3][196]  ( .D(n11052), .CK(N28803), .Q(n2512), .QN(
        n6949) );
  DFF_X1 \CACHE_MEM_reg[3][195]  ( .D(n11051), .CK(N28803), .Q(n2499), .QN(
        n6965) );
  DFF_X1 \CACHE_MEM_reg[3][194]  ( .D(n11050), .CK(N28803), .Q(n2484), .QN(
        n6981) );
  DFF_X1 \CACHE_MEM_reg[3][193]  ( .D(n11049), .CK(N28803), .Q(n2471), .QN(
        n6997) );
  DFF_X1 \CACHE_MEM_reg[3][192]  ( .D(n11048), .CK(N28803), .Q(n2460), .QN(
        n7013) );
  DFF_X1 \CACHE_MEM_reg[3][191]  ( .D(n11047), .CK(N28803), .Q(n3329), .QN(
        n7029) );
  DFF_X1 \CACHE_MEM_reg[3][190]  ( .D(n11046), .CK(N28803), .Q(n3318), .QN(
        n7045) );
  DFF_X1 \CACHE_MEM_reg[3][189]  ( .D(n11045), .CK(N28803), .Q(n3301), .QN(
        n7061) );
  DFF_X1 \CACHE_MEM_reg[3][188]  ( .D(n11044), .CK(N28803), .Q(n3290), .QN(
        n7077) );
  DFF_X1 \CACHE_MEM_reg[3][187]  ( .D(n11043), .CK(N28803), .Q(n3268), .QN(
        n7093) );
  DFF_X1 \CACHE_MEM_reg[3][186]  ( .D(n11042), .CK(N28803), .Q(n3257), .QN(
        n7109) );
  DFF_X1 \CACHE_MEM_reg[3][185]  ( .D(n11041), .CK(N28803), .Q(n3244), .QN(
        n7125) );
  DFF_X1 \CACHE_MEM_reg[3][184]  ( .D(n11040), .CK(N28803), .Q(n3229), .QN(
        n7141) );
  DFF_X1 \CACHE_MEM_reg[3][183]  ( .D(n11039), .CK(N28803), .Q(n3216), .QN(
        n7157) );
  DFF_X1 \CACHE_MEM_reg[3][182]  ( .D(n11038), .CK(N28803), .Q(n3205), .QN(
        n7173) );
  DFF_X1 \CACHE_MEM_reg[3][181]  ( .D(n11037), .CK(N28803), .Q(n3188), .QN(
        n7189) );
  DFF_X1 \CACHE_MEM_reg[3][180]  ( .D(n11036), .CK(N28803), .Q(n3177), .QN(
        n7205) );
  DFF_X1 \CACHE_MEM_reg[3][179]  ( .D(n11035), .CK(N28803), .Q(n3160), .QN(
        n7221) );
  DFF_X1 \CACHE_MEM_reg[3][178]  ( .D(n11034), .CK(N28803), .Q(n3149), .QN(
        n7237) );
  DFF_X1 \CACHE_MEM_reg[3][177]  ( .D(n11033), .CK(N28803), .Q(n3136), .QN(
        n7253) );
  DFF_X1 \CACHE_MEM_reg[3][176]  ( .D(n11032), .CK(N28803), .Q(n3116), .QN(
        n7269) );
  DFF_X1 \CACHE_MEM_reg[3][175]  ( .D(n11031), .CK(N28803), .Q(n3103), .QN(
        n7285) );
  DFF_X1 \CACHE_MEM_reg[3][174]  ( .D(n11030), .CK(N28803), .Q(n3092), .QN(
        n7301) );
  DFF_X1 \CACHE_MEM_reg[3][173]  ( .D(n11029), .CK(N28803), .Q(n3075), .QN(
        n7317) );
  DFF_X1 \CACHE_MEM_reg[3][172]  ( .D(n11028), .CK(N28803), .Q(n3064), .QN(
        n7333) );
  DFF_X1 \CACHE_MEM_reg[3][171]  ( .D(n11027), .CK(N28803), .Q(n3047), .QN(
        n7349) );
  DFF_X1 \CACHE_MEM_reg[3][170]  ( .D(n11026), .CK(N28803), .Q(n3036), .QN(
        n7365) );
  DFF_X1 \CACHE_MEM_reg[3][169]  ( .D(n11025), .CK(N28803), .Q(n3023), .QN(
        n7381) );
  DFF_X1 \CACHE_MEM_reg[3][168]  ( .D(n11024), .CK(N28803), .Q(n3008), .QN(
        n7397) );
  DFF_X1 \CACHE_MEM_reg[3][167]  ( .D(n11023), .CK(N28803), .Q(n2995), .QN(
        n7413) );
  DFF_X1 \CACHE_MEM_reg[3][166]  ( .D(n11022), .CK(N28803), .Q(n2984), .QN(
        n7429) );
  DFF_X1 \CACHE_MEM_reg[3][165]  ( .D(n11021), .CK(N28803), .Q(n2962), .QN(
        n7445) );
  DFF_X1 \CACHE_MEM_reg[3][164]  ( .D(n11020), .CK(N28803), .Q(n2951), .QN(
        n7461) );
  DFF_X1 \CACHE_MEM_reg[3][163]  ( .D(n11019), .CK(N28803), .Q(n2934), .QN(
        n7477) );
  DFF_X1 \CACHE_MEM_reg[3][162]  ( .D(n11018), .CK(N28803), .Q(n2923), .QN(
        n7493) );
  DFF_X1 \CACHE_MEM_reg[3][161]  ( .D(n11017), .CK(N28803), .Q(n2910), .QN(
        n7509) );
  DFF_X1 \CACHE_MEM_reg[3][160]  ( .D(n11016), .CK(N28803), .Q(n2895), .QN(
        n7525) );
  DFF_X1 \CACHE_MEM_reg[3][159]  ( .D(n11015), .CK(N28803), .Q(n3334), .QN(
        n7541) );
  DFF_X1 \CACHE_MEM_reg[3][158]  ( .D(n11014), .CK(N28803), .Q(n3342), .QN(
        n7557) );
  DFF_X1 \CACHE_MEM_reg[3][157]  ( .D(n11013), .CK(N28803), .Q(n3306), .QN(
        n7573) );
  DFF_X1 \CACHE_MEM_reg[3][156]  ( .D(n11012), .CK(N28803), .Q(n3293), .QN(
        n7589) );
  DFF_X1 \CACHE_MEM_reg[3][155]  ( .D(n11011), .CK(N28803), .Q(n3282), .QN(
        n7605) );
  DFF_X1 \CACHE_MEM_reg[3][154]  ( .D(n11010), .CK(N28803), .Q(n3260), .QN(
        n7621) );
  DFF_X1 \CACHE_MEM_reg[3][153]  ( .D(n11009), .CK(N28803), .Q(n3249), .QN(
        n7637) );
  DFF_X1 \CACHE_MEM_reg[3][152]  ( .D(n11008), .CK(N28803), .Q(n3232), .QN(
        n7653) );
  DFF_X1 \CACHE_MEM_reg[3][151]  ( .D(n11007), .CK(N28803), .Q(n3221), .QN(
        n7669) );
  DFF_X1 \CACHE_MEM_reg[3][150]  ( .D(n11006), .CK(N28803), .Q(n3208), .QN(
        n7685) );
  DFF_X1 \CACHE_MEM_reg[3][149]  ( .D(n11005), .CK(N28803), .Q(n3193), .QN(
        n7701) );
  DFF_X1 \CACHE_MEM_reg[3][148]  ( .D(n11004), .CK(N28803), .Q(n3180), .QN(
        n7717) );
  DFF_X1 \CACHE_MEM_reg[3][147]  ( .D(n11003), .CK(N28803), .Q(n3169), .QN(
        n7733) );
  DFF_X1 \CACHE_MEM_reg[3][146]  ( .D(n11002), .CK(N28803), .Q(n3152), .QN(
        n7749) );
  DFF_X1 \CACHE_MEM_reg[3][145]  ( .D(n11001), .CK(N28803), .Q(n3141), .QN(
        n7765) );
  DFF_X1 \CACHE_MEM_reg[3][144]  ( .D(n11000), .CK(N28803), .Q(n3119), .QN(
        n7781) );
  DFF_X1 \CACHE_MEM_reg[3][143]  ( .D(n10999), .CK(N28803), .Q(n3108), .QN(
        n7797) );
  DFF_X1 \CACHE_MEM_reg[3][142]  ( .D(n10998), .CK(N28803), .Q(n3095), .QN(
        n7813) );
  DFF_X1 \CACHE_MEM_reg[3][141]  ( .D(n10997), .CK(N28803), .Q(n3080), .QN(
        n7829) );
  DFF_X1 \CACHE_MEM_reg[3][140]  ( .D(n10996), .CK(N28803), .Q(n3067), .QN(
        n7845) );
  DFF_X1 \CACHE_MEM_reg[3][139]  ( .D(n10995), .CK(N28803), .Q(n3056), .QN(
        n7861) );
  DFF_X1 \CACHE_MEM_reg[3][138]  ( .D(n10994), .CK(N28803), .Q(n3039), .QN(
        n7877) );
  DFF_X1 \CACHE_MEM_reg[3][137]  ( .D(n10993), .CK(N28803), .Q(n3028), .QN(
        n7893) );
  DFF_X1 \CACHE_MEM_reg[3][136]  ( .D(n10992), .CK(N28803), .Q(n3011), .QN(
        n7909) );
  DFF_X1 \CACHE_MEM_reg[3][135]  ( .D(n10991), .CK(N28803), .Q(n3000), .QN(
        n7925) );
  DFF_X1 \CACHE_MEM_reg[3][134]  ( .D(n10990), .CK(N28803), .Q(n2987), .QN(
        n7941) );
  DFF_X1 \CACHE_MEM_reg[3][133]  ( .D(n10989), .CK(N28803), .Q(n2967), .QN(
        n7957) );
  DFF_X1 \CACHE_MEM_reg[3][132]  ( .D(n10988), .CK(N28803), .Q(n2954), .QN(
        n7973) );
  DFF_X1 \CACHE_MEM_reg[3][131]  ( .D(n10987), .CK(N28803), .Q(n2943), .QN(
        n7989) );
  DFF_X1 \CACHE_MEM_reg[3][130]  ( .D(n10986), .CK(N28803), .Q(n2926), .QN(
        n8005) );
  DFF_X1 \CACHE_MEM_reg[3][129]  ( .D(n10985), .CK(N28803), .Q(n2915), .QN(
        n8021) );
  DFF_X1 \CACHE_MEM_reg[3][128]  ( .D(n10984), .CK(N28803), .Q(n2898), .QN(
        n8037) );
  DFF_X1 \CACHE_MEM_reg[3][127]  ( .D(n10983), .CK(N28803), .Q(n1993), .QN(
        n8053) );
  DFF_X1 \CACHE_MEM_reg[3][126]  ( .D(n10982), .CK(N28803), .Q(n1980), .QN(
        n8069) );
  DFF_X1 \CACHE_MEM_reg[3][125]  ( .D(n10981), .CK(N28803), .Q(n1960), .QN(
        n8085) );
  DFF_X1 \CACHE_MEM_reg[3][124]  ( .D(n10980), .CK(N28803), .Q(n1944), .QN(
        n8101) );
  DFF_X1 \CACHE_MEM_reg[3][123]  ( .D(n10979), .CK(N28803), .Q(n1919), .QN(
        n8117) );
  DFF_X1 \CACHE_MEM_reg[3][122]  ( .D(n10978), .CK(N28803), .Q(n1903), .QN(
        n8133) );
  DFF_X1 \CACHE_MEM_reg[3][121]  ( .D(n10977), .CK(N28803), .Q(n1883), .QN(
        n8149) );
  DFF_X1 \CACHE_MEM_reg[3][120]  ( .D(n10976), .CK(N28803), .Q(n1867), .QN(
        n8165) );
  DFF_X1 \CACHE_MEM_reg[3][119]  ( .D(n10975), .CK(N28803), .Q(n1847), .QN(
        n8181) );
  DFF_X1 \CACHE_MEM_reg[3][118]  ( .D(n10974), .CK(N28803), .Q(n1831), .QN(
        n8197) );
  DFF_X1 \CACHE_MEM_reg[3][117]  ( .D(n10973), .CK(N28803), .Q(n1811), .QN(
        n8213) );
  DFF_X1 \CACHE_MEM_reg[3][116]  ( .D(n10972), .CK(N28803), .Q(n1795), .QN(
        n8229) );
  DFF_X1 \CACHE_MEM_reg[3][115]  ( .D(n10971), .CK(N28803), .Q(n1770), .QN(
        n8245) );
  DFF_X1 \CACHE_MEM_reg[3][114]  ( .D(n10970), .CK(N28803), .Q(n1754), .QN(
        n8261) );
  DFF_X1 \CACHE_MEM_reg[3][113]  ( .D(n10969), .CK(N28803), .Q(n1734), .QN(
        n8277) );
  DFF_X1 \CACHE_MEM_reg[3][112]  ( .D(n10968), .CK(N28803), .Q(n1718), .QN(
        n8293) );
  DFF_X1 \CACHE_MEM_reg[3][111]  ( .D(n10967), .CK(N28803), .Q(n1698), .QN(
        n8309) );
  DFF_X1 \CACHE_MEM_reg[3][110]  ( .D(n10966), .CK(N28803), .Q(n1682), .QN(
        n8325) );
  DFF_X1 \CACHE_MEM_reg[3][109]  ( .D(n10965), .CK(N28803), .Q(n1662), .QN(
        n8341) );
  DFF_X1 \CACHE_MEM_reg[3][108]  ( .D(n10964), .CK(N28803), .Q(n1646), .QN(
        n8357) );
  DFF_X1 \CACHE_MEM_reg[3][107]  ( .D(n10963), .CK(N28803), .Q(n1621), .QN(
        n8373) );
  DFF_X1 \CACHE_MEM_reg[3][106]  ( .D(n10962), .CK(N28803), .Q(n1605), .QN(
        n8389) );
  DFF_X1 \CACHE_MEM_reg[3][105]  ( .D(n10961), .CK(N28803), .Q(n1585), .QN(
        n8405) );
  DFF_X1 \CACHE_MEM_reg[3][104]  ( .D(n10960), .CK(N28803), .Q(n1569), .QN(
        n8421) );
  DFF_X1 \CACHE_MEM_reg[3][103]  ( .D(n10959), .CK(N28803), .Q(n1549), .QN(
        n8437) );
  DFF_X1 \CACHE_MEM_reg[3][102]  ( .D(n10958), .CK(N28803), .Q(n1533), .QN(
        n8453) );
  DFF_X1 \CACHE_MEM_reg[3][101]  ( .D(n10957), .CK(N28803), .Q(n1513), .QN(
        n8469) );
  DFF_X1 \CACHE_MEM_reg[3][100]  ( .D(n10956), .CK(N28803), .Q(n1497), .QN(
        n8485) );
  DFF_X1 \CACHE_MEM_reg[3][99]  ( .D(n10955), .CK(N28803), .Q(n1472), .QN(
        n8501) );
  DFF_X1 \CACHE_MEM_reg[3][98]  ( .D(n10954), .CK(N28803), .Q(n1456), .QN(
        n8517) );
  DFF_X1 \CACHE_MEM_reg[3][97]  ( .D(n10953), .CK(N28803), .Q(n1436), .QN(
        n8533) );
  DFF_X1 \CACHE_MEM_reg[3][96]  ( .D(n10952), .CK(N28803), .Q(n1420), .QN(
        n8549) );
  DFF_X1 \CACHE_MEM_reg[3][95]  ( .D(n10951), .CK(N28803), .Q(n1996), .QN(
        n8565) );
  DFF_X1 \CACHE_MEM_reg[3][94]  ( .D(n10950), .CK(N28803), .Q(n1985), .QN(
        n8581) );
  DFF_X1 \CACHE_MEM_reg[3][93]  ( .D(n10949), .CK(N28803), .Q(n1965), .QN(
        n8597) );
  DFF_X1 \CACHE_MEM_reg[3][92]  ( .D(n10948), .CK(N28803), .Q(n1949), .QN(
        n8613) );
  DFF_X1 \CACHE_MEM_reg[3][91]  ( .D(n10947), .CK(N28803), .Q(n1924), .QN(
        n8629) );
  DFF_X1 \CACHE_MEM_reg[3][90]  ( .D(n10946), .CK(N28803), .Q(n1908), .QN(
        n8645) );
  DFF_X1 \CACHE_MEM_reg[3][89]  ( .D(n10945), .CK(N28803), .Q(n1888), .QN(
        n8661) );
  DFF_X1 \CACHE_MEM_reg[3][88]  ( .D(n10944), .CK(N28803), .Q(n1872), .QN(
        n8677) );
  DFF_X1 \CACHE_MEM_reg[3][87]  ( .D(n10943), .CK(N28803), .Q(n1852), .QN(
        n8693) );
  DFF_X1 \CACHE_MEM_reg[3][86]  ( .D(n10942), .CK(N28803), .Q(n1836), .QN(
        n8709) );
  DFF_X1 \CACHE_MEM_reg[3][85]  ( .D(n10941), .CK(N28803), .Q(n1816), .QN(
        n8725) );
  DFF_X1 \CACHE_MEM_reg[3][84]  ( .D(n10940), .CK(N28803), .Q(n1800), .QN(
        n8741) );
  DFF_X1 \CACHE_MEM_reg[3][83]  ( .D(n10939), .CK(N28803), .Q(n1775), .QN(
        n8757) );
  DFF_X1 \CACHE_MEM_reg[3][82]  ( .D(n10938), .CK(N28803), .Q(n1759), .QN(
        n8773) );
  DFF_X1 \CACHE_MEM_reg[3][81]  ( .D(n10937), .CK(N28803), .Q(n1739), .QN(
        n8789) );
  DFF_X1 \CACHE_MEM_reg[3][80]  ( .D(n10936), .CK(N28803), .Q(n1723), .QN(
        n8805) );
  DFF_X1 \CACHE_MEM_reg[3][79]  ( .D(n10935), .CK(N28803), .Q(n1703), .QN(
        n8821) );
  DFF_X1 \CACHE_MEM_reg[3][78]  ( .D(n10934), .CK(N28803), .Q(n1687), .QN(
        n8837) );
  DFF_X1 \CACHE_MEM_reg[3][77]  ( .D(n10933), .CK(N28803), .Q(n1667), .QN(
        n8853) );
  DFF_X1 \CACHE_MEM_reg[3][76]  ( .D(n10932), .CK(N28803), .Q(n1651), .QN(
        n8869) );
  DFF_X1 \CACHE_MEM_reg[3][75]  ( .D(n10931), .CK(N28803), .Q(n1626), .QN(
        n8885) );
  DFF_X1 \CACHE_MEM_reg[3][74]  ( .D(n10930), .CK(N28803), .Q(n1610), .QN(
        n8901) );
  DFF_X1 \CACHE_MEM_reg[3][73]  ( .D(n10929), .CK(N28803), .Q(n1590), .QN(
        n8917) );
  DFF_X1 \CACHE_MEM_reg[3][72]  ( .D(n10928), .CK(N28803), .Q(n1574), .QN(
        n8933) );
  DFF_X1 \CACHE_MEM_reg[3][71]  ( .D(n10927), .CK(N28803), .Q(n1554), .QN(
        n8949) );
  DFF_X1 \CACHE_MEM_reg[3][70]  ( .D(n10926), .CK(N28803), .Q(n1538), .QN(
        n8965) );
  DFF_X1 \CACHE_MEM_reg[3][69]  ( .D(n10925), .CK(N28803), .Q(n1518), .QN(
        n8981) );
  DFF_X1 \CACHE_MEM_reg[3][68]  ( .D(n10924), .CK(N28803), .Q(n1502), .QN(
        n8997) );
  DFF_X1 \CACHE_MEM_reg[3][67]  ( .D(n10923), .CK(N28803), .Q(n1477), .QN(
        n9013) );
  DFF_X1 \CACHE_MEM_reg[3][66]  ( .D(n10922), .CK(N28803), .Q(n1461), .QN(
        n9029) );
  DFF_X1 \CACHE_MEM_reg[3][65]  ( .D(n10921), .CK(N28803), .Q(n1441), .QN(
        n9045) );
  DFF_X1 \CACHE_MEM_reg[3][64]  ( .D(n10920), .CK(N28803), .Q(n1425), .QN(
        n9061) );
  DFF_X1 \CACHE_MEM_reg[3][63]  ( .D(n10919), .CK(N28803), .Q(n2440), .QN(
        n9077) );
  DFF_X1 \CACHE_MEM_reg[3][62]  ( .D(n10918), .CK(N28803), .Q(n2427), .QN(
        n9093) );
  DFF_X1 \CACHE_MEM_reg[3][61]  ( .D(n10917), .CK(N28803), .Q(n2412), .QN(
        n9109) );
  DFF_X1 \CACHE_MEM_reg[3][60]  ( .D(n10916), .CK(N28803), .Q(n2399), .QN(
        n9125) );
  DFF_X1 \CACHE_MEM_reg[3][59]  ( .D(n10915), .CK(N28803), .Q(n2388), .QN(
        n9141) );
  DFF_X1 \CACHE_MEM_reg[3][58]  ( .D(n10914), .CK(N28803), .Q(n2366), .QN(
        n9157) );
  DFF_X1 \CACHE_MEM_reg[3][57]  ( .D(n10913), .CK(N28803), .Q(n2355), .QN(
        n9173) );
  DFF_X1 \CACHE_MEM_reg[3][56]  ( .D(n10912), .CK(N28803), .Q(n2338), .QN(
        n9189) );
  DFF_X1 \CACHE_MEM_reg[3][55]  ( .D(n10911), .CK(N28803), .Q(n2327), .QN(
        n9205) );
  DFF_X1 \CACHE_MEM_reg[3][54]  ( .D(n10910), .CK(N28803), .Q(n2314), .QN(
        n9221) );
  DFF_X1 \CACHE_MEM_reg[3][53]  ( .D(n10909), .CK(N28803), .Q(n2299), .QN(
        n9237) );
  DFF_X1 \CACHE_MEM_reg[3][52]  ( .D(n10908), .CK(N28803), .Q(n2286), .QN(
        n9253) );
  DFF_X1 \CACHE_MEM_reg[3][51]  ( .D(n10907), .CK(N28803), .Q(n2275), .QN(
        n9269) );
  DFF_X1 \CACHE_MEM_reg[3][50]  ( .D(n10906), .CK(N28803), .Q(n2258), .QN(
        n9285) );
  DFF_X1 \CACHE_MEM_reg[3][49]  ( .D(n10905), .CK(N28803), .Q(n2247), .QN(
        n9301) );
  DFF_X1 \CACHE_MEM_reg[3][48]  ( .D(n10904), .CK(N28803), .Q(n2225), .QN(
        n9317) );
  DFF_X1 \CACHE_MEM_reg[3][47]  ( .D(n10903), .CK(N28803), .Q(n2214), .QN(
        n9333) );
  DFF_X1 \CACHE_MEM_reg[3][46]  ( .D(n10902), .CK(N28803), .Q(n2201), .QN(
        n9349) );
  DFF_X1 \CACHE_MEM_reg[3][45]  ( .D(n10901), .CK(N28803), .Q(n2186), .QN(
        n9365) );
  DFF_X1 \CACHE_MEM_reg[3][44]  ( .D(n10900), .CK(N28803), .Q(n2173), .QN(
        n9381) );
  DFF_X1 \CACHE_MEM_reg[3][43]  ( .D(n10899), .CK(N28803), .Q(n2162), .QN(
        n9397) );
  DFF_X1 \CACHE_MEM_reg[3][42]  ( .D(n10898), .CK(N28803), .Q(n2145), .QN(
        n9413) );
  DFF_X1 \CACHE_MEM_reg[3][41]  ( .D(n10897), .CK(N28803), .Q(n2134), .QN(
        n9429) );
  DFF_X1 \CACHE_MEM_reg[3][40]  ( .D(n10896), .CK(N28803), .Q(n2117), .QN(
        n9445) );
  DFF_X1 \CACHE_MEM_reg[3][39]  ( .D(n10895), .CK(N28803), .Q(n2106), .QN(
        n9461) );
  DFF_X1 \CACHE_MEM_reg[3][38]  ( .D(n10894), .CK(N28803), .Q(n2093), .QN(
        n9477) );
  DFF_X1 \CACHE_MEM_reg[3][37]  ( .D(n10893), .CK(N28803), .Q(n2073), .QN(
        n9493) );
  DFF_X1 \CACHE_MEM_reg[3][36]  ( .D(n10892), .CK(N28803), .Q(n2060), .QN(
        n9509) );
  DFF_X1 \CACHE_MEM_reg[3][35]  ( .D(n10891), .CK(N28803), .Q(n2049), .QN(
        n9525) );
  DFF_X1 \CACHE_MEM_reg[3][34]  ( .D(n10890), .CK(N28803), .Q(n2032), .QN(
        n9541) );
  DFF_X1 \CACHE_MEM_reg[3][33]  ( .D(n10889), .CK(N28803), .Q(n2021), .QN(
        n9557) );
  DFF_X1 \CACHE_MEM_reg[3][32]  ( .D(n10888), .CK(N28803), .Q(n2004), .QN(
        n9573) );
  DFF_X1 \CACHE_MEM_reg[3][31]  ( .D(n10887), .CK(N28803), .Q(n2443), .QN(
        n9589) );
  DFF_X1 \CACHE_MEM_reg[3][30]  ( .D(n10886), .CK(N28803), .Q(n2432), .QN(
        n9605) );
  DFF_X1 \CACHE_MEM_reg[3][29]  ( .D(n10885), .CK(N28803), .Q(n2415), .QN(
        n9621) );
  DFF_X1 \CACHE_MEM_reg[3][28]  ( .D(n10884), .CK(N28803), .Q(n2404), .QN(
        n9637) );
  DFF_X1 \CACHE_MEM_reg[3][27]  ( .D(n10883), .CK(N28803), .Q(n2391), .QN(
        n9653) );
  DFF_X1 \CACHE_MEM_reg[3][26]  ( .D(n10882), .CK(N28803), .Q(n2371), .QN(
        n9669) );
  DFF_X1 \CACHE_MEM_reg[3][25]  ( .D(n10881), .CK(N28803), .Q(n2358), .QN(
        n9685) );
  DFF_X1 \CACHE_MEM_reg[3][24]  ( .D(n10880), .CK(N28803), .Q(n2347), .QN(
        n9701) );
  DFF_X1 \CACHE_MEM_reg[3][23]  ( .D(n10879), .CK(N28803), .Q(n2330), .QN(
        n9717) );
  DFF_X1 \CACHE_MEM_reg[3][22]  ( .D(n10878), .CK(N28803), .Q(n2319), .QN(
        n9733) );
  DFF_X1 \CACHE_MEM_reg[3][21]  ( .D(n10877), .CK(N28803), .Q(n2302), .QN(
        n9749) );
  DFF_X1 \CACHE_MEM_reg[3][20]  ( .D(n10876), .CK(N28803), .Q(n2291), .QN(
        n9765) );
  DFF_X1 \CACHE_MEM_reg[3][19]  ( .D(n10875), .CK(N28803), .Q(n2278), .QN(
        n9781) );
  DFF_X1 \CACHE_MEM_reg[3][18]  ( .D(n10874), .CK(N28803), .Q(n2263), .QN(
        n9797) );
  DFF_X1 \CACHE_MEM_reg[3][17]  ( .D(n10873), .CK(N28803), .Q(n2250), .QN(
        n9813) );
  DFF_X1 \CACHE_MEM_reg[3][16]  ( .D(n10872), .CK(N28803), .Q(n2239), .QN(
        n9829) );
  DFF_X1 \CACHE_MEM_reg[3][15]  ( .D(n10871), .CK(N28803), .Q(n2217), .QN(
        n9845) );
  DFF_X1 \CACHE_MEM_reg[3][14]  ( .D(n10870), .CK(N28803), .Q(n2206), .QN(
        n9861) );
  DFF_X1 \CACHE_MEM_reg[3][13]  ( .D(n10869), .CK(N28803), .Q(n2189), .QN(
        n9877) );
  DFF_X1 \CACHE_MEM_reg[3][12]  ( .D(n10868), .CK(N28803), .Q(n2178), .QN(
        n9893) );
  DFF_X1 \CACHE_MEM_reg[3][11]  ( .D(n10867), .CK(N28803), .Q(n2165), .QN(
        n9909) );
  DFF_X1 \CACHE_MEM_reg[3][10]  ( .D(n10866), .CK(N28803), .Q(n2150), .QN(
        n9925) );
  DFF_X1 \CACHE_MEM_reg[3][9]  ( .D(n10865), .CK(N28803), .Q(n2137), .QN(n9941) );
  DFF_X1 \CACHE_MEM_reg[3][8]  ( .D(n10864), .CK(N28803), .Q(n2126), .QN(n9957) );
  DFF_X1 \CACHE_MEM_reg[3][7]  ( .D(n10863), .CK(N28803), .Q(n2109), .QN(n9973) );
  DFF_X1 \CACHE_MEM_reg[3][6]  ( .D(n10862), .CK(N28803), .Q(n2098), .QN(n9989) );
  DFF_X1 \CACHE_MEM_reg[3][5]  ( .D(n10861), .CK(N28803), .Q(n2076), .QN(
        n10005) );
  DFF_X1 \CACHE_MEM_reg[3][4]  ( .D(n10860), .CK(N28803), .Q(n2065), .QN(
        n10021) );
  DFF_X1 \CACHE_MEM_reg[3][3]  ( .D(n10859), .CK(N28803), .Q(n2052), .QN(
        n10037) );
  DFF_X1 \CACHE_MEM_reg[3][2]  ( .D(n10858), .CK(N28803), .Q(n2037), .QN(
        n10053) );
  DFF_X1 \CACHE_MEM_reg[3][1]  ( .D(n10857), .CK(N28803), .Q(n2024), .QN(
        n10069) );
  DFF_X1 \CACHE_MEM_reg[3][0]  ( .D(n10856), .CK(N28803), .Q(n2013), .QN(
        n10085) );
  DFF_X1 \CACHE_MEM_reg[2][255]  ( .D(n10855), .CK(N28803), .QN(n6001) );
  DFF_X1 \CACHE_MEM_reg[2][254]  ( .D(n10854), .CK(N28803), .QN(n6017) );
  DFF_X1 \CACHE_MEM_reg[2][253]  ( .D(n10853), .CK(N28803), .QN(n6033) );
  DFF_X1 \CACHE_MEM_reg[2][252]  ( .D(n10852), .CK(N28803), .QN(n6049) );
  DFF_X1 \CACHE_MEM_reg[2][251]  ( .D(n10851), .CK(N28803), .QN(n6065) );
  DFF_X1 \CACHE_MEM_reg[2][250]  ( .D(n10850), .CK(N28803), .QN(n6081) );
  DFF_X1 \CACHE_MEM_reg[2][249]  ( .D(n10849), .CK(N28803), .QN(n6097) );
  DFF_X1 \CACHE_MEM_reg[2][248]  ( .D(n10848), .CK(N28803), .QN(n6113) );
  DFF_X1 \CACHE_MEM_reg[2][247]  ( .D(n10847), .CK(N28803), .QN(n6129) );
  DFF_X1 \CACHE_MEM_reg[2][246]  ( .D(n10846), .CK(N28803), .QN(n6145) );
  DFF_X1 \CACHE_MEM_reg[2][245]  ( .D(n10845), .CK(N28803), .QN(n6161) );
  DFF_X1 \CACHE_MEM_reg[2][244]  ( .D(n10844), .CK(N28803), .QN(n6177) );
  DFF_X1 \CACHE_MEM_reg[2][243]  ( .D(n10843), .CK(N28803), .QN(n6193) );
  DFF_X1 \CACHE_MEM_reg[2][242]  ( .D(n10842), .CK(N28803), .QN(n6209) );
  DFF_X1 \CACHE_MEM_reg[2][241]  ( .D(n10841), .CK(N28803), .QN(n6225) );
  DFF_X1 \CACHE_MEM_reg[2][240]  ( .D(n10840), .CK(N28803), .QN(n6241) );
  DFF_X1 \CACHE_MEM_reg[2][239]  ( .D(n10839), .CK(N28803), .QN(n6257) );
  DFF_X1 \CACHE_MEM_reg[2][238]  ( .D(n10838), .CK(N28803), .QN(n6273) );
  DFF_X1 \CACHE_MEM_reg[2][237]  ( .D(n10837), .CK(N28803), .QN(n6289) );
  DFF_X1 \CACHE_MEM_reg[2][236]  ( .D(n10836), .CK(N28803), .QN(n6305) );
  DFF_X1 \CACHE_MEM_reg[2][235]  ( .D(n10835), .CK(N28803), .QN(n6321) );
  DFF_X1 \CACHE_MEM_reg[2][234]  ( .D(n10834), .CK(N28803), .QN(n6337) );
  DFF_X1 \CACHE_MEM_reg[2][233]  ( .D(n10833), .CK(N28803), .QN(n6353) );
  DFF_X1 \CACHE_MEM_reg[2][232]  ( .D(n10832), .CK(N28803), .QN(n6369) );
  DFF_X1 \CACHE_MEM_reg[2][231]  ( .D(n10831), .CK(N28803), .QN(n6385) );
  DFF_X1 \CACHE_MEM_reg[2][230]  ( .D(n10830), .CK(N28803), .QN(n6401) );
  DFF_X1 \CACHE_MEM_reg[2][229]  ( .D(n10829), .CK(N28803), .QN(n6417) );
  DFF_X1 \CACHE_MEM_reg[2][228]  ( .D(n10828), .CK(N28803), .QN(n6433) );
  DFF_X1 \CACHE_MEM_reg[2][227]  ( .D(n10827), .CK(N28803), .QN(n6449) );
  DFF_X1 \CACHE_MEM_reg[2][226]  ( .D(n10826), .CK(N28803), .QN(n6465) );
  DFF_X1 \CACHE_MEM_reg[2][225]  ( .D(n10825), .CK(N28803), .QN(n6481) );
  DFF_X1 \CACHE_MEM_reg[2][224]  ( .D(n10824), .CK(N28803), .QN(n6497) );
  DFF_X1 \CACHE_MEM_reg[2][223]  ( .D(n10823), .CK(N28803), .QN(n6513) );
  DFF_X1 \CACHE_MEM_reg[2][222]  ( .D(n10822), .CK(N28803), .QN(n6529) );
  DFF_X1 \CACHE_MEM_reg[2][221]  ( .D(n10821), .CK(N28803), .QN(n6545) );
  DFF_X1 \CACHE_MEM_reg[2][220]  ( .D(n10820), .CK(N28803), .QN(n6561) );
  DFF_X1 \CACHE_MEM_reg[2][219]  ( .D(n10819), .CK(N28803), .QN(n6577) );
  DFF_X1 \CACHE_MEM_reg[2][218]  ( .D(n10818), .CK(N28803), .QN(n6593) );
  DFF_X1 \CACHE_MEM_reg[2][217]  ( .D(n10817), .CK(N28803), .QN(n6609) );
  DFF_X1 \CACHE_MEM_reg[2][216]  ( .D(n10816), .CK(N28803), .QN(n6625) );
  DFF_X1 \CACHE_MEM_reg[2][215]  ( .D(n10815), .CK(N28803), .QN(n6641) );
  DFF_X1 \CACHE_MEM_reg[2][214]  ( .D(n10814), .CK(N28803), .QN(n6657) );
  DFF_X1 \CACHE_MEM_reg[2][213]  ( .D(n10813), .CK(N28803), .QN(n6673) );
  DFF_X1 \CACHE_MEM_reg[2][212]  ( .D(n10812), .CK(N28803), .QN(n6689) );
  DFF_X1 \CACHE_MEM_reg[2][211]  ( .D(n10811), .CK(N28803), .QN(n6705) );
  DFF_X1 \CACHE_MEM_reg[2][210]  ( .D(n10810), .CK(N28803), .QN(n6721) );
  DFF_X1 \CACHE_MEM_reg[2][209]  ( .D(n10809), .CK(N28803), .QN(n6737) );
  DFF_X1 \CACHE_MEM_reg[2][208]  ( .D(n10808), .CK(N28803), .QN(n6753) );
  DFF_X1 \CACHE_MEM_reg[2][207]  ( .D(n10807), .CK(N28803), .QN(n6769) );
  DFF_X1 \CACHE_MEM_reg[2][206]  ( .D(n10806), .CK(N28803), .QN(n6785) );
  DFF_X1 \CACHE_MEM_reg[2][205]  ( .D(n10805), .CK(N28803), .QN(n6801) );
  DFF_X1 \CACHE_MEM_reg[2][204]  ( .D(n10804), .CK(N28803), .QN(n6817) );
  DFF_X1 \CACHE_MEM_reg[2][203]  ( .D(n10803), .CK(N28803), .QN(n6833) );
  DFF_X1 \CACHE_MEM_reg[2][202]  ( .D(n10802), .CK(N28803), .QN(n6849) );
  DFF_X1 \CACHE_MEM_reg[2][201]  ( .D(n10801), .CK(N28803), .QN(n6865) );
  DFF_X1 \CACHE_MEM_reg[2][200]  ( .D(n10800), .CK(N28803), .QN(n6881) );
  DFF_X1 \CACHE_MEM_reg[2][199]  ( .D(n10799), .CK(N28803), .QN(n6897) );
  DFF_X1 \CACHE_MEM_reg[2][198]  ( .D(n10798), .CK(N28803), .QN(n6913) );
  DFF_X1 \CACHE_MEM_reg[2][197]  ( .D(n10797), .CK(N28803), .QN(n6929) );
  DFF_X1 \CACHE_MEM_reg[2][196]  ( .D(n10796), .CK(N28803), .QN(n6945) );
  DFF_X1 \CACHE_MEM_reg[2][195]  ( .D(n10795), .CK(N28803), .QN(n6961) );
  DFF_X1 \CACHE_MEM_reg[2][194]  ( .D(n10794), .CK(N28803), .QN(n6977) );
  DFF_X1 \CACHE_MEM_reg[2][193]  ( .D(n10793), .CK(N28803), .QN(n6993) );
  DFF_X1 \CACHE_MEM_reg[2][192]  ( .D(n10792), .CK(N28803), .QN(n7009) );
  DFF_X1 \CACHE_MEM_reg[2][191]  ( .D(n10791), .CK(N28803), .QN(n7025) );
  DFF_X1 \CACHE_MEM_reg[2][190]  ( .D(n10790), .CK(N28803), .QN(n7041) );
  DFF_X1 \CACHE_MEM_reg[2][189]  ( .D(n10789), .CK(N28803), .QN(n7057) );
  DFF_X1 \CACHE_MEM_reg[2][188]  ( .D(n10788), .CK(N28803), .QN(n7073) );
  DFF_X1 \CACHE_MEM_reg[2][187]  ( .D(n10787), .CK(N28803), .QN(n7089) );
  DFF_X1 \CACHE_MEM_reg[2][186]  ( .D(n10786), .CK(N28803), .QN(n7105) );
  DFF_X1 \CACHE_MEM_reg[2][185]  ( .D(n10785), .CK(N28803), .QN(n7121) );
  DFF_X1 \CACHE_MEM_reg[2][184]  ( .D(n10784), .CK(N28803), .QN(n7137) );
  DFF_X1 \CACHE_MEM_reg[2][183]  ( .D(n10783), .CK(N28803), .QN(n7153) );
  DFF_X1 \CACHE_MEM_reg[2][182]  ( .D(n10782), .CK(N28803), .QN(n7169) );
  DFF_X1 \CACHE_MEM_reg[2][181]  ( .D(n10781), .CK(N28803), .QN(n7185) );
  DFF_X1 \CACHE_MEM_reg[2][180]  ( .D(n10780), .CK(N28803), .QN(n7201) );
  DFF_X1 \CACHE_MEM_reg[2][179]  ( .D(n10779), .CK(N28803), .QN(n7217) );
  DFF_X1 \CACHE_MEM_reg[2][178]  ( .D(n10778), .CK(N28803), .QN(n7233) );
  DFF_X1 \CACHE_MEM_reg[2][177]  ( .D(n10777), .CK(N28803), .QN(n7249) );
  DFF_X1 \CACHE_MEM_reg[2][176]  ( .D(n10776), .CK(N28803), .QN(n7265) );
  DFF_X1 \CACHE_MEM_reg[2][175]  ( .D(n10775), .CK(N28803), .QN(n7281) );
  DFF_X1 \CACHE_MEM_reg[2][174]  ( .D(n10774), .CK(N28803), .QN(n7297) );
  DFF_X1 \CACHE_MEM_reg[2][173]  ( .D(n10773), .CK(N28803), .QN(n7313) );
  DFF_X1 \CACHE_MEM_reg[2][172]  ( .D(n10772), .CK(N28803), .QN(n7329) );
  DFF_X1 \CACHE_MEM_reg[2][171]  ( .D(n10771), .CK(N28803), .QN(n7345) );
  DFF_X1 \CACHE_MEM_reg[2][170]  ( .D(n10770), .CK(N28803), .QN(n7361) );
  DFF_X1 \CACHE_MEM_reg[2][169]  ( .D(n10769), .CK(N28803), .QN(n7377) );
  DFF_X1 \CACHE_MEM_reg[2][168]  ( .D(n10768), .CK(N28803), .QN(n7393) );
  DFF_X1 \CACHE_MEM_reg[2][167]  ( .D(n10767), .CK(N28803), .QN(n7409) );
  DFF_X1 \CACHE_MEM_reg[2][166]  ( .D(n10766), .CK(N28803), .QN(n7425) );
  DFF_X1 \CACHE_MEM_reg[2][165]  ( .D(n10765), .CK(N28803), .QN(n7441) );
  DFF_X1 \CACHE_MEM_reg[2][164]  ( .D(n10764), .CK(N28803), .QN(n7457) );
  DFF_X1 \CACHE_MEM_reg[2][163]  ( .D(n10763), .CK(N28803), .QN(n7473) );
  DFF_X1 \CACHE_MEM_reg[2][162]  ( .D(n10762), .CK(N28803), .QN(n7489) );
  DFF_X1 \CACHE_MEM_reg[2][161]  ( .D(n10761), .CK(N28803), .QN(n7505) );
  DFF_X1 \CACHE_MEM_reg[2][160]  ( .D(n10760), .CK(N28803), .QN(n7521) );
  DFF_X1 \CACHE_MEM_reg[2][159]  ( .D(n10759), .CK(N28803), .QN(n7537) );
  DFF_X1 \CACHE_MEM_reg[2][158]  ( .D(n10758), .CK(N28803), .QN(n7553) );
  DFF_X1 \CACHE_MEM_reg[2][157]  ( .D(n10757), .CK(N28803), .QN(n7569) );
  DFF_X1 \CACHE_MEM_reg[2][156]  ( .D(n10756), .CK(N28803), .QN(n7585) );
  DFF_X1 \CACHE_MEM_reg[2][155]  ( .D(n10755), .CK(N28803), .QN(n7601) );
  DFF_X1 \CACHE_MEM_reg[2][154]  ( .D(n10754), .CK(N28803), .QN(n7617) );
  DFF_X1 \CACHE_MEM_reg[2][153]  ( .D(n10753), .CK(N28803), .QN(n7633) );
  DFF_X1 \CACHE_MEM_reg[2][152]  ( .D(n10752), .CK(N28803), .QN(n7649) );
  DFF_X1 \CACHE_MEM_reg[2][151]  ( .D(n10751), .CK(N28803), .QN(n7665) );
  DFF_X1 \CACHE_MEM_reg[2][150]  ( .D(n10750), .CK(N28803), .QN(n7681) );
  DFF_X1 \CACHE_MEM_reg[2][149]  ( .D(n10749), .CK(N28803), .QN(n7697) );
  DFF_X1 \CACHE_MEM_reg[2][148]  ( .D(n10748), .CK(N28803), .QN(n7713) );
  DFF_X1 \CACHE_MEM_reg[2][147]  ( .D(n10747), .CK(N28803), .QN(n7729) );
  DFF_X1 \CACHE_MEM_reg[2][146]  ( .D(n10746), .CK(N28803), .QN(n7745) );
  DFF_X1 \CACHE_MEM_reg[2][145]  ( .D(n10745), .CK(N28803), .QN(n7761) );
  DFF_X1 \CACHE_MEM_reg[2][144]  ( .D(n10744), .CK(N28803), .QN(n7777) );
  DFF_X1 \CACHE_MEM_reg[2][143]  ( .D(n10743), .CK(N28803), .QN(n7793) );
  DFF_X1 \CACHE_MEM_reg[2][142]  ( .D(n10742), .CK(N28803), .QN(n7809) );
  DFF_X1 \CACHE_MEM_reg[2][141]  ( .D(n10741), .CK(N28803), .QN(n7825) );
  DFF_X1 \CACHE_MEM_reg[2][140]  ( .D(n10740), .CK(N28803), .QN(n7841) );
  DFF_X1 \CACHE_MEM_reg[2][139]  ( .D(n10739), .CK(N28803), .QN(n7857) );
  DFF_X1 \CACHE_MEM_reg[2][138]  ( .D(n10738), .CK(N28803), .QN(n7873) );
  DFF_X1 \CACHE_MEM_reg[2][137]  ( .D(n10737), .CK(N28803), .QN(n7889) );
  DFF_X1 \CACHE_MEM_reg[2][136]  ( .D(n10736), .CK(N28803), .QN(n7905) );
  DFF_X1 \CACHE_MEM_reg[2][135]  ( .D(n10735), .CK(N28803), .QN(n7921) );
  DFF_X1 \CACHE_MEM_reg[2][134]  ( .D(n10734), .CK(N28803), .QN(n7937) );
  DFF_X1 \CACHE_MEM_reg[2][133]  ( .D(n10733), .CK(N28803), .QN(n7953) );
  DFF_X1 \CACHE_MEM_reg[2][132]  ( .D(n10732), .CK(N28803), .QN(n7969) );
  DFF_X1 \CACHE_MEM_reg[2][131]  ( .D(n10731), .CK(N28803), .QN(n7985) );
  DFF_X1 \CACHE_MEM_reg[2][130]  ( .D(n10730), .CK(N28803), .QN(n8001) );
  DFF_X1 \CACHE_MEM_reg[2][129]  ( .D(n10729), .CK(N28803), .QN(n8017) );
  DFF_X1 \CACHE_MEM_reg[2][128]  ( .D(n10728), .CK(N28803), .QN(n8033) );
  DFF_X1 \CACHE_MEM_reg[2][127]  ( .D(n10727), .CK(N28803), .QN(n8049) );
  DFF_X1 \CACHE_MEM_reg[2][126]  ( .D(n10726), .CK(N28803), .QN(n8065) );
  DFF_X1 \CACHE_MEM_reg[2][125]  ( .D(n10725), .CK(N28803), .QN(n8081) );
  DFF_X1 \CACHE_MEM_reg[2][124]  ( .D(n10724), .CK(N28803), .QN(n8097) );
  DFF_X1 \CACHE_MEM_reg[2][123]  ( .D(n10723), .CK(N28803), .QN(n8113) );
  DFF_X1 \CACHE_MEM_reg[2][122]  ( .D(n10722), .CK(N28803), .QN(n8129) );
  DFF_X1 \CACHE_MEM_reg[2][121]  ( .D(n10721), .CK(N28803), .QN(n8145) );
  DFF_X1 \CACHE_MEM_reg[2][120]  ( .D(n10720), .CK(N28803), .QN(n8161) );
  DFF_X1 \CACHE_MEM_reg[2][119]  ( .D(n10719), .CK(N28803), .QN(n8177) );
  DFF_X1 \CACHE_MEM_reg[2][118]  ( .D(n10718), .CK(N28803), .QN(n8193) );
  DFF_X1 \CACHE_MEM_reg[2][117]  ( .D(n10717), .CK(N28803), .QN(n8209) );
  DFF_X1 \CACHE_MEM_reg[2][116]  ( .D(n10716), .CK(N28803), .QN(n8225) );
  DFF_X1 \CACHE_MEM_reg[2][115]  ( .D(n10715), .CK(N28803), .QN(n8241) );
  DFF_X1 \CACHE_MEM_reg[2][114]  ( .D(n10714), .CK(N28803), .QN(n8257) );
  DFF_X1 \CACHE_MEM_reg[2][113]  ( .D(n10713), .CK(N28803), .QN(n8273) );
  DFF_X1 \CACHE_MEM_reg[2][112]  ( .D(n10712), .CK(N28803), .QN(n8289) );
  DFF_X1 \CACHE_MEM_reg[2][111]  ( .D(n10711), .CK(N28803), .QN(n8305) );
  DFF_X1 \CACHE_MEM_reg[2][110]  ( .D(n10710), .CK(N28803), .QN(n8321) );
  DFF_X1 \CACHE_MEM_reg[2][109]  ( .D(n10709), .CK(N28803), .QN(n8337) );
  DFF_X1 \CACHE_MEM_reg[2][108]  ( .D(n10708), .CK(N28803), .QN(n8353) );
  DFF_X1 \CACHE_MEM_reg[2][107]  ( .D(n10707), .CK(N28803), .QN(n8369) );
  DFF_X1 \CACHE_MEM_reg[2][106]  ( .D(n10706), .CK(N28803), .QN(n8385) );
  DFF_X1 \CACHE_MEM_reg[2][105]  ( .D(n10705), .CK(N28803), .QN(n8401) );
  DFF_X1 \CACHE_MEM_reg[2][104]  ( .D(n10704), .CK(N28803), .QN(n8417) );
  DFF_X1 \CACHE_MEM_reg[2][103]  ( .D(n10703), .CK(N28803), .QN(n8433) );
  DFF_X1 \CACHE_MEM_reg[2][102]  ( .D(n10702), .CK(N28803), .QN(n8449) );
  DFF_X1 \CACHE_MEM_reg[2][101]  ( .D(n10701), .CK(N28803), .QN(n8465) );
  DFF_X1 \CACHE_MEM_reg[2][100]  ( .D(n10700), .CK(N28803), .QN(n8481) );
  DFF_X1 \CACHE_MEM_reg[2][99]  ( .D(n10699), .CK(N28803), .QN(n8497) );
  DFF_X1 \CACHE_MEM_reg[2][98]  ( .D(n10698), .CK(N28803), .QN(n8513) );
  DFF_X1 \CACHE_MEM_reg[2][97]  ( .D(n10697), .CK(N28803), .QN(n8529) );
  DFF_X1 \CACHE_MEM_reg[2][96]  ( .D(n10696), .CK(N28803), .QN(n8545) );
  DFF_X1 \CACHE_MEM_reg[2][95]  ( .D(n10695), .CK(N28803), .QN(n8561) );
  DFF_X1 \CACHE_MEM_reg[2][94]  ( .D(n10694), .CK(N28803), .QN(n8577) );
  DFF_X1 \CACHE_MEM_reg[2][93]  ( .D(n10693), .CK(N28803), .QN(n8593) );
  DFF_X1 \CACHE_MEM_reg[2][92]  ( .D(n10692), .CK(N28803), .QN(n8609) );
  DFF_X1 \CACHE_MEM_reg[2][91]  ( .D(n10691), .CK(N28803), .QN(n8625) );
  DFF_X1 \CACHE_MEM_reg[2][90]  ( .D(n10690), .CK(N28803), .QN(n8641) );
  DFF_X1 \CACHE_MEM_reg[2][89]  ( .D(n10689), .CK(N28803), .QN(n8657) );
  DFF_X1 \CACHE_MEM_reg[2][88]  ( .D(n10688), .CK(N28803), .QN(n8673) );
  DFF_X1 \CACHE_MEM_reg[2][87]  ( .D(n10687), .CK(N28803), .QN(n8689) );
  DFF_X1 \CACHE_MEM_reg[2][86]  ( .D(n10686), .CK(N28803), .QN(n8705) );
  DFF_X1 \CACHE_MEM_reg[2][85]  ( .D(n10685), .CK(N28803), .QN(n8721) );
  DFF_X1 \CACHE_MEM_reg[2][84]  ( .D(n10684), .CK(N28803), .QN(n8737) );
  DFF_X1 \CACHE_MEM_reg[2][83]  ( .D(n10683), .CK(N28803), .QN(n8753) );
  DFF_X1 \CACHE_MEM_reg[2][82]  ( .D(n10682), .CK(N28803), .QN(n8769) );
  DFF_X1 \CACHE_MEM_reg[2][81]  ( .D(n10681), .CK(N28803), .QN(n8785) );
  DFF_X1 \CACHE_MEM_reg[2][80]  ( .D(n10680), .CK(N28803), .QN(n8801) );
  DFF_X1 \CACHE_MEM_reg[2][79]  ( .D(n10679), .CK(N28803), .QN(n8817) );
  DFF_X1 \CACHE_MEM_reg[2][78]  ( .D(n10678), .CK(N28803), .QN(n8833) );
  DFF_X1 \CACHE_MEM_reg[2][77]  ( .D(n10677), .CK(N28803), .QN(n8849) );
  DFF_X1 \CACHE_MEM_reg[2][76]  ( .D(n10676), .CK(N28803), .QN(n8865) );
  DFF_X1 \CACHE_MEM_reg[2][75]  ( .D(n10675), .CK(N28803), .QN(n8881) );
  DFF_X1 \CACHE_MEM_reg[2][74]  ( .D(n10674), .CK(N28803), .QN(n8897) );
  DFF_X1 \CACHE_MEM_reg[2][73]  ( .D(n10673), .CK(N28803), .QN(n8913) );
  DFF_X1 \CACHE_MEM_reg[2][72]  ( .D(n10672), .CK(N28803), .QN(n8929) );
  DFF_X1 \CACHE_MEM_reg[2][71]  ( .D(n10671), .CK(N28803), .QN(n8945) );
  DFF_X1 \CACHE_MEM_reg[2][70]  ( .D(n10670), .CK(N28803), .QN(n8961) );
  DFF_X1 \CACHE_MEM_reg[2][69]  ( .D(n10669), .CK(N28803), .QN(n8977) );
  DFF_X1 \CACHE_MEM_reg[2][68]  ( .D(n10668), .CK(N28803), .QN(n8993) );
  DFF_X1 \CACHE_MEM_reg[2][67]  ( .D(n10667), .CK(N28803), .QN(n9009) );
  DFF_X1 \CACHE_MEM_reg[2][66]  ( .D(n10666), .CK(N28803), .QN(n9025) );
  DFF_X1 \CACHE_MEM_reg[2][65]  ( .D(n10665), .CK(N28803), .QN(n9041) );
  DFF_X1 \CACHE_MEM_reg[2][64]  ( .D(n10664), .CK(N28803), .QN(n9057) );
  DFF_X1 \CACHE_MEM_reg[2][63]  ( .D(n10663), .CK(N28803), .QN(n9073) );
  DFF_X1 \CACHE_MEM_reg[2][62]  ( .D(n10662), .CK(N28803), .QN(n9089) );
  DFF_X1 \CACHE_MEM_reg[2][61]  ( .D(n10661), .CK(N28803), .QN(n9105) );
  DFF_X1 \CACHE_MEM_reg[2][60]  ( .D(n10660), .CK(N28803), .QN(n9121) );
  DFF_X1 \CACHE_MEM_reg[2][59]  ( .D(n10659), .CK(N28803), .QN(n9137) );
  DFF_X1 \CACHE_MEM_reg[2][58]  ( .D(n10658), .CK(N28803), .QN(n9153) );
  DFF_X1 \CACHE_MEM_reg[2][57]  ( .D(n10657), .CK(N28803), .QN(n9169) );
  DFF_X1 \CACHE_MEM_reg[2][56]  ( .D(n10656), .CK(N28803), .QN(n9185) );
  DFF_X1 \CACHE_MEM_reg[2][55]  ( .D(n10655), .CK(N28803), .QN(n9201) );
  DFF_X1 \CACHE_MEM_reg[2][54]  ( .D(n10654), .CK(N28803), .QN(n9217) );
  DFF_X1 \CACHE_MEM_reg[2][53]  ( .D(n10653), .CK(N28803), .QN(n9233) );
  DFF_X1 \CACHE_MEM_reg[2][52]  ( .D(n10652), .CK(N28803), .QN(n9249) );
  DFF_X1 \CACHE_MEM_reg[2][51]  ( .D(n10651), .CK(N28803), .QN(n9265) );
  DFF_X1 \CACHE_MEM_reg[2][50]  ( .D(n10650), .CK(N28803), .QN(n9281) );
  DFF_X1 \CACHE_MEM_reg[2][49]  ( .D(n10649), .CK(N28803), .QN(n9297) );
  DFF_X1 \CACHE_MEM_reg[2][48]  ( .D(n10648), .CK(N28803), .QN(n9313) );
  DFF_X1 \CACHE_MEM_reg[2][47]  ( .D(n10647), .CK(N28803), .QN(n9329) );
  DFF_X1 \CACHE_MEM_reg[2][46]  ( .D(n10646), .CK(N28803), .QN(n9345) );
  DFF_X1 \CACHE_MEM_reg[2][45]  ( .D(n10645), .CK(N28803), .QN(n9361) );
  DFF_X1 \CACHE_MEM_reg[2][44]  ( .D(n10644), .CK(N28803), .QN(n9377) );
  DFF_X1 \CACHE_MEM_reg[2][43]  ( .D(n10643), .CK(N28803), .QN(n9393) );
  DFF_X1 \CACHE_MEM_reg[2][42]  ( .D(n10642), .CK(N28803), .QN(n9409) );
  DFF_X1 \CACHE_MEM_reg[2][41]  ( .D(n10641), .CK(N28803), .QN(n9425) );
  DFF_X1 \CACHE_MEM_reg[2][40]  ( .D(n10640), .CK(N28803), .QN(n9441) );
  DFF_X1 \CACHE_MEM_reg[2][39]  ( .D(n10639), .CK(N28803), .QN(n9457) );
  DFF_X1 \CACHE_MEM_reg[2][38]  ( .D(n10638), .CK(N28803), .QN(n9473) );
  DFF_X1 \CACHE_MEM_reg[2][37]  ( .D(n10637), .CK(N28803), .QN(n9489) );
  DFF_X1 \CACHE_MEM_reg[2][36]  ( .D(n10636), .CK(N28803), .QN(n9505) );
  DFF_X1 \CACHE_MEM_reg[2][35]  ( .D(n10635), .CK(N28803), .QN(n9521) );
  DFF_X1 \CACHE_MEM_reg[2][34]  ( .D(n10634), .CK(N28803), .QN(n9537) );
  DFF_X1 \CACHE_MEM_reg[2][33]  ( .D(n10633), .CK(N28803), .QN(n9553) );
  DFF_X1 \CACHE_MEM_reg[2][32]  ( .D(n10632), .CK(N28803), .QN(n9569) );
  DFF_X1 \CACHE_MEM_reg[2][31]  ( .D(n10631), .CK(N28803), .QN(n9585) );
  DFF_X1 \CACHE_MEM_reg[2][30]  ( .D(n10630), .CK(N28803), .QN(n9601) );
  DFF_X1 \CACHE_MEM_reg[2][29]  ( .D(n10629), .CK(N28803), .QN(n9617) );
  DFF_X1 \CACHE_MEM_reg[2][28]  ( .D(n10628), .CK(N28803), .QN(n9633) );
  DFF_X1 \CACHE_MEM_reg[2][27]  ( .D(n10627), .CK(N28803), .QN(n9649) );
  DFF_X1 \CACHE_MEM_reg[2][26]  ( .D(n10626), .CK(N28803), .QN(n9665) );
  DFF_X1 \CACHE_MEM_reg[2][25]  ( .D(n10625), .CK(N28803), .QN(n9681) );
  DFF_X1 \CACHE_MEM_reg[2][24]  ( .D(n10624), .CK(N28803), .QN(n9697) );
  DFF_X1 \CACHE_MEM_reg[2][23]  ( .D(n10623), .CK(N28803), .QN(n9713) );
  DFF_X1 \CACHE_MEM_reg[2][22]  ( .D(n10622), .CK(N28803), .QN(n9729) );
  DFF_X1 \CACHE_MEM_reg[2][21]  ( .D(n10621), .CK(N28803), .QN(n9745) );
  DFF_X1 \CACHE_MEM_reg[2][20]  ( .D(n10620), .CK(N28803), .QN(n9761) );
  DFF_X1 \CACHE_MEM_reg[2][19]  ( .D(n10619), .CK(N28803), .QN(n9777) );
  DFF_X1 \CACHE_MEM_reg[2][18]  ( .D(n10618), .CK(N28803), .QN(n9793) );
  DFF_X1 \CACHE_MEM_reg[2][17]  ( .D(n10617), .CK(N28803), .QN(n9809) );
  DFF_X1 \CACHE_MEM_reg[2][16]  ( .D(n10616), .CK(N28803), .QN(n9825) );
  DFF_X1 \CACHE_MEM_reg[2][15]  ( .D(n10615), .CK(N28803), .QN(n9841) );
  DFF_X1 \CACHE_MEM_reg[2][14]  ( .D(n10614), .CK(N28803), .QN(n9857) );
  DFF_X1 \CACHE_MEM_reg[2][13]  ( .D(n10613), .CK(N28803), .QN(n9873) );
  DFF_X1 \CACHE_MEM_reg[2][12]  ( .D(n10612), .CK(N28803), .QN(n9889) );
  DFF_X1 \CACHE_MEM_reg[2][11]  ( .D(n10611), .CK(N28803), .QN(n9905) );
  DFF_X1 \CACHE_MEM_reg[2][10]  ( .D(n10610), .CK(N28803), .QN(n9921) );
  DFF_X1 \CACHE_MEM_reg[2][9]  ( .D(n10609), .CK(N28803), .QN(n9937) );
  DFF_X1 \CACHE_MEM_reg[2][8]  ( .D(n10608), .CK(N28803), .QN(n9953) );
  DFF_X1 \CACHE_MEM_reg[2][7]  ( .D(n10607), .CK(N28803), .QN(n9969) );
  DFF_X1 \CACHE_MEM_reg[2][6]  ( .D(n10606), .CK(N28803), .QN(n9985) );
  DFF_X1 \CACHE_MEM_reg[2][5]  ( .D(n10605), .CK(N28803), .QN(n10001) );
  DFF_X1 \CACHE_MEM_reg[2][4]  ( .D(n10604), .CK(N28803), .QN(n10017) );
  DFF_X1 \CACHE_MEM_reg[2][3]  ( .D(n10603), .CK(N28803), .QN(n10033) );
  DFF_X1 \CACHE_MEM_reg[2][2]  ( .D(n10602), .CK(N28803), .QN(n10049) );
  DFF_X1 \CACHE_MEM_reg[2][1]  ( .D(n10601), .CK(N28803), .QN(n10065) );
  DFF_X1 \CACHE_MEM_reg[2][0]  ( .D(n10600), .CK(N28803), .QN(n10081) );
  DFF_X1 \CACHE_MEM_reg[1][255]  ( .D(n10599), .CK(N28803), .Q(n167), .QN(
        n5997) );
  DFF_X1 \CACHE_MEM_reg[1][254]  ( .D(n10598), .CK(N28803), .Q(n155), .QN(
        n6013) );
  DFF_X1 \CACHE_MEM_reg[1][253]  ( .D(n10597), .CK(N28803), .Q(n146), .QN(
        n6029) );
  DFF_X1 \CACHE_MEM_reg[1][252]  ( .D(n10596), .CK(N28803), .Q(n137), .QN(
        n6045) );
  DFF_X1 \CACHE_MEM_reg[1][251]  ( .D(n10595), .CK(N28803), .Q(n128), .QN(
        n6061) );
  DFF_X1 \CACHE_MEM_reg[1][250]  ( .D(n10594), .CK(N28803), .Q(n119), .QN(
        n6077) );
  DFF_X1 \CACHE_MEM_reg[1][249]  ( .D(n10593), .CK(N28803), .Q(n110), .QN(
        n6093) );
  DFF_X1 \CACHE_MEM_reg[1][248]  ( .D(n10592), .CK(N28803), .Q(n101), .QN(
        n6109) );
  DFF_X1 \CACHE_MEM_reg[1][247]  ( .D(n10591), .CK(N28803), .Q(n92), .QN(n6125) );
  DFF_X1 \CACHE_MEM_reg[1][246]  ( .D(n10590), .CK(N28803), .Q(n83), .QN(n6141) );
  DFF_X1 \CACHE_MEM_reg[1][245]  ( .D(n10589), .CK(N28803), .Q(n65), .QN(n6157) );
  DFF_X1 \CACHE_MEM_reg[1][244]  ( .D(n10588), .CK(N28803), .Q(n62), .QN(n6173) );
  DFF_X1 \CACHE_MEM_reg[1][243]  ( .D(n10587), .CK(N28803), .Q(n59), .QN(n6189) );
  DFF_X1 \CACHE_MEM_reg[1][242]  ( .D(n10586), .CK(N28803), .Q(n56), .QN(n6205) );
  DFF_X1 \CACHE_MEM_reg[1][241]  ( .D(n10585), .CK(N28803), .Q(n53), .QN(n6221) );
  DFF_X1 \CACHE_MEM_reg[1][240]  ( .D(n10584), .CK(N28803), .Q(n50), .QN(n6237) );
  DFF_X1 \CACHE_MEM_reg[1][239]  ( .D(n10583), .CK(N28803), .Q(n47), .QN(n6253) );
  DFF_X1 \CACHE_MEM_reg[1][238]  ( .D(n10582), .CK(N28803), .Q(n44), .QN(n6269) );
  DFF_X1 \CACHE_MEM_reg[1][237]  ( .D(n10581), .CK(N28803), .Q(n41), .QN(n6285) );
  DFF_X1 \CACHE_MEM_reg[1][236]  ( .D(n10580), .CK(N28803), .Q(n38), .QN(n6301) );
  DFF_X1 \CACHE_MEM_reg[1][235]  ( .D(n10579), .CK(N28803), .Q(n35), .QN(n6317) );
  DFF_X1 \CACHE_MEM_reg[1][234]  ( .D(n10578), .CK(N28803), .Q(n32), .QN(n6333) );
  DFF_X1 \CACHE_MEM_reg[1][233]  ( .D(n10577), .CK(N28803), .Q(n29), .QN(n6349) );
  DFF_X1 \CACHE_MEM_reg[1][232]  ( .D(n10576), .CK(N28803), .Q(n26), .QN(n6365) );
  DFF_X1 \CACHE_MEM_reg[1][231]  ( .D(n10575), .CK(N28803), .Q(n23), .QN(n6381) );
  DFF_X1 \CACHE_MEM_reg[1][230]  ( .D(n10574), .CK(N28803), .Q(n20), .QN(n6397) );
  DFF_X1 \CACHE_MEM_reg[1][229]  ( .D(n10573), .CK(N28803), .Q(n17), .QN(n6413) );
  DFF_X1 \CACHE_MEM_reg[1][228]  ( .D(n10572), .CK(N28803), .Q(n14), .QN(n6429) );
  DFF_X1 \CACHE_MEM_reg[1][227]  ( .D(n10571), .CK(N28803), .Q(n11), .QN(n6445) );
  DFF_X1 \CACHE_MEM_reg[1][226]  ( .D(n10570), .CK(N28803), .Q(n8), .QN(n6461)
         );
  DFF_X1 \CACHE_MEM_reg[1][225]  ( .D(n10569), .CK(N28803), .Q(n5), .QN(n6477)
         );
  DFF_X1 \CACHE_MEM_reg[1][224]  ( .D(n10568), .CK(N28803), .Q(n2), .QN(n6493)
         );
  DFF_X1 \CACHE_MEM_reg[1][223]  ( .D(n10567), .CK(N28803), .Q(n2879), .QN(
        n6509) );
  DFF_X1 \CACHE_MEM_reg[1][222]  ( .D(n10566), .CK(N28803), .Q(n2862), .QN(
        n6525) );
  DFF_X1 \CACHE_MEM_reg[1][221]  ( .D(n10565), .CK(N28803), .Q(n2851), .QN(
        n6541) );
  DFF_X1 \CACHE_MEM_reg[1][220]  ( .D(n10564), .CK(N28803), .Q(n2838), .QN(
        n6557) );
  DFF_X1 \CACHE_MEM_reg[1][219]  ( .D(n10563), .CK(N28803), .Q(n2818), .QN(
        n6573) );
  DFF_X1 \CACHE_MEM_reg[1][218]  ( .D(n10562), .CK(N28803), .Q(n2805), .QN(
        n6589) );
  DFF_X1 \CACHE_MEM_reg[1][217]  ( .D(n10561), .CK(N28803), .Q(n2794), .QN(
        n6605) );
  DFF_X1 \CACHE_MEM_reg[1][216]  ( .D(n10560), .CK(N28803), .Q(n2777), .QN(
        n6621) );
  DFF_X1 \CACHE_MEM_reg[1][215]  ( .D(n10559), .CK(N28803), .Q(n2766), .QN(
        n6637) );
  DFF_X1 \CACHE_MEM_reg[1][214]  ( .D(n10558), .CK(N28803), .Q(n2749), .QN(
        n6653) );
  DFF_X1 \CACHE_MEM_reg[1][213]  ( .D(n10557), .CK(N28803), .Q(n2738), .QN(
        n6669) );
  DFF_X1 \CACHE_MEM_reg[1][212]  ( .D(n10556), .CK(N28803), .Q(n2725), .QN(
        n6685) );
  DFF_X1 \CACHE_MEM_reg[1][211]  ( .D(n10555), .CK(N28803), .Q(n2710), .QN(
        n6701) );
  DFF_X1 \CACHE_MEM_reg[1][210]  ( .D(n10554), .CK(N28803), .Q(n2697), .QN(
        n6717) );
  DFF_X1 \CACHE_MEM_reg[1][209]  ( .D(n10553), .CK(N28803), .Q(n2686), .QN(
        n6733) );
  DFF_X1 \CACHE_MEM_reg[1][208]  ( .D(n10552), .CK(N28803), .Q(n2669), .QN(
        n6749) );
  DFF_X1 \CACHE_MEM_reg[1][207]  ( .D(n10551), .CK(N28803), .Q(n2656), .QN(
        n6765) );
  DFF_X1 \CACHE_MEM_reg[1][206]  ( .D(n10550), .CK(N28803), .Q(n2645), .QN(
        n6781) );
  DFF_X1 \CACHE_MEM_reg[1][205]  ( .D(n10549), .CK(N28803), .Q(n2628), .QN(
        n6797) );
  DFF_X1 \CACHE_MEM_reg[1][204]  ( .D(n10548), .CK(N28803), .Q(n2617), .QN(
        n6813) );
  DFF_X1 \CACHE_MEM_reg[1][203]  ( .D(n10547), .CK(N28803), .Q(n2600), .QN(
        n6829) );
  DFF_X1 \CACHE_MEM_reg[1][202]  ( .D(n10546), .CK(N28803), .Q(n2589), .QN(
        n6845) );
  DFF_X1 \CACHE_MEM_reg[1][201]  ( .D(n10545), .CK(N28803), .Q(n2576), .QN(
        n6861) );
  DFF_X1 \CACHE_MEM_reg[1][200]  ( .D(n10544), .CK(N28803), .Q(n2561), .QN(
        n6877) );
  DFF_X1 \CACHE_MEM_reg[1][199]  ( .D(n10543), .CK(N28803), .Q(n2548), .QN(
        n6893) );
  DFF_X1 \CACHE_MEM_reg[1][198]  ( .D(n10542), .CK(N28803), .Q(n2537), .QN(
        n6909) );
  DFF_X1 \CACHE_MEM_reg[1][197]  ( .D(n10541), .CK(N28803), .Q(n2515), .QN(
        n6925) );
  DFF_X1 \CACHE_MEM_reg[1][196]  ( .D(n10540), .CK(N28803), .Q(n2504), .QN(
        n6941) );
  DFF_X1 \CACHE_MEM_reg[1][195]  ( .D(n10539), .CK(N28803), .Q(n2487), .QN(
        n6957) );
  DFF_X1 \CACHE_MEM_reg[1][194]  ( .D(n10538), .CK(N28803), .Q(n2476), .QN(
        n6973) );
  DFF_X1 \CACHE_MEM_reg[1][193]  ( .D(n10537), .CK(N28803), .Q(n2463), .QN(
        n6989) );
  DFF_X1 \CACHE_MEM_reg[1][192]  ( .D(n10536), .CK(N28803), .Q(n2448), .QN(
        n7005) );
  DFF_X1 \CACHE_MEM_reg[1][191]  ( .D(n10535), .CK(N28803), .Q(n3321), .QN(
        n7021) );
  DFF_X1 \CACHE_MEM_reg[1][190]  ( .D(n10534), .CK(N28803), .Q(n158), .QN(
        n7037) );
  DFF_X1 \CACHE_MEM_reg[1][189]  ( .D(n10533), .CK(N28803), .Q(n149), .QN(
        n7053) );
  DFF_X1 \CACHE_MEM_reg[1][188]  ( .D(n10532), .CK(N28803), .Q(n140), .QN(
        n7069) );
  DFF_X1 \CACHE_MEM_reg[1][187]  ( .D(n10531), .CK(N28803), .Q(n131), .QN(
        n7085) );
  DFF_X1 \CACHE_MEM_reg[1][186]  ( .D(n10530), .CK(N28803), .Q(n122), .QN(
        n7101) );
  DFF_X1 \CACHE_MEM_reg[1][185]  ( .D(n10529), .CK(N28803), .Q(n113), .QN(
        n7117) );
  DFF_X1 \CACHE_MEM_reg[1][184]  ( .D(n10528), .CK(N28803), .Q(n104), .QN(
        n7133) );
  DFF_X1 \CACHE_MEM_reg[1][183]  ( .D(n10527), .CK(N28803), .Q(n95), .QN(n7149) );
  DFF_X1 \CACHE_MEM_reg[1][182]  ( .D(n10526), .CK(N28803), .Q(n86), .QN(n7165) );
  DFF_X1 \CACHE_MEM_reg[1][181]  ( .D(n10525), .CK(N28803), .Q(n76), .QN(n7181) );
  DFF_X1 \CACHE_MEM_reg[1][180]  ( .D(n10524), .CK(N28803), .Q(n63), .QN(n7197) );
  DFF_X1 \CACHE_MEM_reg[1][179]  ( .D(n10523), .CK(N28803), .Q(n60), .QN(n7213) );
  DFF_X1 \CACHE_MEM_reg[1][178]  ( .D(n10522), .CK(N28803), .Q(n57), .QN(n7229) );
  DFF_X1 \CACHE_MEM_reg[1][177]  ( .D(n10521), .CK(N28803), .Q(n54), .QN(n7245) );
  DFF_X1 \CACHE_MEM_reg[1][176]  ( .D(n10520), .CK(N28803), .Q(n51), .QN(n7261) );
  DFF_X1 \CACHE_MEM_reg[1][175]  ( .D(n10519), .CK(N28803), .Q(n48), .QN(n7277) );
  DFF_X1 \CACHE_MEM_reg[1][174]  ( .D(n10518), .CK(N28803), .Q(n45), .QN(n7293) );
  DFF_X1 \CACHE_MEM_reg[1][173]  ( .D(n10517), .CK(N28803), .Q(n42), .QN(n7309) );
  DFF_X1 \CACHE_MEM_reg[1][172]  ( .D(n10516), .CK(N28803), .Q(n39), .QN(n7325) );
  DFF_X1 \CACHE_MEM_reg[1][171]  ( .D(n10515), .CK(N28803), .Q(n36), .QN(n7341) );
  DFF_X1 \CACHE_MEM_reg[1][170]  ( .D(n10514), .CK(N28803), .Q(n33), .QN(n7357) );
  DFF_X1 \CACHE_MEM_reg[1][169]  ( .D(n10513), .CK(N28803), .Q(n30), .QN(n7373) );
  DFF_X1 \CACHE_MEM_reg[1][168]  ( .D(n10512), .CK(N28803), .Q(n27), .QN(n7389) );
  DFF_X1 \CACHE_MEM_reg[1][167]  ( .D(n10511), .CK(N28803), .Q(n24), .QN(n7405) );
  DFF_X1 \CACHE_MEM_reg[1][166]  ( .D(n10510), .CK(N28803), .Q(n21), .QN(n7421) );
  DFF_X1 \CACHE_MEM_reg[1][165]  ( .D(n10509), .CK(N28803), .Q(n18), .QN(n7437) );
  DFF_X1 \CACHE_MEM_reg[1][164]  ( .D(n10508), .CK(N28803), .Q(n15), .QN(n7453) );
  DFF_X1 \CACHE_MEM_reg[1][163]  ( .D(n10507), .CK(N28803), .Q(n12), .QN(n7469) );
  DFF_X1 \CACHE_MEM_reg[1][162]  ( .D(n10506), .CK(N28803), .Q(n9), .QN(n7485)
         );
  DFF_X1 \CACHE_MEM_reg[1][161]  ( .D(n10505), .CK(N28803), .Q(n6), .QN(n7501)
         );
  DFF_X1 \CACHE_MEM_reg[1][160]  ( .D(n10504), .CK(N28803), .Q(n3), .QN(n7517)
         );
  DFF_X1 \CACHE_MEM_reg[1][159]  ( .D(n10503), .CK(N28803), .Q(n3326), .QN(
        n7533) );
  DFF_X1 \CACHE_MEM_reg[1][158]  ( .D(n10502), .CK(N28803), .Q(n3309), .QN(
        n7549) );
  DFF_X1 \CACHE_MEM_reg[1][157]  ( .D(n10501), .CK(N28803), .Q(n3298), .QN(
        n7565) );
  DFF_X1 \CACHE_MEM_reg[1][156]  ( .D(n10500), .CK(N28803), .Q(n3285), .QN(
        n7581) );
  DFF_X1 \CACHE_MEM_reg[1][155]  ( .D(n10499), .CK(N28803), .Q(n3265), .QN(
        n7597) );
  DFF_X1 \CACHE_MEM_reg[1][154]  ( .D(n10498), .CK(N28803), .Q(n3252), .QN(
        n7613) );
  DFF_X1 \CACHE_MEM_reg[1][153]  ( .D(n10497), .CK(N28803), .Q(n3241), .QN(
        n7629) );
  DFF_X1 \CACHE_MEM_reg[1][152]  ( .D(n10496), .CK(N28803), .Q(n3224), .QN(
        n7645) );
  DFF_X1 \CACHE_MEM_reg[1][151]  ( .D(n10495), .CK(N28803), .Q(n3213), .QN(
        n7661) );
  DFF_X1 \CACHE_MEM_reg[1][150]  ( .D(n10494), .CK(N28803), .Q(n3196), .QN(
        n7677) );
  DFF_X1 \CACHE_MEM_reg[1][149]  ( .D(n10493), .CK(N28803), .Q(n3185), .QN(
        n7693) );
  DFF_X1 \CACHE_MEM_reg[1][148]  ( .D(n10492), .CK(N28803), .Q(n3172), .QN(
        n7709) );
  DFF_X1 \CACHE_MEM_reg[1][147]  ( .D(n10491), .CK(N28803), .Q(n3157), .QN(
        n7725) );
  DFF_X1 \CACHE_MEM_reg[1][146]  ( .D(n10490), .CK(N28803), .Q(n3144), .QN(
        n7741) );
  DFF_X1 \CACHE_MEM_reg[1][145]  ( .D(n10489), .CK(N28803), .Q(n3133), .QN(
        n7757) );
  DFF_X1 \CACHE_MEM_reg[1][144]  ( .D(n10488), .CK(N28803), .Q(n3111), .QN(
        n7773) );
  DFF_X1 \CACHE_MEM_reg[1][143]  ( .D(n10487), .CK(N28803), .Q(n3100), .QN(
        n7789) );
  DFF_X1 \CACHE_MEM_reg[1][142]  ( .D(n10486), .CK(N28803), .Q(n3083), .QN(
        n7805) );
  DFF_X1 \CACHE_MEM_reg[1][141]  ( .D(n10485), .CK(N28803), .Q(n3072), .QN(
        n7821) );
  DFF_X1 \CACHE_MEM_reg[1][140]  ( .D(n10484), .CK(N28803), .Q(n3059), .QN(
        n7837) );
  DFF_X1 \CACHE_MEM_reg[1][139]  ( .D(n10483), .CK(N28803), .Q(n3044), .QN(
        n7853) );
  DFF_X1 \CACHE_MEM_reg[1][138]  ( .D(n10482), .CK(N28803), .Q(n3031), .QN(
        n7869) );
  DFF_X1 \CACHE_MEM_reg[1][137]  ( .D(n10481), .CK(N28803), .Q(n3020), .QN(
        n7885) );
  DFF_X1 \CACHE_MEM_reg[1][136]  ( .D(n10480), .CK(N28803), .Q(n3003), .QN(
        n7901) );
  DFF_X1 \CACHE_MEM_reg[1][135]  ( .D(n10479), .CK(N28803), .Q(n2992), .QN(
        n7917) );
  DFF_X1 \CACHE_MEM_reg[1][134]  ( .D(n10478), .CK(N28803), .Q(n2970), .QN(
        n7933) );
  DFF_X1 \CACHE_MEM_reg[1][133]  ( .D(n10477), .CK(N28803), .Q(n2959), .QN(
        n7949) );
  DFF_X1 \CACHE_MEM_reg[1][132]  ( .D(n10476), .CK(N28803), .Q(n2946), .QN(
        n7965) );
  DFF_X1 \CACHE_MEM_reg[1][131]  ( .D(n10475), .CK(N28803), .Q(n2931), .QN(
        n7981) );
  DFF_X1 \CACHE_MEM_reg[1][130]  ( .D(n10474), .CK(N28803), .Q(n2918), .QN(
        n7997) );
  DFF_X1 \CACHE_MEM_reg[1][129]  ( .D(n10473), .CK(N28803), .Q(n2907), .QN(
        n8013) );
  DFF_X1 \CACHE_MEM_reg[1][128]  ( .D(n10472), .CK(N28803), .Q(n2890), .QN(
        n8029) );
  DFF_X1 \CACHE_MEM_reg[1][127]  ( .D(n10471), .CK(N28803), .Q(n161), .QN(
        n8045) );
  DFF_X1 \CACHE_MEM_reg[1][126]  ( .D(n10470), .CK(N28803), .Q(n1968), .QN(
        n8061) );
  DFF_X1 \CACHE_MEM_reg[1][125]  ( .D(n10469), .CK(N28803), .Q(n1952), .QN(
        n8077) );
  DFF_X1 \CACHE_MEM_reg[1][124]  ( .D(n10468), .CK(N28803), .Q(n1927), .QN(
        n8093) );
  DFF_X1 \CACHE_MEM_reg[1][123]  ( .D(n10467), .CK(N28803), .Q(n1911), .QN(
        n8109) );
  DFF_X1 \CACHE_MEM_reg[1][122]  ( .D(n10466), .CK(N28803), .Q(n1891), .QN(
        n8125) );
  DFF_X1 \CACHE_MEM_reg[1][121]  ( .D(n10465), .CK(N28803), .Q(n1875), .QN(
        n8141) );
  DFF_X1 \CACHE_MEM_reg[1][120]  ( .D(n10464), .CK(N28803), .Q(n1855), .QN(
        n8157) );
  DFF_X1 \CACHE_MEM_reg[1][119]  ( .D(n10463), .CK(N28803), .Q(n1839), .QN(
        n8173) );
  DFF_X1 \CACHE_MEM_reg[1][118]  ( .D(n10462), .CK(N28803), .Q(n1819), .QN(
        n8189) );
  DFF_X1 \CACHE_MEM_reg[1][117]  ( .D(n10461), .CK(N28803), .Q(n1803), .QN(
        n8205) );
  DFF_X1 \CACHE_MEM_reg[1][116]  ( .D(n10460), .CK(N28803), .Q(n1778), .QN(
        n8221) );
  DFF_X1 \CACHE_MEM_reg[1][115]  ( .D(n10459), .CK(N28803), .Q(n1762), .QN(
        n8237) );
  DFF_X1 \CACHE_MEM_reg[1][114]  ( .D(n10458), .CK(N28803), .Q(n1742), .QN(
        n8253) );
  DFF_X1 \CACHE_MEM_reg[1][113]  ( .D(n10457), .CK(N28803), .Q(n1726), .QN(
        n8269) );
  DFF_X1 \CACHE_MEM_reg[1][112]  ( .D(n10456), .CK(N28803), .Q(n1706), .QN(
        n8285) );
  DFF_X1 \CACHE_MEM_reg[1][111]  ( .D(n10455), .CK(N28803), .Q(n1690), .QN(
        n8301) );
  DFF_X1 \CACHE_MEM_reg[1][110]  ( .D(n10454), .CK(N28803), .Q(n1670), .QN(
        n8317) );
  DFF_X1 \CACHE_MEM_reg[1][109]  ( .D(n10453), .CK(N28803), .Q(n1654), .QN(
        n8333) );
  DFF_X1 \CACHE_MEM_reg[1][108]  ( .D(n10452), .CK(N28803), .Q(n1629), .QN(
        n8349) );
  DFF_X1 \CACHE_MEM_reg[1][107]  ( .D(n10451), .CK(N28803), .Q(n1613), .QN(
        n8365) );
  DFF_X1 \CACHE_MEM_reg[1][106]  ( .D(n10450), .CK(N28803), .Q(n1593), .QN(
        n8381) );
  DFF_X1 \CACHE_MEM_reg[1][105]  ( .D(n10449), .CK(N28803), .Q(n1577), .QN(
        n8397) );
  DFF_X1 \CACHE_MEM_reg[1][104]  ( .D(n10448), .CK(N28803), .Q(n1557), .QN(
        n8413) );
  DFF_X1 \CACHE_MEM_reg[1][103]  ( .D(n10447), .CK(N28803), .Q(n1541), .QN(
        n8429) );
  DFF_X1 \CACHE_MEM_reg[1][102]  ( .D(n10446), .CK(N28803), .Q(n1521), .QN(
        n8445) );
  DFF_X1 \CACHE_MEM_reg[1][101]  ( .D(n10445), .CK(N28803), .Q(n1505), .QN(
        n8461) );
  DFF_X1 \CACHE_MEM_reg[1][100]  ( .D(n10444), .CK(N28803), .Q(n1480), .QN(
        n8477) );
  DFF_X1 \CACHE_MEM_reg[1][99]  ( .D(n10443), .CK(N28803), .Q(n1464), .QN(
        n8493) );
  DFF_X1 \CACHE_MEM_reg[1][98]  ( .D(n10442), .CK(N28803), .Q(n1444), .QN(
        n8509) );
  DFF_X1 \CACHE_MEM_reg[1][97]  ( .D(n10441), .CK(N28803), .Q(n1428), .QN(
        n8525) );
  DFF_X1 \CACHE_MEM_reg[1][96]  ( .D(n10440), .CK(N28803), .Q(n1408), .QN(
        n8541) );
  DFF_X1 \CACHE_MEM_reg[1][95]  ( .D(n10439), .CK(N28803), .Q(n1988), .QN(
        n8557) );
  DFF_X1 \CACHE_MEM_reg[1][94]  ( .D(n10438), .CK(N28803), .Q(n1977), .QN(
        n8573) );
  DFF_X1 \CACHE_MEM_reg[1][93]  ( .D(n10437), .CK(N28803), .Q(n1957), .QN(
        n8589) );
  DFF_X1 \CACHE_MEM_reg[1][92]  ( .D(n10436), .CK(N28803), .Q(n1941), .QN(
        n8605) );
  DFF_X1 \CACHE_MEM_reg[1][91]  ( .D(n10435), .CK(N28803), .Q(n1916), .QN(
        n8621) );
  DFF_X1 \CACHE_MEM_reg[1][90]  ( .D(n10434), .CK(N28803), .Q(n1900), .QN(
        n8637) );
  DFF_X1 \CACHE_MEM_reg[1][89]  ( .D(n10433), .CK(N28803), .Q(n1880), .QN(
        n8653) );
  DFF_X1 \CACHE_MEM_reg[1][88]  ( .D(n10432), .CK(N28803), .Q(n1864), .QN(
        n8669) );
  DFF_X1 \CACHE_MEM_reg[1][87]  ( .D(n10431), .CK(N28803), .Q(n1844), .QN(
        n8685) );
  DFF_X1 \CACHE_MEM_reg[1][86]  ( .D(n10430), .CK(N28803), .Q(n1828), .QN(
        n8701) );
  DFF_X1 \CACHE_MEM_reg[1][85]  ( .D(n10429), .CK(N28803), .Q(n1808), .QN(
        n8717) );
  DFF_X1 \CACHE_MEM_reg[1][84]  ( .D(n10428), .CK(N28803), .Q(n1792), .QN(
        n8733) );
  DFF_X1 \CACHE_MEM_reg[1][83]  ( .D(n10427), .CK(N28803), .Q(n1767), .QN(
        n8749) );
  DFF_X1 \CACHE_MEM_reg[1][82]  ( .D(n10426), .CK(N28803), .Q(n1751), .QN(
        n8765) );
  DFF_X1 \CACHE_MEM_reg[1][81]  ( .D(n10425), .CK(N28803), .Q(n1731), .QN(
        n8781) );
  DFF_X1 \CACHE_MEM_reg[1][80]  ( .D(n10424), .CK(N28803), .Q(n1715), .QN(
        n8797) );
  DFF_X1 \CACHE_MEM_reg[1][79]  ( .D(n10423), .CK(N28803), .Q(n1695), .QN(
        n8813) );
  DFF_X1 \CACHE_MEM_reg[1][78]  ( .D(n10422), .CK(N28803), .Q(n1679), .QN(
        n8829) );
  DFF_X1 \CACHE_MEM_reg[1][77]  ( .D(n10421), .CK(N28803), .Q(n1659), .QN(
        n8845) );
  DFF_X1 \CACHE_MEM_reg[1][76]  ( .D(n10420), .CK(N28803), .Q(n1643), .QN(
        n8861) );
  DFF_X1 \CACHE_MEM_reg[1][75]  ( .D(n10419), .CK(N28803), .Q(n1618), .QN(
        n8877) );
  DFF_X1 \CACHE_MEM_reg[1][74]  ( .D(n10418), .CK(N28803), .Q(n1602), .QN(
        n8893) );
  DFF_X1 \CACHE_MEM_reg[1][73]  ( .D(n10417), .CK(N28803), .Q(n1582), .QN(
        n8909) );
  DFF_X1 \CACHE_MEM_reg[1][72]  ( .D(n10416), .CK(N28803), .Q(n1566), .QN(
        n8925) );
  DFF_X1 \CACHE_MEM_reg[1][71]  ( .D(n10415), .CK(N28803), .Q(n1546), .QN(
        n8941) );
  DFF_X1 \CACHE_MEM_reg[1][70]  ( .D(n10414), .CK(N28803), .Q(n1530), .QN(
        n8957) );
  DFF_X1 \CACHE_MEM_reg[1][69]  ( .D(n10413), .CK(N28803), .Q(n1510), .QN(
        n8973) );
  DFF_X1 \CACHE_MEM_reg[1][68]  ( .D(n10412), .CK(N28803), .Q(n1494), .QN(
        n8989) );
  DFF_X1 \CACHE_MEM_reg[1][67]  ( .D(n10411), .CK(N28803), .Q(n1469), .QN(
        n9005) );
  DFF_X1 \CACHE_MEM_reg[1][66]  ( .D(n10410), .CK(N28803), .Q(n1453), .QN(
        n9021) );
  DFF_X1 \CACHE_MEM_reg[1][65]  ( .D(n10409), .CK(N28803), .Q(n1433), .QN(
        n9037) );
  DFF_X1 \CACHE_MEM_reg[1][64]  ( .D(n10408), .CK(N28803), .Q(n1417), .QN(
        n9053) );
  DFF_X1 \CACHE_MEM_reg[1][63]  ( .D(n10407), .CK(N28803), .Q(n164), .QN(n9069) );
  DFF_X1 \CACHE_MEM_reg[1][62]  ( .D(n10406), .CK(N28803), .Q(n152), .QN(n9085) );
  DFF_X1 \CACHE_MEM_reg[1][61]  ( .D(n10405), .CK(N28803), .Q(n143), .QN(n9101) );
  DFF_X1 \CACHE_MEM_reg[1][60]  ( .D(n10404), .CK(N28803), .Q(n134), .QN(n9117) );
  DFF_X1 \CACHE_MEM_reg[1][59]  ( .D(n10403), .CK(N28803), .Q(n125), .QN(n9133) );
  DFF_X1 \CACHE_MEM_reg[1][58]  ( .D(n10402), .CK(N28803), .Q(n116), .QN(n9149) );
  DFF_X1 \CACHE_MEM_reg[1][57]  ( .D(n10401), .CK(N28803), .Q(n107), .QN(n9165) );
  DFF_X1 \CACHE_MEM_reg[1][56]  ( .D(n10400), .CK(N28803), .Q(n98), .QN(n9181)
         );
  DFF_X1 \CACHE_MEM_reg[1][55]  ( .D(n10399), .CK(N28803), .Q(n89), .QN(n9197)
         );
  DFF_X1 \CACHE_MEM_reg[1][54]  ( .D(n10398), .CK(N28803), .Q(n80), .QN(n9213)
         );
  DFF_X1 \CACHE_MEM_reg[1][53]  ( .D(n10397), .CK(N28803), .Q(n64), .QN(n9229)
         );
  DFF_X1 \CACHE_MEM_reg[1][52]  ( .D(n10396), .CK(N28803), .Q(n61), .QN(n9245)
         );
  DFF_X1 \CACHE_MEM_reg[1][51]  ( .D(n10395), .CK(N28803), .Q(n58), .QN(n9261)
         );
  DFF_X1 \CACHE_MEM_reg[1][50]  ( .D(n10394), .CK(N28803), .Q(n55), .QN(n9277)
         );
  DFF_X1 \CACHE_MEM_reg[1][49]  ( .D(n10393), .CK(N28803), .Q(n52), .QN(n9293)
         );
  DFF_X1 \CACHE_MEM_reg[1][48]  ( .D(n10392), .CK(N28803), .Q(n49), .QN(n9309)
         );
  DFF_X1 \CACHE_MEM_reg[1][47]  ( .D(n10391), .CK(N28803), .Q(n46), .QN(n9325)
         );
  DFF_X1 \CACHE_MEM_reg[1][46]  ( .D(n10390), .CK(N28803), .Q(n43), .QN(n9341)
         );
  DFF_X1 \CACHE_MEM_reg[1][45]  ( .D(n10389), .CK(N28803), .Q(n40), .QN(n9357)
         );
  DFF_X1 \CACHE_MEM_reg[1][44]  ( .D(n10388), .CK(N28803), .Q(n37), .QN(n9373)
         );
  DFF_X1 \CACHE_MEM_reg[1][43]  ( .D(n10387), .CK(N28803), .Q(n34), .QN(n9389)
         );
  DFF_X1 \CACHE_MEM_reg[1][42]  ( .D(n10386), .CK(N28803), .Q(n31), .QN(n9405)
         );
  DFF_X1 \CACHE_MEM_reg[1][41]  ( .D(n10385), .CK(N28803), .Q(n28), .QN(n9421)
         );
  DFF_X1 \CACHE_MEM_reg[1][40]  ( .D(n10384), .CK(N28803), .Q(n25), .QN(n9437)
         );
  DFF_X1 \CACHE_MEM_reg[1][39]  ( .D(n10383), .CK(N28803), .Q(n22), .QN(n9453)
         );
  DFF_X1 \CACHE_MEM_reg[1][38]  ( .D(n10382), .CK(N28803), .Q(n19), .QN(n9469)
         );
  DFF_X1 \CACHE_MEM_reg[1][37]  ( .D(n10381), .CK(N28803), .Q(n16), .QN(n9485)
         );
  DFF_X1 \CACHE_MEM_reg[1][36]  ( .D(n10380), .CK(N28803), .Q(n13), .QN(n9501)
         );
  DFF_X1 \CACHE_MEM_reg[1][35]  ( .D(n10379), .CK(N28803), .Q(n10), .QN(n9517)
         );
  DFF_X1 \CACHE_MEM_reg[1][34]  ( .D(n10378), .CK(N28803), .Q(n7), .QN(n9533)
         );
  DFF_X1 \CACHE_MEM_reg[1][33]  ( .D(n10377), .CK(N28803), .Q(n4), .QN(n9549)
         );
  DFF_X1 \CACHE_MEM_reg[1][32]  ( .D(n10376), .CK(N28803), .Q(n1), .QN(n9565)
         );
  DFF_X1 \CACHE_MEM_reg[1][31]  ( .D(n10375), .CK(N28803), .Q(n2435), .QN(
        n9581) );
  DFF_X1 \CACHE_MEM_reg[1][30]  ( .D(n10374), .CK(N28803), .Q(n2424), .QN(
        n9597) );
  DFF_X1 \CACHE_MEM_reg[1][29]  ( .D(n10373), .CK(N28803), .Q(n2407), .QN(
        n9613) );
  DFF_X1 \CACHE_MEM_reg[1][28]  ( .D(n10372), .CK(N28803), .Q(n2396), .QN(
        n9629) );
  DFF_X1 \CACHE_MEM_reg[1][27]  ( .D(n10371), .CK(N28803), .Q(n2374), .QN(
        n9645) );
  DFF_X1 \CACHE_MEM_reg[1][26]  ( .D(n10370), .CK(N28803), .Q(n2363), .QN(
        n9661) );
  DFF_X1 \CACHE_MEM_reg[1][25]  ( .D(n10369), .CK(N28803), .Q(n2350), .QN(
        n9677) );
  DFF_X1 \CACHE_MEM_reg[1][24]  ( .D(n10368), .CK(N28803), .Q(n2335), .QN(
        n9693) );
  DFF_X1 \CACHE_MEM_reg[1][23]  ( .D(n10367), .CK(N28803), .Q(n2322), .QN(
        n9709) );
  DFF_X1 \CACHE_MEM_reg[1][22]  ( .D(n10366), .CK(N28803), .Q(n2311), .QN(
        n9725) );
  DFF_X1 \CACHE_MEM_reg[1][21]  ( .D(n10365), .CK(N28803), .Q(n2294), .QN(
        n9741) );
  DFF_X1 \CACHE_MEM_reg[1][20]  ( .D(n10364), .CK(N28803), .Q(n2283), .QN(
        n9757) );
  DFF_X1 \CACHE_MEM_reg[1][19]  ( .D(n10363), .CK(N28803), .Q(n2266), .QN(
        n9773) );
  DFF_X1 \CACHE_MEM_reg[1][18]  ( .D(n10362), .CK(N28803), .Q(n2255), .QN(
        n9789) );
  DFF_X1 \CACHE_MEM_reg[1][17]  ( .D(n10361), .CK(N28803), .Q(n2242), .QN(
        n9805) );
  DFF_X1 \CACHE_MEM_reg[1][16]  ( .D(n10360), .CK(N28803), .Q(n2222), .QN(
        n9821) );
  DFF_X1 \CACHE_MEM_reg[1][15]  ( .D(n10359), .CK(N28803), .Q(n2209), .QN(
        n9837) );
  DFF_X1 \CACHE_MEM_reg[1][14]  ( .D(n10358), .CK(N28803), .Q(n2198), .QN(
        n9853) );
  DFF_X1 \CACHE_MEM_reg[1][13]  ( .D(n10357), .CK(N28803), .Q(n2181), .QN(
        n9869) );
  DFF_X1 \CACHE_MEM_reg[1][12]  ( .D(n10356), .CK(N28803), .Q(n2170), .QN(
        n9885) );
  DFF_X1 \CACHE_MEM_reg[1][11]  ( .D(n10355), .CK(N28803), .Q(n2153), .QN(
        n9901) );
  DFF_X1 \CACHE_MEM_reg[1][10]  ( .D(n10354), .CK(N28803), .Q(n2142), .QN(
        n9917) );
  DFF_X1 \CACHE_MEM_reg[1][9]  ( .D(n10353), .CK(N28803), .Q(n2129), .QN(n9933) );
  DFF_X1 \CACHE_MEM_reg[1][8]  ( .D(n10352), .CK(N28803), .Q(n2114), .QN(n9949) );
  DFF_X1 \CACHE_MEM_reg[1][7]  ( .D(n10351), .CK(N28803), .Q(n2101), .QN(n9965) );
  DFF_X1 \CACHE_MEM_reg[1][6]  ( .D(n10350), .CK(N28803), .Q(n2090), .QN(n9981) );
  DFF_X1 \CACHE_MEM_reg[1][5]  ( .D(n10349), .CK(N28803), .Q(n2068), .QN(n9997) );
  DFF_X1 \CACHE_MEM_reg[1][4]  ( .D(n10348), .CK(N28803), .Q(n2057), .QN(
        n10013) );
  DFF_X1 \CACHE_MEM_reg[1][3]  ( .D(n10347), .CK(N28803), .Q(n2040), .QN(
        n10029) );
  DFF_X1 \CACHE_MEM_reg[1][2]  ( .D(n10346), .CK(N28803), .Q(n2029), .QN(
        n10045) );
  DFF_X1 \CACHE_MEM_reg[1][1]  ( .D(n10345), .CK(N28803), .Q(n2016), .QN(
        n10061) );
  DFF_X1 \CACHE_MEM_reg[1][0]  ( .D(n10344), .CK(N28803), .Q(n2001), .QN(
        n10077) );
  DFF_X1 \CACHE_MEM_reg[0][255]  ( .D(n10343), .CK(N28803), .QN(n5993) );
  DFF_X1 \CACHE_MEM_reg[0][254]  ( .D(n10342), .CK(N28803), .QN(n6009) );
  DFF_X1 \CACHE_MEM_reg[0][253]  ( .D(n10341), .CK(N28803), .QN(n6025) );
  DFF_X1 \CACHE_MEM_reg[0][252]  ( .D(n10340), .CK(N28803), .QN(n6041) );
  DFF_X1 \CACHE_MEM_reg[0][251]  ( .D(n10339), .CK(N28803), .QN(n6057) );
  DFF_X1 \CACHE_MEM_reg[0][250]  ( .D(n10338), .CK(N28803), .QN(n6073) );
  DFF_X1 \CACHE_MEM_reg[0][249]  ( .D(n10337), .CK(N28803), .QN(n6089) );
  DFF_X1 \CACHE_MEM_reg[0][248]  ( .D(n10336), .CK(N28803), .QN(n6105) );
  DFF_X1 \CACHE_MEM_reg[0][247]  ( .D(n10335), .CK(N28803), .QN(n6121) );
  DFF_X1 \CACHE_MEM_reg[0][246]  ( .D(n10334), .CK(N28803), .QN(n6137) );
  DFF_X1 \CACHE_MEM_reg[0][245]  ( .D(n10333), .CK(N28803), .QN(n6153) );
  DFF_X1 \CACHE_MEM_reg[0][244]  ( .D(n10332), .CK(N28803), .QN(n6169) );
  DFF_X1 \CACHE_MEM_reg[0][243]  ( .D(n10331), .CK(N28803), .QN(n6185) );
  DFF_X1 \CACHE_MEM_reg[0][242]  ( .D(n10330), .CK(N28803), .QN(n6201) );
  DFF_X1 \CACHE_MEM_reg[0][241]  ( .D(n10329), .CK(N28803), .QN(n6217) );
  DFF_X1 \CACHE_MEM_reg[0][240]  ( .D(n10328), .CK(N28803), .QN(n6233) );
  DFF_X1 \CACHE_MEM_reg[0][239]  ( .D(n10327), .CK(N28803), .QN(n6249) );
  DFF_X1 \CACHE_MEM_reg[0][238]  ( .D(n10326), .CK(N28803), .QN(n6265) );
  DFF_X1 \CACHE_MEM_reg[0][237]  ( .D(n10325), .CK(N28803), .QN(n6281) );
  DFF_X1 \CACHE_MEM_reg[0][236]  ( .D(n10324), .CK(N28803), .QN(n6297) );
  DFF_X1 \CACHE_MEM_reg[0][235]  ( .D(n10323), .CK(N28803), .QN(n6313) );
  DFF_X1 \CACHE_MEM_reg[0][234]  ( .D(n10322), .CK(N28803), .QN(n6329) );
  DFF_X1 \CACHE_MEM_reg[0][233]  ( .D(n10321), .CK(N28803), .QN(n6345) );
  DFF_X1 \CACHE_MEM_reg[0][232]  ( .D(n10320), .CK(N28803), .QN(n6361) );
  DFF_X1 \CACHE_MEM_reg[0][231]  ( .D(n10319), .CK(N28803), .QN(n6377) );
  DFF_X1 \CACHE_MEM_reg[0][230]  ( .D(n10318), .CK(N28803), .QN(n6393) );
  DFF_X1 \CACHE_MEM_reg[0][229]  ( .D(n10317), .CK(N28803), .QN(n6409) );
  DFF_X1 \CACHE_MEM_reg[0][228]  ( .D(n10316), .CK(N28803), .QN(n6425) );
  DFF_X1 \CACHE_MEM_reg[0][227]  ( .D(n10315), .CK(N28803), .QN(n6441) );
  DFF_X1 \CACHE_MEM_reg[0][226]  ( .D(n10314), .CK(N28803), .QN(n6457) );
  DFF_X1 \CACHE_MEM_reg[0][225]  ( .D(n10313), .CK(N28803), .QN(n6473) );
  DFF_X1 \CACHE_MEM_reg[0][224]  ( .D(n10312), .CK(N28803), .QN(n6489) );
  DFF_X1 \CACHE_MEM_reg[0][223]  ( .D(n10311), .CK(N28803), .QN(n6505) );
  DFF_X1 \CACHE_MEM_reg[0][222]  ( .D(n10310), .CK(N28803), .QN(n6521) );
  DFF_X1 \CACHE_MEM_reg[0][221]  ( .D(n10309), .CK(N28803), .QN(n6537) );
  DFF_X1 \CACHE_MEM_reg[0][220]  ( .D(n10308), .CK(N28803), .QN(n6553) );
  DFF_X1 \CACHE_MEM_reg[0][219]  ( .D(n10307), .CK(N28803), .QN(n6569) );
  DFF_X1 \CACHE_MEM_reg[0][218]  ( .D(n10306), .CK(N28803), .QN(n6585) );
  DFF_X1 \CACHE_MEM_reg[0][217]  ( .D(n10305), .CK(N28803), .QN(n6601) );
  DFF_X1 \CACHE_MEM_reg[0][216]  ( .D(n10304), .CK(N28803), .QN(n6617) );
  DFF_X1 \CACHE_MEM_reg[0][215]  ( .D(n10303), .CK(N28803), .QN(n6633) );
  DFF_X1 \CACHE_MEM_reg[0][214]  ( .D(n10302), .CK(N28803), .QN(n6649) );
  DFF_X1 \CACHE_MEM_reg[0][213]  ( .D(n10301), .CK(N28803), .QN(n6665) );
  DFF_X1 \CACHE_MEM_reg[0][212]  ( .D(n10300), .CK(N28803), .QN(n6681) );
  DFF_X1 \CACHE_MEM_reg[0][211]  ( .D(n10299), .CK(N28803), .QN(n6697) );
  DFF_X1 \CACHE_MEM_reg[0][210]  ( .D(n10298), .CK(N28803), .QN(n6713) );
  DFF_X1 \CACHE_MEM_reg[0][209]  ( .D(n10297), .CK(N28803), .QN(n6729) );
  DFF_X1 \CACHE_MEM_reg[0][208]  ( .D(n10296), .CK(N28803), .QN(n6745) );
  DFF_X1 \CACHE_MEM_reg[0][207]  ( .D(n10295), .CK(N28803), .QN(n6761) );
  DFF_X1 \CACHE_MEM_reg[0][206]  ( .D(n10294), .CK(N28803), .QN(n6777) );
  DFF_X1 \CACHE_MEM_reg[0][205]  ( .D(n10293), .CK(N28803), .QN(n6793) );
  DFF_X1 \CACHE_MEM_reg[0][204]  ( .D(n10292), .CK(N28803), .QN(n6809) );
  DFF_X1 \CACHE_MEM_reg[0][203]  ( .D(n10291), .CK(N28803), .QN(n6825) );
  DFF_X1 \CACHE_MEM_reg[0][202]  ( .D(n10290), .CK(N28803), .QN(n6841) );
  DFF_X1 \CACHE_MEM_reg[0][201]  ( .D(n10289), .CK(N28803), .QN(n6857) );
  DFF_X1 \CACHE_MEM_reg[0][200]  ( .D(n10288), .CK(N28803), .QN(n6873) );
  DFF_X1 \CACHE_MEM_reg[0][199]  ( .D(n10287), .CK(N28803), .QN(n6889) );
  DFF_X1 \CACHE_MEM_reg[0][198]  ( .D(n10286), .CK(N28803), .QN(n6905) );
  DFF_X1 \CACHE_MEM_reg[0][197]  ( .D(n10285), .CK(N28803), .QN(n6921) );
  DFF_X1 \CACHE_MEM_reg[0][196]  ( .D(n10284), .CK(N28803), .QN(n6937) );
  DFF_X1 \CACHE_MEM_reg[0][195]  ( .D(n10283), .CK(N28803), .QN(n6953) );
  DFF_X1 \CACHE_MEM_reg[0][194]  ( .D(n10282), .CK(N28803), .QN(n6969) );
  DFF_X1 \CACHE_MEM_reg[0][193]  ( .D(n10281), .CK(N28803), .QN(n6985) );
  DFF_X1 \CACHE_MEM_reg[0][192]  ( .D(n10280), .CK(N28803), .QN(n7001) );
  DFF_X1 \CACHE_MEM_reg[0][191]  ( .D(n10279), .CK(N28803), .QN(n7017) );
  DFF_X1 \CACHE_MEM_reg[0][190]  ( .D(n10278), .CK(N28803), .QN(n7033) );
  DFF_X1 \CACHE_MEM_reg[0][189]  ( .D(n10277), .CK(N28803), .QN(n7049) );
  DFF_X1 \CACHE_MEM_reg[0][188]  ( .D(n10276), .CK(N28803), .QN(n7065) );
  DFF_X1 \CACHE_MEM_reg[0][187]  ( .D(n10275), .CK(N28803), .QN(n7081) );
  DFF_X1 \CACHE_MEM_reg[0][186]  ( .D(n10274), .CK(N28803), .QN(n7097) );
  DFF_X1 \CACHE_MEM_reg[0][185]  ( .D(n10273), .CK(N28803), .QN(n7113) );
  DFF_X1 \CACHE_MEM_reg[0][184]  ( .D(n10272), .CK(N28803), .QN(n7129) );
  DFF_X1 \CACHE_MEM_reg[0][183]  ( .D(n10271), .CK(N28803), .QN(n7145) );
  DFF_X1 \CACHE_MEM_reg[0][182]  ( .D(n10270), .CK(N28803), .QN(n7161) );
  DFF_X1 \CACHE_MEM_reg[0][181]  ( .D(n10269), .CK(N28803), .QN(n7177) );
  DFF_X1 \CACHE_MEM_reg[0][180]  ( .D(n10268), .CK(N28803), .QN(n7193) );
  DFF_X1 \CACHE_MEM_reg[0][179]  ( .D(n10267), .CK(N28803), .QN(n7209) );
  DFF_X1 \CACHE_MEM_reg[0][178]  ( .D(n10266), .CK(N28803), .QN(n7225) );
  DFF_X1 \CACHE_MEM_reg[0][177]  ( .D(n10265), .CK(N28803), .QN(n7241) );
  DFF_X1 \CACHE_MEM_reg[0][176]  ( .D(n10264), .CK(N28803), .QN(n7257) );
  DFF_X1 \CACHE_MEM_reg[0][175]  ( .D(n10263), .CK(N28803), .QN(n7273) );
  DFF_X1 \CACHE_MEM_reg[0][174]  ( .D(n10262), .CK(N28803), .QN(n7289) );
  DFF_X1 \CACHE_MEM_reg[0][173]  ( .D(n10261), .CK(N28803), .QN(n7305) );
  DFF_X1 \CACHE_MEM_reg[0][172]  ( .D(n10260), .CK(N28803), .QN(n7321) );
  DFF_X1 \CACHE_MEM_reg[0][171]  ( .D(n10259), .CK(N28803), .QN(n7337) );
  DFF_X1 \CACHE_MEM_reg[0][170]  ( .D(n10258), .CK(N28803), .QN(n7353) );
  DFF_X1 \CACHE_MEM_reg[0][169]  ( .D(n10257), .CK(N28803), .QN(n7369) );
  DFF_X1 \CACHE_MEM_reg[0][168]  ( .D(n10256), .CK(N28803), .QN(n7385) );
  DFF_X1 \CACHE_MEM_reg[0][167]  ( .D(n10255), .CK(N28803), .QN(n7401) );
  DFF_X1 \CACHE_MEM_reg[0][166]  ( .D(n10254), .CK(N28803), .QN(n7417) );
  DFF_X1 \CACHE_MEM_reg[0][165]  ( .D(n10253), .CK(N28803), .QN(n7433) );
  DFF_X1 \CACHE_MEM_reg[0][164]  ( .D(n10252), .CK(N28803), .QN(n7449) );
  DFF_X1 \CACHE_MEM_reg[0][163]  ( .D(n10251), .CK(N28803), .QN(n7465) );
  DFF_X1 \CACHE_MEM_reg[0][162]  ( .D(n10250), .CK(N28803), .QN(n7481) );
  DFF_X1 \CACHE_MEM_reg[0][161]  ( .D(n10249), .CK(N28803), .QN(n7497) );
  DFF_X1 \CACHE_MEM_reg[0][160]  ( .D(n10248), .CK(N28803), .QN(n7513) );
  DFF_X1 \CACHE_MEM_reg[0][159]  ( .D(n10247), .CK(N28803), .QN(n7529) );
  DFF_X1 \CACHE_MEM_reg[0][158]  ( .D(n10246), .CK(N28803), .QN(n7545) );
  DFF_X1 \CACHE_MEM_reg[0][157]  ( .D(n10245), .CK(N28803), .QN(n7561) );
  DFF_X1 \CACHE_MEM_reg[0][156]  ( .D(n10244), .CK(N28803), .QN(n7577) );
  DFF_X1 \CACHE_MEM_reg[0][155]  ( .D(n10243), .CK(N28803), .QN(n7593) );
  DFF_X1 \CACHE_MEM_reg[0][154]  ( .D(n10242), .CK(N28803), .QN(n7609) );
  DFF_X1 \CACHE_MEM_reg[0][153]  ( .D(n10241), .CK(N28803), .QN(n7625) );
  DFF_X1 \CACHE_MEM_reg[0][152]  ( .D(n10240), .CK(N28803), .QN(n7641) );
  DFF_X1 \CACHE_MEM_reg[0][151]  ( .D(n10239), .CK(N28803), .QN(n7657) );
  DFF_X1 \CACHE_MEM_reg[0][150]  ( .D(n10238), .CK(N28803), .QN(n7673) );
  DFF_X1 \CACHE_MEM_reg[0][149]  ( .D(n10237), .CK(N28803), .QN(n7689) );
  DFF_X1 \CACHE_MEM_reg[0][148]  ( .D(n10236), .CK(N28803), .QN(n7705) );
  DFF_X1 \CACHE_MEM_reg[0][147]  ( .D(n10235), .CK(N28803), .QN(n7721) );
  DFF_X1 \CACHE_MEM_reg[0][146]  ( .D(n10234), .CK(N28803), .QN(n7737) );
  DFF_X1 \CACHE_MEM_reg[0][145]  ( .D(n10233), .CK(N28803), .QN(n7753) );
  DFF_X1 \CACHE_MEM_reg[0][144]  ( .D(n10232), .CK(N28803), .QN(n7769) );
  DFF_X1 \CACHE_MEM_reg[0][143]  ( .D(n10231), .CK(N28803), .QN(n7785) );
  DFF_X1 \CACHE_MEM_reg[0][142]  ( .D(n10230), .CK(N28803), .QN(n7801) );
  DFF_X1 \CACHE_MEM_reg[0][141]  ( .D(n10229), .CK(N28803), .QN(n7817) );
  DFF_X1 \CACHE_MEM_reg[0][140]  ( .D(n10228), .CK(N28803), .QN(n7833) );
  DFF_X1 \CACHE_MEM_reg[0][139]  ( .D(n10227), .CK(N28803), .QN(n7849) );
  DFF_X1 \CACHE_MEM_reg[0][138]  ( .D(n10226), .CK(N28803), .QN(n7865) );
  DFF_X1 \CACHE_MEM_reg[0][137]  ( .D(n10225), .CK(N28803), .QN(n7881) );
  DFF_X1 \CACHE_MEM_reg[0][136]  ( .D(n10224), .CK(N28803), .QN(n7897) );
  DFF_X1 \CACHE_MEM_reg[0][135]  ( .D(n10223), .CK(N28803), .QN(n7913) );
  DFF_X1 \CACHE_MEM_reg[0][134]  ( .D(n10222), .CK(N28803), .QN(n7929) );
  DFF_X1 \CACHE_MEM_reg[0][133]  ( .D(n10221), .CK(N28803), .QN(n7945) );
  DFF_X1 \CACHE_MEM_reg[0][132]  ( .D(n10220), .CK(N28803), .QN(n7961) );
  DFF_X1 \CACHE_MEM_reg[0][131]  ( .D(n10219), .CK(N28803), .QN(n7977) );
  DFF_X1 \CACHE_MEM_reg[0][130]  ( .D(n10218), .CK(N28803), .QN(n7993) );
  DFF_X1 \CACHE_MEM_reg[0][129]  ( .D(n10217), .CK(N28803), .QN(n8009) );
  DFF_X1 \CACHE_MEM_reg[0][128]  ( .D(n10216), .CK(N28803), .QN(n8025) );
  DFF_X1 \CACHE_MEM_reg[0][127]  ( .D(n10215), .CK(N28803), .QN(n8041) );
  DFF_X1 \CACHE_MEM_reg[0][126]  ( .D(n10214), .CK(N28803), .QN(n8057) );
  DFF_X1 \CACHE_MEM_reg[0][125]  ( .D(n10213), .CK(N28803), .QN(n8073) );
  DFF_X1 \CACHE_MEM_reg[0][124]  ( .D(n10212), .CK(N28803), .QN(n8089) );
  DFF_X1 \CACHE_MEM_reg[0][123]  ( .D(n10211), .CK(N28803), .QN(n8105) );
  DFF_X1 \CACHE_MEM_reg[0][122]  ( .D(n10210), .CK(N28803), .QN(n8121) );
  DFF_X1 \CACHE_MEM_reg[0][121]  ( .D(n10209), .CK(N28803), .QN(n8137) );
  DFF_X1 \CACHE_MEM_reg[0][120]  ( .D(n10208), .CK(N28803), .QN(n8153) );
  DFF_X1 \CACHE_MEM_reg[0][119]  ( .D(n10207), .CK(N28803), .QN(n8169) );
  DFF_X1 \CACHE_MEM_reg[0][118]  ( .D(n10206), .CK(N28803), .QN(n8185) );
  DFF_X1 \CACHE_MEM_reg[0][117]  ( .D(n10205), .CK(N28803), .QN(n8201) );
  DFF_X1 \CACHE_MEM_reg[0][116]  ( .D(n10204), .CK(N28803), .QN(n8217) );
  DFF_X1 \CACHE_MEM_reg[0][115]  ( .D(n10203), .CK(N28803), .QN(n8233) );
  DFF_X1 \CACHE_MEM_reg[0][114]  ( .D(n10202), .CK(N28803), .QN(n8249) );
  DFF_X1 \CACHE_MEM_reg[0][113]  ( .D(n10201), .CK(N28803), .QN(n8265) );
  DFF_X1 \CACHE_MEM_reg[0][112]  ( .D(n10200), .CK(N28803), .QN(n8281) );
  DFF_X1 \CACHE_MEM_reg[0][111]  ( .D(n10199), .CK(N28803), .QN(n8297) );
  DFF_X1 \CACHE_MEM_reg[0][110]  ( .D(n10198), .CK(N28803), .QN(n8313) );
  DFF_X1 \CACHE_MEM_reg[0][109]  ( .D(n10197), .CK(N28803), .QN(n8329) );
  DFF_X1 \CACHE_MEM_reg[0][108]  ( .D(n10196), .CK(N28803), .QN(n8345) );
  DFF_X1 \CACHE_MEM_reg[0][107]  ( .D(n10195), .CK(N28803), .QN(n8361) );
  DFF_X1 \CACHE_MEM_reg[0][106]  ( .D(n10194), .CK(N28803), .QN(n8377) );
  DFF_X1 \CACHE_MEM_reg[0][105]  ( .D(n10193), .CK(N28803), .QN(n8393) );
  DFF_X1 \CACHE_MEM_reg[0][104]  ( .D(n10192), .CK(N28803), .QN(n8409) );
  DFF_X1 \CACHE_MEM_reg[0][103]  ( .D(n10191), .CK(N28803), .QN(n8425) );
  DFF_X1 \CACHE_MEM_reg[0][102]  ( .D(n10190), .CK(N28803), .QN(n8441) );
  DFF_X1 \CACHE_MEM_reg[0][101]  ( .D(n10189), .CK(N28803), .QN(n8457) );
  DFF_X1 \CACHE_MEM_reg[0][100]  ( .D(n10188), .CK(N28803), .QN(n8473) );
  DFF_X1 \CACHE_MEM_reg[0][99]  ( .D(n10187), .CK(N28803), .QN(n8489) );
  DFF_X1 \CACHE_MEM_reg[0][98]  ( .D(n10186), .CK(N28803), .QN(n8505) );
  DFF_X1 \CACHE_MEM_reg[0][97]  ( .D(n10185), .CK(N28803), .QN(n8521) );
  DFF_X1 \CACHE_MEM_reg[0][96]  ( .D(n10184), .CK(N28803), .QN(n8537) );
  DFF_X1 \CACHE_MEM_reg[0][95]  ( .D(n10183), .CK(N28803), .QN(n8553) );
  DFF_X1 \CACHE_MEM_reg[0][94]  ( .D(n10182), .CK(N28803), .QN(n8569) );
  DFF_X1 \CACHE_MEM_reg[0][93]  ( .D(n10181), .CK(N28803), .QN(n8585) );
  DFF_X1 \CACHE_MEM_reg[0][92]  ( .D(n10180), .CK(N28803), .QN(n8601) );
  DFF_X1 \CACHE_MEM_reg[0][91]  ( .D(n10179), .CK(N28803), .QN(n8617) );
  DFF_X1 \CACHE_MEM_reg[0][90]  ( .D(n10178), .CK(N28803), .QN(n8633) );
  DFF_X1 \CACHE_MEM_reg[0][89]  ( .D(n10177), .CK(N28803), .QN(n8649) );
  DFF_X1 \CACHE_MEM_reg[0][88]  ( .D(n10176), .CK(N28803), .QN(n8665) );
  DFF_X1 \CACHE_MEM_reg[0][87]  ( .D(n10175), .CK(N28803), .QN(n8681) );
  DFF_X1 \CACHE_MEM_reg[0][86]  ( .D(n10174), .CK(N28803), .QN(n8697) );
  DFF_X1 \CACHE_MEM_reg[0][85]  ( .D(n10173), .CK(N28803), .QN(n8713) );
  DFF_X1 \CACHE_MEM_reg[0][84]  ( .D(n10172), .CK(N28803), .QN(n8729) );
  DFF_X1 \CACHE_MEM_reg[0][83]  ( .D(n10171), .CK(N28803), .QN(n8745) );
  DFF_X1 \CACHE_MEM_reg[0][82]  ( .D(n10170), .CK(N28803), .QN(n8761) );
  DFF_X1 \CACHE_MEM_reg[0][81]  ( .D(n10169), .CK(N28803), .QN(n8777) );
  DFF_X1 \CACHE_MEM_reg[0][80]  ( .D(n10168), .CK(N28803), .QN(n8793) );
  DFF_X1 \CACHE_MEM_reg[0][79]  ( .D(n10167), .CK(N28803), .QN(n8809) );
  DFF_X1 \CACHE_MEM_reg[0][78]  ( .D(n10166), .CK(N28803), .QN(n8825) );
  DFF_X1 \CACHE_MEM_reg[0][77]  ( .D(n10165), .CK(N28803), .QN(n8841) );
  DFF_X1 \CACHE_MEM_reg[0][76]  ( .D(n10164), .CK(N28803), .QN(n8857) );
  DFF_X1 \CACHE_MEM_reg[0][75]  ( .D(n10163), .CK(N28803), .QN(n8873) );
  DFF_X1 \CACHE_MEM_reg[0][74]  ( .D(n10162), .CK(N28803), .QN(n8889) );
  DFF_X1 \CACHE_MEM_reg[0][73]  ( .D(n10161), .CK(N28803), .QN(n8905) );
  DFF_X1 \CACHE_MEM_reg[0][72]  ( .D(n10160), .CK(N28803), .QN(n8921) );
  DFF_X1 \CACHE_MEM_reg[0][71]  ( .D(n10159), .CK(N28803), .QN(n8937) );
  DFF_X1 \CACHE_MEM_reg[0][70]  ( .D(n10158), .CK(N28803), .QN(n8953) );
  DFF_X1 \CACHE_MEM_reg[0][69]  ( .D(n10157), .CK(N28803), .QN(n8969) );
  DFF_X1 \CACHE_MEM_reg[0][68]  ( .D(n10156), .CK(N28803), .QN(n8985) );
  DFF_X1 \CACHE_MEM_reg[0][67]  ( .D(n10155), .CK(N28803), .QN(n9001) );
  DFF_X1 \CACHE_MEM_reg[0][66]  ( .D(n10154), .CK(N28803), .QN(n9017) );
  DFF_X1 \CACHE_MEM_reg[0][65]  ( .D(n10153), .CK(N28803), .QN(n9033) );
  DFF_X1 \CACHE_MEM_reg[0][64]  ( .D(n10152), .CK(N28803), .QN(n9049) );
  DFF_X1 \CACHE_MEM_reg[0][63]  ( .D(n10151), .CK(N28803), .QN(n9065) );
  DFF_X1 \CACHE_MEM_reg[0][62]  ( .D(n10150), .CK(N28803), .QN(n9081) );
  DFF_X1 \CACHE_MEM_reg[0][61]  ( .D(n10149), .CK(N28803), .QN(n9097) );
  DFF_X1 \CACHE_MEM_reg[0][60]  ( .D(n10148), .CK(N28803), .QN(n9113) );
  DFF_X1 \CACHE_MEM_reg[0][59]  ( .D(n10147), .CK(N28803), .QN(n9129) );
  DFF_X1 \CACHE_MEM_reg[0][58]  ( .D(n10146), .CK(N28803), .QN(n9145) );
  DFF_X1 \CACHE_MEM_reg[0][57]  ( .D(n10145), .CK(N28803), .QN(n9161) );
  DFF_X1 \CACHE_MEM_reg[0][56]  ( .D(n10144), .CK(N28803), .QN(n9177) );
  DFF_X1 \CACHE_MEM_reg[0][55]  ( .D(n10143), .CK(N28803), .QN(n9193) );
  DFF_X1 \CACHE_MEM_reg[0][54]  ( .D(n10142), .CK(N28803), .QN(n9209) );
  DFF_X1 \CACHE_MEM_reg[0][53]  ( .D(n10141), .CK(N28803), .QN(n9225) );
  DFF_X1 \CACHE_MEM_reg[0][52]  ( .D(n10140), .CK(N28803), .QN(n9241) );
  DFF_X1 \CACHE_MEM_reg[0][51]  ( .D(n10139), .CK(N28803), .QN(n9257) );
  DFF_X1 \CACHE_MEM_reg[0][50]  ( .D(n10138), .CK(N28803), .QN(n9273) );
  DFF_X1 \CACHE_MEM_reg[0][49]  ( .D(n10137), .CK(N28803), .QN(n9289) );
  DFF_X1 \CACHE_MEM_reg[0][48]  ( .D(n10136), .CK(N28803), .QN(n9305) );
  DFF_X1 \CACHE_MEM_reg[0][47]  ( .D(n10135), .CK(N28803), .QN(n9321) );
  DFF_X1 \CACHE_MEM_reg[0][46]  ( .D(n10134), .CK(N28803), .QN(n9337) );
  DFF_X1 \CACHE_MEM_reg[0][45]  ( .D(n10133), .CK(N28803), .QN(n9353) );
  DFF_X1 \CACHE_MEM_reg[0][44]  ( .D(n10132), .CK(N28803), .QN(n9369) );
  DFF_X1 \CACHE_MEM_reg[0][43]  ( .D(n10131), .CK(N28803), .QN(n9385) );
  DFF_X1 \CACHE_MEM_reg[0][42]  ( .D(n10130), .CK(N28803), .QN(n9401) );
  DFF_X1 \CACHE_MEM_reg[0][41]  ( .D(n10129), .CK(N28803), .QN(n9417) );
  DFF_X1 \CACHE_MEM_reg[0][40]  ( .D(n10128), .CK(N28803), .QN(n9433) );
  DFF_X1 \CACHE_MEM_reg[0][39]  ( .D(n10127), .CK(N28803), .QN(n9449) );
  DFF_X1 \CACHE_MEM_reg[0][38]  ( .D(n10126), .CK(N28803), .QN(n9465) );
  DFF_X1 \CACHE_MEM_reg[0][37]  ( .D(n10125), .CK(N28803), .QN(n9481) );
  DFF_X1 \CACHE_MEM_reg[0][36]  ( .D(n10124), .CK(N28803), .QN(n9497) );
  DFF_X1 \CACHE_MEM_reg[0][35]  ( .D(n10123), .CK(N28803), .QN(n9513) );
  DFF_X1 \CACHE_MEM_reg[0][34]  ( .D(n10122), .CK(N28803), .QN(n9529) );
  DFF_X1 \CACHE_MEM_reg[0][33]  ( .D(n10121), .CK(N28803), .QN(n9545) );
  DFF_X1 \CACHE_MEM_reg[0][32]  ( .D(n10120), .CK(N28803), .QN(n9561) );
  DFF_X1 \CACHE_MEM_reg[0][31]  ( .D(n10119), .CK(N28803), .QN(n9577) );
  DFF_X1 \CACHE_MEM_reg[0][30]  ( .D(n10118), .CK(N28803), .QN(n9593) );
  DFF_X1 \CACHE_MEM_reg[0][29]  ( .D(n10117), .CK(N28803), .QN(n9609) );
  DFF_X1 \CACHE_MEM_reg[0][28]  ( .D(n10116), .CK(N28803), .QN(n9625) );
  DFF_X1 \CACHE_MEM_reg[0][27]  ( .D(n10115), .CK(N28803), .QN(n9641) );
  DFF_X1 \CACHE_MEM_reg[0][26]  ( .D(n10114), .CK(N28803), .QN(n9657) );
  DFF_X1 \CACHE_MEM_reg[0][25]  ( .D(n10113), .CK(N28803), .QN(n9673) );
  DFF_X1 \CACHE_MEM_reg[0][24]  ( .D(n10112), .CK(N28803), .QN(n9689) );
  DFF_X1 \CACHE_MEM_reg[0][23]  ( .D(n10111), .CK(N28803), .QN(n9705) );
  DFF_X1 \CACHE_MEM_reg[0][22]  ( .D(n10110), .CK(N28803), .QN(n9721) );
  DFF_X1 \CACHE_MEM_reg[0][21]  ( .D(n10109), .CK(N28803), .QN(n9737) );
  DFF_X1 \CACHE_MEM_reg[0][20]  ( .D(n10108), .CK(N28803), .QN(n9753) );
  DFF_X1 \CACHE_MEM_reg[0][19]  ( .D(n10107), .CK(N28803), .QN(n9769) );
  DFF_X1 \CACHE_MEM_reg[0][18]  ( .D(n10106), .CK(N28803), .QN(n9785) );
  DFF_X1 \CACHE_MEM_reg[0][17]  ( .D(n10105), .CK(N28803), .QN(n9801) );
  DFF_X1 \CACHE_MEM_reg[0][16]  ( .D(n10104), .CK(N28803), .QN(n9817) );
  DFF_X1 \CACHE_MEM_reg[0][15]  ( .D(n10103), .CK(N28803), .QN(n9833) );
  DFF_X1 \CACHE_MEM_reg[0][14]  ( .D(n10102), .CK(N28803), .QN(n9849) );
  DFF_X1 \CACHE_MEM_reg[0][13]  ( .D(n10101), .CK(N28803), .QN(n9865) );
  DFF_X1 \CACHE_MEM_reg[0][12]  ( .D(n10100), .CK(N28803), .QN(n9881) );
  DFF_X1 \CACHE_MEM_reg[0][11]  ( .D(n10099), .CK(N28803), .QN(n9897) );
  DFF_X1 \CACHE_MEM_reg[0][10]  ( .D(n10098), .CK(N28803), .QN(n9913) );
  DFF_X1 \CACHE_MEM_reg[0][9]  ( .D(n10097), .CK(N28803), .QN(n9929) );
  DFF_X1 \CACHE_MEM_reg[0][8]  ( .D(n10096), .CK(N28803), .QN(n9945) );
  DFF_X1 \CACHE_MEM_reg[0][7]  ( .D(n10095), .CK(N28803), .QN(n9961) );
  DFF_X1 \CACHE_MEM_reg[0][6]  ( .D(n10094), .CK(N28803), .QN(n9977) );
  DFF_X1 \CACHE_MEM_reg[0][5]  ( .D(n10093), .CK(N28803), .QN(n9993) );
  DFF_X1 \CACHE_MEM_reg[0][4]  ( .D(n10092), .CK(N28803), .QN(n10009) );
  DFF_X1 \CACHE_MEM_reg[0][3]  ( .D(n10091), .CK(N28803), .QN(n10025) );
  DFF_X1 \CACHE_MEM_reg[0][2]  ( .D(n10090), .CK(N28803), .QN(n10041) );
  DFF_X1 \CACHE_MEM_reg[0][1]  ( .D(n10089), .CK(N28803), .QN(n10057) );
  DFF_X1 \CACHE_MEM_reg[0][0]  ( .D(n10088), .CK(N28803), .QN(n10073) );
  NAND2_X1 U5184 ( .A1(n14978), .A2(n1169), .ZN(n14185) );
  NAND2_X1 U5336 ( .A1(n14976), .A2(n1334), .ZN(n14188) );
  NAND2_X1 U5488 ( .A1(n14976), .A2(n1483), .ZN(n14191) );
  NAND2_X1 U5640 ( .A1(n14976), .A2(n1632), .ZN(n14194) );
  NAND2_X1 U5792 ( .A1(n14976), .A2(n1781), .ZN(n14197) );
  NAND2_X1 U5944 ( .A1(n14977), .A2(n1930), .ZN(n14200) );
  NAND2_X1 U6096 ( .A1(n14977), .A2(n2079), .ZN(n14203) );
  NAND2_X1 U6248 ( .A1(n14977), .A2(n2228), .ZN(n14206) );
  NAND2_X1 U6400 ( .A1(n14977), .A2(n2377), .ZN(n14209) );
  NAND2_X1 U6552 ( .A1(n14977), .A2(n2526), .ZN(n14212) );
  NAND2_X1 U6704 ( .A1(n14977), .A2(n2675), .ZN(n14215) );
  NAND2_X1 U6856 ( .A1(n14977), .A2(n2824), .ZN(n14218) );
  NAND2_X1 U7008 ( .A1(n14978), .A2(n2973), .ZN(n14221) );
  NAND2_X1 U7160 ( .A1(n14978), .A2(n3122), .ZN(n14224) );
  NAND2_X1 U7312 ( .A1(n14978), .A2(n3271), .ZN(n14227) );
  NAND2_X1 U7464 ( .A1(n14978), .A2(n3420), .ZN(n14230) );
  NAND2_X1 U7616 ( .A1(n14978), .A2(n3569), .ZN(n14233) );
  NAND2_X1 U7768 ( .A1(n14978), .A2(n3718), .ZN(n14236) );
  NAND2_X1 U7920 ( .A1(n14979), .A2(n3867), .ZN(n14239) );
  NAND2_X1 U8072 ( .A1(n14979), .A2(n4016), .ZN(n14242) );
  NAND2_X1 U8224 ( .A1(n14979), .A2(n4165), .ZN(n14245) );
  NAND2_X1 U8376 ( .A1(n14979), .A2(n4314), .ZN(n14248) );
  NAND2_X1 U8528 ( .A1(n14979), .A2(n4463), .ZN(n14251) );
  NAND2_X1 U8680 ( .A1(n14979), .A2(n4612), .ZN(n14254) );
  NAND2_X1 U8832 ( .A1(n14979), .A2(n4761), .ZN(n14257) );
  NAND2_X1 U8984 ( .A1(n14980), .A2(n4910), .ZN(n14260) );
  NAND2_X1 U9136 ( .A1(n14980), .A2(n5059), .ZN(n14263) );
  NAND2_X1 U9288 ( .A1(n14980), .A2(n5208), .ZN(n14266) );
  NAND2_X1 U9440 ( .A1(n14980), .A2(n5357), .ZN(n14269) );
  NAND2_X1 U9592 ( .A1(n14980), .A2(n5506), .ZN(n14272) );
  NAND2_X1 U9744 ( .A1(n14980), .A2(n5655), .ZN(n14275) );
  NAND2_X1 U9896 ( .A1(n14975), .A2(n5804), .ZN(n14278) );
  NAND2_X1 U9902 ( .A1(n1125), .A2(n14987), .ZN(n1180) );
  NAND2_X1 U9912 ( .A1(n1107), .A2(n14987), .ZN(n1189) );
  NAND2_X1 U9922 ( .A1(n1161), .A2(n14987), .ZN(n1198) );
  NAND2_X1 U9932 ( .A1(n1143), .A2(n14987), .ZN(n1207) );
  NAND2_X1 U9943 ( .A1(n1116), .A2(n14987), .ZN(n1220) );
  NAND2_X1 U9953 ( .A1(n1094), .A2(n14987), .ZN(n1229) );
  NAND2_X1 U9963 ( .A1(n1152), .A2(n14987), .ZN(n1238) );
  NAND2_X1 U9973 ( .A1(n1134), .A2(n14987), .ZN(n1247) );
  NAND2_X1 U9985 ( .A1(n14985), .A2(n1125), .ZN(n1260) );
  NAND2_X1 U9996 ( .A1(n14985), .A2(n1107), .ZN(n1269) );
  NAND2_X1 U10007 ( .A1(n14985), .A2(n1161), .ZN(n1278) );
  NAND2_X1 U10018 ( .A1(n14985), .A2(n1143), .ZN(n1287) );
  NAND2_X1 U10030 ( .A1(n14985), .A2(n1116), .ZN(n1300) );
  NAND2_X1 U10041 ( .A1(n14985), .A2(n1094), .ZN(n1309) );
  NAND2_X1 U10052 ( .A1(n14986), .A2(n1152), .ZN(n1318) );
  NAND2_X1 U10063 ( .A1(n14986), .A2(n1134), .ZN(n1327) );
  NAND2_X1 U10069 ( .A1(ADDR[2]), .A2(n5952), .ZN(n501) );
  NAND2_X1 U10070 ( .A1(n5953), .A2(n14982), .ZN(n959) );
  DFFRS_X2 \DATA_OUT_reg[31]  ( .D(n14279), .CK(N28803), .RN(n14277), .SN(
        n14278), .Q(DATA_OUT[31]), .QN(n5991) );
  DFFRS_X2 \DATA_OUT_reg[30]  ( .D(n14276), .CK(N28803), .RN(n14274), .SN(
        n14275), .Q(DATA_OUT[30]), .QN(n5990) );
  DFFRS_X2 \DATA_OUT_reg[29]  ( .D(n14273), .CK(N28803), .RN(n14271), .SN(
        n14272), .Q(DATA_OUT[29]), .QN(n5989) );
  DFFRS_X2 \DATA_OUT_reg[28]  ( .D(n14270), .CK(N28803), .RN(n14268), .SN(
        n14269), .Q(DATA_OUT[28]), .QN(n5988) );
  DFFRS_X2 \DATA_OUT_reg[27]  ( .D(n14267), .CK(N28803), .RN(n14265), .SN(
        n14266), .Q(DATA_OUT[27]), .QN(n5987) );
  DFFRS_X2 \DATA_OUT_reg[26]  ( .D(n14264), .CK(N28803), .RN(n14262), .SN(
        n14263), .Q(DATA_OUT[26]), .QN(n5986) );
  DFFRS_X2 \DATA_OUT_reg[25]  ( .D(n14261), .CK(N28803), .RN(n14259), .SN(
        n14260), .Q(DATA_OUT[25]), .QN(n5985) );
  DFFRS_X2 \DATA_OUT_reg[24]  ( .D(n14258), .CK(N28803), .RN(n14256), .SN(
        n14257), .Q(DATA_OUT[24]), .QN(n5984) );
  DFFRS_X2 \DATA_OUT_reg[23]  ( .D(n14255), .CK(N28803), .RN(n14253), .SN(
        n14254), .Q(DATA_OUT[23]), .QN(n5983) );
  DFFRS_X2 \DATA_OUT_reg[22]  ( .D(n14252), .CK(N28803), .RN(n14250), .SN(
        n14251), .Q(DATA_OUT[22]), .QN(n5982) );
  DFFRS_X2 \DATA_OUT_reg[21]  ( .D(n14249), .CK(N28803), .RN(n14247), .SN(
        n14248), .Q(DATA_OUT[21]), .QN(n5981) );
  DFFRS_X2 \DATA_OUT_reg[20]  ( .D(n14246), .CK(N28803), .RN(n14244), .SN(
        n14245), .Q(DATA_OUT[20]), .QN(n5980) );
  DFFRS_X2 \DATA_OUT_reg[19]  ( .D(n14243), .CK(N28803), .RN(n14241), .SN(
        n14242), .Q(DATA_OUT[19]), .QN(n5979) );
  DFFRS_X2 \DATA_OUT_reg[18]  ( .D(n14240), .CK(N28803), .RN(n14238), .SN(
        n14239), .Q(DATA_OUT[18]), .QN(n5978) );
  DFFRS_X2 \DATA_OUT_reg[17]  ( .D(n14237), .CK(N28803), .RN(n14235), .SN(
        n14236), .Q(DATA_OUT[17]), .QN(n5977) );
  DFFRS_X2 \DATA_OUT_reg[16]  ( .D(n14234), .CK(N28803), .RN(n14232), .SN(
        n14233), .Q(DATA_OUT[16]), .QN(n5976) );
  DFFRS_X2 \DATA_OUT_reg[15]  ( .D(n14231), .CK(N28803), .RN(n14229), .SN(
        n14230), .Q(DATA_OUT[15]), .QN(n5975) );
  DFFRS_X2 \DATA_OUT_reg[14]  ( .D(n14228), .CK(N28803), .RN(n14226), .SN(
        n14227), .Q(DATA_OUT[14]), .QN(n5974) );
  DFFRS_X2 \DATA_OUT_reg[13]  ( .D(n14225), .CK(N28803), .RN(n14223), .SN(
        n14224), .Q(DATA_OUT[13]), .QN(n5973) );
  DFFRS_X2 \DATA_OUT_reg[12]  ( .D(n14222), .CK(N28803), .RN(n14220), .SN(
        n14221), .Q(DATA_OUT[12]), .QN(n5972) );
  DFFRS_X2 \DATA_OUT_reg[11]  ( .D(n14219), .CK(N28803), .RN(n14217), .SN(
        n14218), .Q(DATA_OUT[11]), .QN(n5971) );
  DFFRS_X2 \DATA_OUT_reg[10]  ( .D(n14216), .CK(N28803), .RN(n14214), .SN(
        n14215), .Q(DATA_OUT[10]), .QN(n5970) );
  DFFRS_X2 \DATA_OUT_reg[9]  ( .D(n14213), .CK(N28803), .RN(n14211), .SN(
        n14212), .Q(DATA_OUT[9]), .QN(n5969) );
  DFFRS_X2 \DATA_OUT_reg[8]  ( .D(n14210), .CK(N28803), .RN(n14208), .SN(
        n14209), .Q(DATA_OUT[8]), .QN(n5968) );
  DFFRS_X2 \DATA_OUT_reg[7]  ( .D(n14207), .CK(N28803), .RN(n14205), .SN(
        n14206), .Q(DATA_OUT[7]), .QN(n5967) );
  DFFRS_X2 \DATA_OUT_reg[6]  ( .D(n14204), .CK(N28803), .RN(n14202), .SN(
        n14203), .Q(DATA_OUT[6]), .QN(n5966) );
  DFFRS_X2 \DATA_OUT_reg[5]  ( .D(n14201), .CK(N28803), .RN(n14199), .SN(
        n14200), .Q(DATA_OUT[5]), .QN(n5965) );
  DFFRS_X2 \DATA_OUT_reg[4]  ( .D(n14198), .CK(N28803), .RN(n14196), .SN(
        n14197), .Q(DATA_OUT[4]), .QN(n5964) );
  DFFRS_X2 \DATA_OUT_reg[3]  ( .D(n14195), .CK(N28803), .RN(n14193), .SN(
        n14194), .Q(DATA_OUT[3]), .QN(n5963) );
  DFFRS_X2 \DATA_OUT_reg[2]  ( .D(n14192), .CK(N28803), .RN(n14190), .SN(
        n14191), .Q(DATA_OUT[2]), .QN(n5962) );
  DFFRS_X2 \DATA_OUT_reg[1]  ( .D(n14189), .CK(N28803), .RN(n14187), .SN(
        n14188), .Q(DATA_OUT[1]), .QN(n5961) );
  DFFRS_X2 \DATA_OUT_reg[0]  ( .D(n14186), .CK(N28803), .RN(n14184), .SN(
        n14185), .Q(DATA_OUT[0]), .QN(n5960) );
  INV_X2 U10089 ( .A(CLK), .ZN(N28803) );
  AND2_X1 U3 ( .A1(n5953), .A2(ADDR[0]), .ZN(n5909) );
  AND2_X1 U4 ( .A1(n5959), .A2(ADDR[0]), .ZN(n5900) );
  AND2_X1 U5 ( .A1(n5953), .A2(ADDR[0]), .ZN(n1025) );
  AND2_X1 U6 ( .A1(n5959), .A2(n14982), .ZN(n5901) );
  AND2_X1 U7 ( .A1(n5959), .A2(ADDR[0]), .ZN(n763) );
  OR3_X1 U8 ( .A1(ADDR[0]), .A2(ADDR[3]), .A3(n14988), .ZN(n435) );
  OR3_X1 U9 ( .A1(ADDR[2]), .A2(ADDR[3]), .A3(ADDR[0]), .ZN(n5906) );
  OR3_X1 U10 ( .A1(ADDR[2]), .A2(ADDR[3]), .A3(ADDR[0]), .ZN(n171) );
  OR3_X1 U11 ( .A1(ADDR[0]), .A2(ADDR[3]), .A3(n14988), .ZN(n5905) );
  AND2_X1 U12 ( .A1(n5953), .A2(ADDR[0]), .ZN(n5908) );
  AND2_X1 U13 ( .A1(n5959), .A2(n14982), .ZN(n697) );
  AND2_X1 U14 ( .A1(n5959), .A2(ADDR[0]), .ZN(n5898) );
  NOR3_X1 U15 ( .A1(OFFSET[3]), .A2(OFFSET[4]), .A3(OFFSET[2]), .ZN(n1094) );
  NOR3_X1 U16 ( .A1(OFFSET[3]), .A2(OFFSET[4]), .A3(n5887), .ZN(n1107) );
  NOR3_X1 U17 ( .A1(OFFSET[2]), .A2(OFFSET[4]), .A3(n5888), .ZN(n1116) );
  NOR3_X1 U18 ( .A1(n5887), .A2(OFFSET[4]), .A3(n5888), .ZN(n1125) );
  NOR2_X1 U19 ( .A1(OFFSET[0]), .A2(OFFSET[1]), .ZN(n1095) );
  NOR2_X1 U20 ( .A1(n1164), .A2(OFFSET[1]), .ZN(n1098) );
  INV_X1 U21 ( .A(N147559), .ZN(n68) );
  INV_X1 U22 ( .A(DATA_IN[1]), .ZN(n69) );
  INV_X1 U23 ( .A(DATA_IN[2]), .ZN(n70) );
  INV_X1 U24 ( .A(DATA_IN[3]), .ZN(n71) );
  INV_X1 U25 ( .A(DATA_IN[4]), .ZN(n72) );
  INV_X1 U26 ( .A(DATA_IN[5]), .ZN(n73) );
  INV_X1 U27 ( .A(DATA_IN[6]), .ZN(n74) );
  INV_X1 U28 ( .A(DATA_IN[7]), .ZN(n75) );
  BUF_X1 U29 ( .A(n175), .Z(n14603) );
  BUF_X1 U30 ( .A(n175), .Z(n14604) );
  BUF_X1 U31 ( .A(n634), .Z(n14494) );
  BUF_X1 U32 ( .A(n634), .Z(n14495) );
  BUF_X1 U33 ( .A(n700), .Z(n14451) );
  BUF_X1 U34 ( .A(n700), .Z(n14452) );
  BUF_X1 U35 ( .A(n962), .Z(n14352) );
  BUF_X1 U36 ( .A(n962), .Z(n14353) );
  BUF_X1 U37 ( .A(n14646), .Z(n14648) );
  BUF_X1 U38 ( .A(n14646), .Z(n14647) );
  BUF_X1 U39 ( .A(n307), .Z(n14597) );
  BUF_X1 U40 ( .A(n307), .Z(n14598) );
  BUF_X1 U41 ( .A(n766), .Z(n14408) );
  BUF_X1 U42 ( .A(n766), .Z(n14409) );
  BUF_X1 U43 ( .A(n831), .Z(n14405) );
  BUF_X1 U44 ( .A(n831), .Z(n14406) );
  BUF_X1 U45 ( .A(n1093), .Z(n14306) );
  BUF_X1 U46 ( .A(n1093), .Z(n14307) );
  BUF_X1 U47 ( .A(n14593), .Z(n14595) );
  BUF_X1 U48 ( .A(n14593), .Z(n14594) );
  BUF_X1 U49 ( .A(n14552), .Z(n14550) );
  BUF_X1 U50 ( .A(n14552), .Z(n14549) );
  BUF_X1 U51 ( .A(n14404), .Z(n14402) );
  BUF_X1 U52 ( .A(n14404), .Z(n14401) );
  AND2_X1 U53 ( .A1(n1094), .A2(n1095), .ZN(n5727) );
  AND2_X1 U54 ( .A1(n1107), .A2(n1101), .ZN(n5729) );
  AND2_X1 U55 ( .A1(n1107), .A2(n1104), .ZN(n5730) );
  AND2_X1 U56 ( .A1(n1116), .A2(n1095), .ZN(n5738) );
  AND2_X1 U57 ( .A1(n1116), .A2(n1098), .ZN(n5739) );
  AND2_X1 U58 ( .A1(n1116), .A2(n1101), .ZN(n5741) );
  AND2_X1 U59 ( .A1(n1116), .A2(n1104), .ZN(n5742) );
  AND2_X1 U60 ( .A1(n1125), .A2(n1095), .ZN(n5746) );
  AND2_X1 U61 ( .A1(n1125), .A2(n1098), .ZN(n5747) );
  AND2_X1 U62 ( .A1(n1125), .A2(n1101), .ZN(n5749) );
  AND2_X1 U63 ( .A1(n1125), .A2(n1104), .ZN(n5750) );
  AND2_X1 U64 ( .A1(n1107), .A2(n1095), .ZN(n5754) );
  AND2_X1 U65 ( .A1(n1107), .A2(n1098), .ZN(n5755) );
  AND2_X1 U66 ( .A1(n1098), .A2(n1094), .ZN(n5757) );
  AND2_X1 U67 ( .A1(n1101), .A2(n1094), .ZN(n5758) );
  AND2_X1 U68 ( .A1(n1104), .A2(n1094), .ZN(n5762) );
  AND2_X1 U69 ( .A1(n1134), .A2(n1104), .ZN(n5763) );
  AND2_X1 U70 ( .A1(n1143), .A2(n1104), .ZN(n5765) );
  AND2_X1 U71 ( .A1(n1152), .A2(n1104), .ZN(n5766) );
  AND2_X1 U72 ( .A1(n1161), .A2(n1104), .ZN(n5774) );
  AND2_X1 U73 ( .A1(n1134), .A2(n1101), .ZN(n5775) );
  AND2_X1 U74 ( .A1(n1143), .A2(n1101), .ZN(n5777) );
  AND2_X1 U75 ( .A1(n1152), .A2(n1101), .ZN(n5778) );
  AND2_X1 U76 ( .A1(n1161), .A2(n1101), .ZN(n5782) );
  AND2_X1 U77 ( .A1(n1134), .A2(n1095), .ZN(n5783) );
  AND2_X1 U78 ( .A1(n1143), .A2(n1095), .ZN(n5785) );
  AND2_X1 U79 ( .A1(n1152), .A2(n1095), .ZN(n5786) );
  AND2_X1 U80 ( .A1(n1161), .A2(n1095), .ZN(n5790) );
  AND2_X1 U81 ( .A1(n1134), .A2(n1098), .ZN(n5791) );
  AND2_X1 U82 ( .A1(n1143), .A2(n1098), .ZN(n5793) );
  AND2_X1 U83 ( .A1(n1152), .A2(n1098), .ZN(n5794) );
  AND2_X1 U84 ( .A1(n1161), .A2(n1098), .ZN(n5798) );
  CLKBUF_X1 U85 ( .A(ADDR[1]), .Z(n14985) );
  CLKBUF_X1 U86 ( .A(ADDR[1]), .Z(n14984) );
  CLKBUF_X1 U87 ( .A(ADDR[1]), .Z(n14983) );
  CLKBUF_X1 U88 ( .A(ADDR[1]), .Z(n14986) );
  INV_X1 U89 ( .A(n241), .ZN(n240) );
  INV_X1 U90 ( .A(n244), .ZN(n243) );
  INV_X1 U91 ( .A(n246), .ZN(n245) );
  INV_X1 U92 ( .A(n248), .ZN(n247) );
  INV_X1 U93 ( .A(n250), .ZN(n249) );
  INV_X1 U94 ( .A(n252), .ZN(n251) );
  INV_X1 U95 ( .A(n503), .ZN(n502) );
  INV_X1 U96 ( .A(n506), .ZN(n505) );
  INV_X1 U97 ( .A(n508), .ZN(n507) );
  INV_X1 U98 ( .A(n510), .ZN(n509) );
  INV_X1 U99 ( .A(n512), .ZN(n511) );
  INV_X1 U100 ( .A(n514), .ZN(n513) );
  INV_X1 U101 ( .A(n568), .ZN(n567) );
  INV_X1 U102 ( .A(n571), .ZN(n570) );
  INV_X1 U103 ( .A(n573), .ZN(n572) );
  INV_X1 U104 ( .A(n575), .ZN(n574) );
  INV_X1 U105 ( .A(n577), .ZN(n576) );
  INV_X1 U106 ( .A(n579), .ZN(n578) );
  INV_X1 U107 ( .A(n1027), .ZN(n1026) );
  INV_X1 U108 ( .A(n1030), .ZN(n1029) );
  INV_X1 U109 ( .A(n1032), .ZN(n1031) );
  INV_X1 U110 ( .A(n1034), .ZN(n1033) );
  INV_X1 U111 ( .A(n1036), .ZN(n1035) );
  INV_X1 U112 ( .A(n1038), .ZN(n1037) );
  INV_X1 U113 ( .A(n227), .ZN(n226) );
  INV_X1 U114 ( .A(n229), .ZN(n228) );
  INV_X1 U115 ( .A(n231), .ZN(n230) );
  INV_X1 U116 ( .A(n233), .ZN(n232) );
  INV_X1 U117 ( .A(n235), .ZN(n234) );
  INV_X1 U118 ( .A(n237), .ZN(n236) );
  INV_X1 U119 ( .A(n359), .ZN(n358) );
  INV_X1 U120 ( .A(n361), .ZN(n360) );
  INV_X1 U121 ( .A(n363), .ZN(n362) );
  INV_X1 U122 ( .A(n365), .ZN(n364) );
  INV_X1 U123 ( .A(n367), .ZN(n366) );
  INV_X1 U124 ( .A(n369), .ZN(n368) );
  INV_X1 U125 ( .A(n686), .ZN(n685) );
  INV_X1 U126 ( .A(n688), .ZN(n687) );
  INV_X1 U127 ( .A(n690), .ZN(n689) );
  INV_X1 U128 ( .A(n692), .ZN(n691) );
  INV_X1 U129 ( .A(n694), .ZN(n693) );
  INV_X1 U130 ( .A(n696), .ZN(n695) );
  INV_X1 U131 ( .A(n752), .ZN(n751) );
  INV_X1 U132 ( .A(n754), .ZN(n753) );
  INV_X1 U133 ( .A(n756), .ZN(n755) );
  INV_X1 U134 ( .A(n758), .ZN(n757) );
  INV_X1 U135 ( .A(n760), .ZN(n759) );
  INV_X1 U136 ( .A(n762), .ZN(n761) );
  INV_X1 U137 ( .A(n818), .ZN(n817) );
  INV_X1 U138 ( .A(n820), .ZN(n819) );
  INV_X1 U139 ( .A(n822), .ZN(n821) );
  INV_X1 U140 ( .A(n824), .ZN(n823) );
  INV_X1 U141 ( .A(n826), .ZN(n825) );
  INV_X1 U142 ( .A(n828), .ZN(n827) );
  INV_X1 U143 ( .A(n883), .ZN(n882) );
  INV_X1 U144 ( .A(n885), .ZN(n884) );
  INV_X1 U145 ( .A(n887), .ZN(n886) );
  INV_X1 U146 ( .A(n889), .ZN(n888) );
  INV_X1 U147 ( .A(n891), .ZN(n890) );
  INV_X1 U148 ( .A(n893), .ZN(n892) );
  INV_X1 U149 ( .A(n1014), .ZN(n1013) );
  INV_X1 U150 ( .A(n1016), .ZN(n1015) );
  INV_X1 U151 ( .A(n1018), .ZN(n1017) );
  INV_X1 U152 ( .A(n1020), .ZN(n1019) );
  INV_X1 U153 ( .A(n1022), .ZN(n1021) );
  INV_X1 U154 ( .A(n1024), .ZN(n1023) );
  INV_X1 U155 ( .A(n1156), .ZN(n1155) );
  INV_X1 U156 ( .A(n1158), .ZN(n1157) );
  INV_X1 U157 ( .A(n1160), .ZN(n1159) );
  INV_X1 U158 ( .A(n1163), .ZN(n1162) );
  INV_X1 U159 ( .A(n1166), .ZN(n1165) );
  INV_X1 U160 ( .A(n1168), .ZN(n1167) );
  INV_X1 U161 ( .A(n437), .ZN(n436) );
  INV_X1 U162 ( .A(n440), .ZN(n439) );
  INV_X1 U163 ( .A(n442), .ZN(n441) );
  INV_X1 U164 ( .A(n444), .ZN(n443) );
  INV_X1 U165 ( .A(n446), .ZN(n445) );
  INV_X1 U166 ( .A(n448), .ZN(n447) );
  INV_X1 U167 ( .A(n895), .ZN(n894) );
  INV_X1 U168 ( .A(n898), .ZN(n897) );
  INV_X1 U169 ( .A(n900), .ZN(n899) );
  INV_X1 U170 ( .A(n902), .ZN(n901) );
  INV_X1 U171 ( .A(n904), .ZN(n903) );
  INV_X1 U172 ( .A(n906), .ZN(n905) );
  INV_X1 U173 ( .A(n254), .ZN(n253) );
  INV_X1 U174 ( .A(n256), .ZN(n255) );
  INV_X1 U175 ( .A(n258), .ZN(n257) );
  INV_X1 U176 ( .A(n260), .ZN(n259) );
  INV_X1 U177 ( .A(n262), .ZN(n261) );
  INV_X1 U178 ( .A(n264), .ZN(n263) );
  INV_X1 U179 ( .A(n266), .ZN(n265) );
  INV_X1 U180 ( .A(n268), .ZN(n267) );
  INV_X1 U181 ( .A(n270), .ZN(n269) );
  INV_X1 U182 ( .A(n272), .ZN(n271) );
  INV_X1 U183 ( .A(n274), .ZN(n273) );
  INV_X1 U184 ( .A(n276), .ZN(n275) );
  INV_X1 U185 ( .A(n278), .ZN(n277) );
  INV_X1 U186 ( .A(n280), .ZN(n279) );
  INV_X1 U187 ( .A(n282), .ZN(n281) );
  INV_X1 U188 ( .A(n284), .ZN(n283) );
  INV_X1 U189 ( .A(n286), .ZN(n285) );
  INV_X1 U190 ( .A(n288), .ZN(n287) );
  INV_X1 U191 ( .A(n290), .ZN(n289) );
  INV_X1 U192 ( .A(n292), .ZN(n291) );
  INV_X1 U193 ( .A(n294), .ZN(n293) );
  INV_X1 U194 ( .A(n296), .ZN(n295) );
  INV_X1 U195 ( .A(n298), .ZN(n297) );
  INV_X1 U196 ( .A(n300), .ZN(n299) );
  INV_X1 U197 ( .A(n302), .ZN(n301) );
  INV_X1 U198 ( .A(n304), .ZN(n303) );
  INV_X1 U199 ( .A(n516), .ZN(n515) );
  INV_X1 U200 ( .A(n518), .ZN(n517) );
  INV_X1 U201 ( .A(n520), .ZN(n519) );
  INV_X1 U202 ( .A(n522), .ZN(n521) );
  INV_X1 U203 ( .A(n524), .ZN(n523) );
  INV_X1 U204 ( .A(n526), .ZN(n525) );
  INV_X1 U205 ( .A(n528), .ZN(n527) );
  INV_X1 U206 ( .A(n530), .ZN(n529) );
  INV_X1 U207 ( .A(n532), .ZN(n531) );
  INV_X1 U208 ( .A(n534), .ZN(n533) );
  INV_X1 U209 ( .A(n536), .ZN(n535) );
  INV_X1 U210 ( .A(n538), .ZN(n537) );
  INV_X1 U211 ( .A(n540), .ZN(n539) );
  INV_X1 U212 ( .A(n542), .ZN(n541) );
  INV_X1 U213 ( .A(n544), .ZN(n543) );
  INV_X1 U214 ( .A(n546), .ZN(n545) );
  INV_X1 U215 ( .A(n548), .ZN(n547) );
  INV_X1 U216 ( .A(n550), .ZN(n549) );
  INV_X1 U217 ( .A(n552), .ZN(n551) );
  INV_X1 U218 ( .A(n554), .ZN(n553) );
  INV_X1 U219 ( .A(n556), .ZN(n555) );
  INV_X1 U220 ( .A(n558), .ZN(n557) );
  INV_X1 U221 ( .A(n560), .ZN(n559) );
  INV_X1 U222 ( .A(n562), .ZN(n561) );
  INV_X1 U223 ( .A(n564), .ZN(n563) );
  INV_X1 U224 ( .A(n566), .ZN(n565) );
  INV_X1 U225 ( .A(n581), .ZN(n580) );
  INV_X1 U226 ( .A(n583), .ZN(n582) );
  INV_X1 U227 ( .A(n585), .ZN(n584) );
  INV_X1 U228 ( .A(n587), .ZN(n586) );
  INV_X1 U229 ( .A(n589), .ZN(n588) );
  INV_X1 U230 ( .A(n591), .ZN(n590) );
  INV_X1 U231 ( .A(n593), .ZN(n592) );
  INV_X1 U232 ( .A(n595), .ZN(n594) );
  INV_X1 U233 ( .A(n597), .ZN(n596) );
  INV_X1 U234 ( .A(n599), .ZN(n598) );
  INV_X1 U235 ( .A(n601), .ZN(n600) );
  INV_X1 U236 ( .A(n603), .ZN(n602) );
  INV_X1 U237 ( .A(n605), .ZN(n604) );
  INV_X1 U238 ( .A(n607), .ZN(n606) );
  INV_X1 U239 ( .A(n609), .ZN(n608) );
  INV_X1 U240 ( .A(n611), .ZN(n610) );
  INV_X1 U241 ( .A(n613), .ZN(n612) );
  INV_X1 U242 ( .A(n615), .ZN(n614) );
  INV_X1 U243 ( .A(n617), .ZN(n616) );
  INV_X1 U244 ( .A(n619), .ZN(n618) );
  INV_X1 U245 ( .A(n621), .ZN(n620) );
  INV_X1 U246 ( .A(n623), .ZN(n622) );
  INV_X1 U247 ( .A(n625), .ZN(n624) );
  INV_X1 U248 ( .A(n627), .ZN(n626) );
  INV_X1 U249 ( .A(n629), .ZN(n628) );
  INV_X1 U250 ( .A(n631), .ZN(n630) );
  INV_X1 U251 ( .A(n1040), .ZN(n1039) );
  INV_X1 U252 ( .A(n1042), .ZN(n1041) );
  INV_X1 U253 ( .A(n1044), .ZN(n1043) );
  INV_X1 U254 ( .A(n1046), .ZN(n1045) );
  INV_X1 U255 ( .A(n1048), .ZN(n1047) );
  INV_X1 U256 ( .A(n1050), .ZN(n1049) );
  INV_X1 U257 ( .A(n1052), .ZN(n1051) );
  INV_X1 U258 ( .A(n1054), .ZN(n1053) );
  INV_X1 U259 ( .A(n1056), .ZN(n1055) );
  INV_X1 U260 ( .A(n1058), .ZN(n1057) );
  INV_X1 U261 ( .A(n1060), .ZN(n1059) );
  INV_X1 U262 ( .A(n1062), .ZN(n1061) );
  INV_X1 U263 ( .A(n1064), .ZN(n1063) );
  INV_X1 U264 ( .A(n1066), .ZN(n1065) );
  INV_X1 U265 ( .A(n1068), .ZN(n1067) );
  INV_X1 U266 ( .A(n1070), .ZN(n1069) );
  INV_X1 U267 ( .A(n1072), .ZN(n1071) );
  INV_X1 U268 ( .A(n1074), .ZN(n1073) );
  INV_X1 U269 ( .A(n1076), .ZN(n1075) );
  INV_X1 U270 ( .A(n1078), .ZN(n1077) );
  INV_X1 U271 ( .A(n1080), .ZN(n1079) );
  INV_X1 U272 ( .A(n1082), .ZN(n1081) );
  INV_X1 U273 ( .A(n1084), .ZN(n1083) );
  INV_X1 U274 ( .A(n1086), .ZN(n1085) );
  INV_X1 U275 ( .A(n1088), .ZN(n1087) );
  INV_X1 U276 ( .A(n1090), .ZN(n1089) );
  INV_X1 U277 ( .A(n410), .ZN(n409) );
  INV_X1 U278 ( .A(n412), .ZN(n411) );
  INV_X1 U279 ( .A(n414), .ZN(n413) );
  INV_X1 U280 ( .A(n416), .ZN(n415) );
  INV_X1 U281 ( .A(n418), .ZN(n417) );
  INV_X1 U282 ( .A(n420), .ZN(n419) );
  INV_X1 U283 ( .A(n422), .ZN(n421) );
  INV_X1 U284 ( .A(n424), .ZN(n423) );
  INV_X1 U285 ( .A(n426), .ZN(n425) );
  INV_X1 U286 ( .A(n428), .ZN(n427) );
  INV_X1 U287 ( .A(n430), .ZN(n429) );
  INV_X1 U288 ( .A(n432), .ZN(n431) );
  INV_X1 U289 ( .A(n434), .ZN(n433) );
  INV_X1 U290 ( .A(n476), .ZN(n475) );
  INV_X1 U291 ( .A(n478), .ZN(n477) );
  INV_X1 U292 ( .A(n480), .ZN(n479) );
  INV_X1 U293 ( .A(n482), .ZN(n481) );
  INV_X1 U294 ( .A(n484), .ZN(n483) );
  INV_X1 U295 ( .A(n486), .ZN(n485) );
  INV_X1 U296 ( .A(n488), .ZN(n487) );
  INV_X1 U297 ( .A(n490), .ZN(n489) );
  INV_X1 U298 ( .A(n492), .ZN(n491) );
  INV_X1 U299 ( .A(n494), .ZN(n493) );
  INV_X1 U300 ( .A(n496), .ZN(n495) );
  INV_X1 U301 ( .A(n498), .ZN(n497) );
  INV_X1 U302 ( .A(n500), .ZN(n499) );
  INV_X1 U303 ( .A(n934), .ZN(n933) );
  INV_X1 U304 ( .A(n936), .ZN(n935) );
  INV_X1 U305 ( .A(n938), .ZN(n937) );
  INV_X1 U306 ( .A(n940), .ZN(n939) );
  INV_X1 U307 ( .A(n942), .ZN(n941) );
  INV_X1 U308 ( .A(n944), .ZN(n943) );
  INV_X1 U309 ( .A(n946), .ZN(n945) );
  INV_X1 U310 ( .A(n948), .ZN(n947) );
  INV_X1 U311 ( .A(n950), .ZN(n949) );
  INV_X1 U312 ( .A(n952), .ZN(n951) );
  INV_X1 U313 ( .A(n954), .ZN(n953) );
  INV_X1 U314 ( .A(n956), .ZN(n955) );
  INV_X1 U315 ( .A(n958), .ZN(n957) );
  INV_X1 U316 ( .A(n370), .ZN(n371) );
  INV_X1 U317 ( .A(n373), .ZN(n374) );
  INV_X1 U318 ( .A(n375), .ZN(n376) );
  INV_X1 U319 ( .A(n377), .ZN(n378) );
  INV_X1 U320 ( .A(n379), .ZN(n380) );
  INV_X1 U321 ( .A(n381), .ZN(n382) );
  INV_X1 U322 ( .A(n79), .ZN(n78) );
  INV_X1 U323 ( .A(n82), .ZN(n81) );
  INV_X1 U324 ( .A(n85), .ZN(n84) );
  INV_X1 U325 ( .A(n88), .ZN(n87) );
  INV_X1 U326 ( .A(n91), .ZN(n90) );
  INV_X1 U327 ( .A(n67), .ZN(n66) );
  INV_X1 U328 ( .A(n133), .ZN(n132) );
  INV_X1 U329 ( .A(n136), .ZN(n135) );
  INV_X1 U330 ( .A(n139), .ZN(n138) );
  INV_X1 U331 ( .A(n142), .ZN(n141) );
  INV_X1 U332 ( .A(n145), .ZN(n144) );
  INV_X1 U333 ( .A(n148), .ZN(n147) );
  INV_X1 U334 ( .A(n151), .ZN(n150) );
  INV_X1 U335 ( .A(n154), .ZN(n153) );
  INV_X1 U336 ( .A(n157), .ZN(n156) );
  INV_X1 U337 ( .A(n160), .ZN(n159) );
  INV_X1 U338 ( .A(n163), .ZN(n162) );
  INV_X1 U339 ( .A(n166), .ZN(n165) );
  INV_X1 U340 ( .A(n169), .ZN(n168) );
  INV_X1 U341 ( .A(n94), .ZN(n93) );
  INV_X1 U342 ( .A(n97), .ZN(n96) );
  INV_X1 U343 ( .A(n100), .ZN(n99) );
  INV_X1 U344 ( .A(n103), .ZN(n102) );
  INV_X1 U345 ( .A(n106), .ZN(n105) );
  INV_X1 U346 ( .A(n109), .ZN(n108) );
  INV_X1 U347 ( .A(n112), .ZN(n111) );
  INV_X1 U348 ( .A(n115), .ZN(n114) );
  INV_X1 U349 ( .A(n118), .ZN(n117) );
  INV_X1 U350 ( .A(n121), .ZN(n120) );
  INV_X1 U351 ( .A(n124), .ZN(n123) );
  INV_X1 U352 ( .A(n127), .ZN(n126) );
  INV_X1 U353 ( .A(n130), .ZN(n129) );
  INV_X1 U354 ( .A(n174), .ZN(n173) );
  INV_X1 U355 ( .A(n177), .ZN(n176) );
  INV_X1 U356 ( .A(n179), .ZN(n178) );
  INV_X1 U357 ( .A(n181), .ZN(n180) );
  INV_X1 U358 ( .A(n183), .ZN(n182) );
  INV_X1 U359 ( .A(n185), .ZN(n184) );
  INV_X1 U360 ( .A(n187), .ZN(n186) );
  INV_X1 U361 ( .A(n189), .ZN(n188) );
  INV_X1 U362 ( .A(n191), .ZN(n190) );
  INV_X1 U363 ( .A(n193), .ZN(n192) );
  INV_X1 U364 ( .A(n195), .ZN(n194) );
  INV_X1 U365 ( .A(n197), .ZN(n196) );
  INV_X1 U366 ( .A(n199), .ZN(n198) );
  INV_X1 U367 ( .A(n201), .ZN(n200) );
  INV_X1 U368 ( .A(n203), .ZN(n202) );
  INV_X1 U369 ( .A(n205), .ZN(n204) );
  INV_X1 U370 ( .A(n207), .ZN(n206) );
  INV_X1 U371 ( .A(n209), .ZN(n208) );
  INV_X1 U372 ( .A(n211), .ZN(n210) );
  INV_X1 U373 ( .A(n213), .ZN(n212) );
  INV_X1 U374 ( .A(n215), .ZN(n214) );
  INV_X1 U375 ( .A(n217), .ZN(n216) );
  INV_X1 U376 ( .A(n219), .ZN(n218) );
  INV_X1 U377 ( .A(n221), .ZN(n220) );
  INV_X1 U378 ( .A(n223), .ZN(n222) );
  INV_X1 U379 ( .A(n225), .ZN(n224) );
  INV_X1 U380 ( .A(n306), .ZN(n305) );
  INV_X1 U381 ( .A(n309), .ZN(n308) );
  INV_X1 U382 ( .A(n311), .ZN(n310) );
  INV_X1 U383 ( .A(n313), .ZN(n312) );
  INV_X1 U384 ( .A(n315), .ZN(n314) );
  INV_X1 U385 ( .A(n317), .ZN(n316) );
  INV_X1 U386 ( .A(n319), .ZN(n318) );
  INV_X1 U387 ( .A(n321), .ZN(n320) );
  INV_X1 U388 ( .A(n323), .ZN(n322) );
  INV_X1 U389 ( .A(n325), .ZN(n324) );
  INV_X1 U390 ( .A(n327), .ZN(n326) );
  INV_X1 U391 ( .A(n329), .ZN(n328) );
  INV_X1 U392 ( .A(n331), .ZN(n330) );
  INV_X1 U393 ( .A(n333), .ZN(n332) );
  INV_X1 U394 ( .A(n335), .ZN(n334) );
  INV_X1 U395 ( .A(n337), .ZN(n336) );
  INV_X1 U396 ( .A(n339), .ZN(n338) );
  INV_X1 U397 ( .A(n341), .ZN(n340) );
  INV_X1 U398 ( .A(n343), .ZN(n342) );
  INV_X1 U399 ( .A(n345), .ZN(n344) );
  INV_X1 U400 ( .A(n347), .ZN(n346) );
  INV_X1 U401 ( .A(n349), .ZN(n348) );
  INV_X1 U402 ( .A(n351), .ZN(n350) );
  INV_X1 U403 ( .A(n353), .ZN(n352) );
  INV_X1 U404 ( .A(n355), .ZN(n354) );
  INV_X1 U405 ( .A(n357), .ZN(n356) );
  INV_X1 U406 ( .A(n398), .ZN(n397) );
  INV_X1 U407 ( .A(n400), .ZN(n399) );
  INV_X1 U408 ( .A(n402), .ZN(n401) );
  INV_X1 U409 ( .A(n404), .ZN(n403) );
  INV_X1 U410 ( .A(n406), .ZN(n405) );
  INV_X1 U411 ( .A(n408), .ZN(n407) );
  INV_X1 U412 ( .A(n450), .ZN(n449) );
  INV_X1 U413 ( .A(n452), .ZN(n451) );
  INV_X1 U414 ( .A(n454), .ZN(n453) );
  INV_X1 U415 ( .A(n456), .ZN(n455) );
  INV_X1 U416 ( .A(n458), .ZN(n457) );
  INV_X1 U417 ( .A(n460), .ZN(n459) );
  INV_X1 U418 ( .A(n462), .ZN(n461) );
  INV_X1 U419 ( .A(n464), .ZN(n463) );
  INV_X1 U420 ( .A(n466), .ZN(n465) );
  INV_X1 U421 ( .A(n468), .ZN(n467) );
  INV_X1 U422 ( .A(n470), .ZN(n469) );
  INV_X1 U423 ( .A(n472), .ZN(n471) );
  INV_X1 U424 ( .A(n474), .ZN(n473) );
  INV_X1 U425 ( .A(n633), .ZN(n632) );
  INV_X1 U426 ( .A(n636), .ZN(n635) );
  INV_X1 U427 ( .A(n638), .ZN(n637) );
  INV_X1 U428 ( .A(n640), .ZN(n639) );
  INV_X1 U429 ( .A(n642), .ZN(n641) );
  INV_X1 U430 ( .A(n644), .ZN(n643) );
  INV_X1 U431 ( .A(n646), .ZN(n645) );
  INV_X1 U432 ( .A(n648), .ZN(n647) );
  INV_X1 U433 ( .A(n650), .ZN(n649) );
  INV_X1 U434 ( .A(n652), .ZN(n651) );
  INV_X1 U435 ( .A(n654), .ZN(n653) );
  INV_X1 U436 ( .A(n656), .ZN(n655) );
  INV_X1 U437 ( .A(n658), .ZN(n657) );
  INV_X1 U438 ( .A(n660), .ZN(n659) );
  INV_X1 U439 ( .A(n662), .ZN(n661) );
  INV_X1 U440 ( .A(n664), .ZN(n663) );
  INV_X1 U441 ( .A(n666), .ZN(n665) );
  INV_X1 U442 ( .A(n668), .ZN(n667) );
  INV_X1 U443 ( .A(n670), .ZN(n669) );
  INV_X1 U444 ( .A(n672), .ZN(n671) );
  INV_X1 U445 ( .A(n674), .ZN(n673) );
  INV_X1 U446 ( .A(n676), .ZN(n675) );
  INV_X1 U447 ( .A(n678), .ZN(n677) );
  INV_X1 U448 ( .A(n680), .ZN(n679) );
  INV_X1 U449 ( .A(n682), .ZN(n681) );
  INV_X1 U450 ( .A(n684), .ZN(n683) );
  INV_X1 U451 ( .A(n699), .ZN(n698) );
  INV_X1 U452 ( .A(n702), .ZN(n701) );
  INV_X1 U453 ( .A(n704), .ZN(n703) );
  INV_X1 U454 ( .A(n706), .ZN(n705) );
  INV_X1 U455 ( .A(n708), .ZN(n707) );
  INV_X1 U456 ( .A(n710), .ZN(n709) );
  INV_X1 U457 ( .A(n712), .ZN(n711) );
  INV_X1 U458 ( .A(n714), .ZN(n713) );
  INV_X1 U459 ( .A(n716), .ZN(n715) );
  INV_X1 U460 ( .A(n718), .ZN(n717) );
  INV_X1 U461 ( .A(n720), .ZN(n719) );
  INV_X1 U462 ( .A(n722), .ZN(n721) );
  INV_X1 U463 ( .A(n724), .ZN(n723) );
  INV_X1 U464 ( .A(n726), .ZN(n725) );
  INV_X1 U465 ( .A(n728), .ZN(n727) );
  INV_X1 U466 ( .A(n730), .ZN(n729) );
  INV_X1 U467 ( .A(n732), .ZN(n731) );
  INV_X1 U468 ( .A(n734), .ZN(n733) );
  INV_X1 U469 ( .A(n736), .ZN(n735) );
  INV_X1 U470 ( .A(n738), .ZN(n737) );
  INV_X1 U471 ( .A(n740), .ZN(n739) );
  INV_X1 U472 ( .A(n742), .ZN(n741) );
  INV_X1 U473 ( .A(n744), .ZN(n743) );
  INV_X1 U474 ( .A(n746), .ZN(n745) );
  INV_X1 U475 ( .A(n748), .ZN(n747) );
  INV_X1 U476 ( .A(n750), .ZN(n749) );
  INV_X1 U477 ( .A(n765), .ZN(n764) );
  INV_X1 U478 ( .A(n768), .ZN(n767) );
  INV_X1 U479 ( .A(n770), .ZN(n769) );
  INV_X1 U480 ( .A(n772), .ZN(n771) );
  INV_X1 U481 ( .A(n774), .ZN(n773) );
  INV_X1 U482 ( .A(n776), .ZN(n775) );
  INV_X1 U483 ( .A(n778), .ZN(n777) );
  INV_X1 U484 ( .A(n780), .ZN(n779) );
  INV_X1 U485 ( .A(n782), .ZN(n781) );
  INV_X1 U486 ( .A(n784), .ZN(n783) );
  INV_X1 U487 ( .A(n786), .ZN(n785) );
  INV_X1 U488 ( .A(n788), .ZN(n787) );
  INV_X1 U489 ( .A(n790), .ZN(n789) );
  INV_X1 U490 ( .A(n792), .ZN(n791) );
  INV_X1 U491 ( .A(n794), .ZN(n793) );
  INV_X1 U492 ( .A(n796), .ZN(n795) );
  INV_X1 U493 ( .A(n798), .ZN(n797) );
  INV_X1 U494 ( .A(n800), .ZN(n799) );
  INV_X1 U495 ( .A(n802), .ZN(n801) );
  INV_X1 U496 ( .A(n804), .ZN(n803) );
  INV_X1 U497 ( .A(n806), .ZN(n805) );
  INV_X1 U498 ( .A(n808), .ZN(n807) );
  INV_X1 U499 ( .A(n810), .ZN(n809) );
  INV_X1 U500 ( .A(n812), .ZN(n811) );
  INV_X1 U501 ( .A(n814), .ZN(n813) );
  INV_X1 U502 ( .A(n816), .ZN(n815) );
  INV_X1 U503 ( .A(n830), .ZN(n829) );
  INV_X1 U504 ( .A(n833), .ZN(n832) );
  INV_X1 U505 ( .A(n835), .ZN(n834) );
  INV_X1 U506 ( .A(n837), .ZN(n836) );
  INV_X1 U507 ( .A(n839), .ZN(n838) );
  INV_X1 U508 ( .A(n841), .ZN(n840) );
  INV_X1 U509 ( .A(n843), .ZN(n842) );
  INV_X1 U510 ( .A(n845), .ZN(n844) );
  INV_X1 U511 ( .A(n847), .ZN(n846) );
  INV_X1 U512 ( .A(n849), .ZN(n848) );
  INV_X1 U513 ( .A(n851), .ZN(n850) );
  INV_X1 U514 ( .A(n853), .ZN(n852) );
  INV_X1 U515 ( .A(n855), .ZN(n854) );
  INV_X1 U516 ( .A(n857), .ZN(n856) );
  INV_X1 U517 ( .A(n859), .ZN(n858) );
  INV_X1 U518 ( .A(n861), .ZN(n860) );
  INV_X1 U519 ( .A(n863), .ZN(n862) );
  INV_X1 U520 ( .A(n865), .ZN(n864) );
  INV_X1 U521 ( .A(n867), .ZN(n866) );
  INV_X1 U522 ( .A(n869), .ZN(n868) );
  INV_X1 U523 ( .A(n871), .ZN(n870) );
  INV_X1 U524 ( .A(n873), .ZN(n872) );
  INV_X1 U525 ( .A(n875), .ZN(n874) );
  INV_X1 U526 ( .A(n877), .ZN(n876) );
  INV_X1 U527 ( .A(n879), .ZN(n878) );
  INV_X1 U528 ( .A(n881), .ZN(n880) );
  INV_X1 U529 ( .A(n908), .ZN(n907) );
  INV_X1 U530 ( .A(n910), .ZN(n909) );
  INV_X1 U531 ( .A(n912), .ZN(n911) );
  INV_X1 U532 ( .A(n914), .ZN(n913) );
  INV_X1 U533 ( .A(n916), .ZN(n915) );
  INV_X1 U534 ( .A(n918), .ZN(n917) );
  INV_X1 U535 ( .A(n920), .ZN(n919) );
  INV_X1 U536 ( .A(n922), .ZN(n921) );
  INV_X1 U537 ( .A(n924), .ZN(n923) );
  INV_X1 U538 ( .A(n926), .ZN(n925) );
  INV_X1 U539 ( .A(n928), .ZN(n927) );
  INV_X1 U540 ( .A(n930), .ZN(n929) );
  INV_X1 U541 ( .A(n932), .ZN(n931) );
  INV_X1 U542 ( .A(n961), .ZN(n960) );
  INV_X1 U543 ( .A(n964), .ZN(n963) );
  INV_X1 U544 ( .A(n966), .ZN(n965) );
  INV_X1 U545 ( .A(n968), .ZN(n967) );
  INV_X1 U546 ( .A(n970), .ZN(n969) );
  INV_X1 U547 ( .A(n972), .ZN(n971) );
  INV_X1 U548 ( .A(n974), .ZN(n973) );
  INV_X1 U549 ( .A(n976), .ZN(n975) );
  INV_X1 U550 ( .A(n978), .ZN(n977) );
  INV_X1 U551 ( .A(n980), .ZN(n979) );
  INV_X1 U552 ( .A(n982), .ZN(n981) );
  INV_X1 U553 ( .A(n984), .ZN(n983) );
  INV_X1 U554 ( .A(n986), .ZN(n985) );
  INV_X1 U555 ( .A(n988), .ZN(n987) );
  INV_X1 U556 ( .A(n990), .ZN(n989) );
  INV_X1 U557 ( .A(n992), .ZN(n991) );
  INV_X1 U558 ( .A(n994), .ZN(n993) );
  INV_X1 U559 ( .A(n996), .ZN(n995) );
  INV_X1 U560 ( .A(n998), .ZN(n997) );
  INV_X1 U561 ( .A(n1000), .ZN(n999) );
  INV_X1 U562 ( .A(n1002), .ZN(n1001) );
  INV_X1 U563 ( .A(n1004), .ZN(n1003) );
  INV_X1 U564 ( .A(n1006), .ZN(n1005) );
  INV_X1 U565 ( .A(n1008), .ZN(n1007) );
  INV_X1 U566 ( .A(n1010), .ZN(n1009) );
  INV_X1 U567 ( .A(n1012), .ZN(n1011) );
  INV_X1 U568 ( .A(n1092), .ZN(n1091) );
  INV_X1 U569 ( .A(n1097), .ZN(n1096) );
  INV_X1 U570 ( .A(n1100), .ZN(n1099) );
  INV_X1 U571 ( .A(n1103), .ZN(n1102) );
  INV_X1 U572 ( .A(n1106), .ZN(n1105) );
  INV_X1 U573 ( .A(n1109), .ZN(n1108) );
  INV_X1 U574 ( .A(n1111), .ZN(n1110) );
  INV_X1 U575 ( .A(n1113), .ZN(n1112) );
  INV_X1 U576 ( .A(n1115), .ZN(n1114) );
  INV_X1 U577 ( .A(n1118), .ZN(n1117) );
  INV_X1 U578 ( .A(n1120), .ZN(n1119) );
  INV_X1 U579 ( .A(n1122), .ZN(n1121) );
  INV_X1 U580 ( .A(n1124), .ZN(n1123) );
  INV_X1 U581 ( .A(n1127), .ZN(n1126) );
  INV_X1 U582 ( .A(n1129), .ZN(n1128) );
  INV_X1 U583 ( .A(n1131), .ZN(n1130) );
  INV_X1 U584 ( .A(n1133), .ZN(n1132) );
  INV_X1 U585 ( .A(n1136), .ZN(n1135) );
  INV_X1 U586 ( .A(n1138), .ZN(n1137) );
  INV_X1 U587 ( .A(n1140), .ZN(n1139) );
  INV_X1 U588 ( .A(n1142), .ZN(n1141) );
  INV_X1 U589 ( .A(n1145), .ZN(n1144) );
  INV_X1 U590 ( .A(n1147), .ZN(n1146) );
  INV_X1 U591 ( .A(n1149), .ZN(n1148) );
  INV_X1 U592 ( .A(n1151), .ZN(n1150) );
  INV_X1 U593 ( .A(n1154), .ZN(n1153) );
  INV_X1 U594 ( .A(n383), .ZN(n384) );
  INV_X1 U595 ( .A(n385), .ZN(n386) );
  INV_X1 U596 ( .A(n387), .ZN(n388) );
  INV_X1 U597 ( .A(n389), .ZN(n390) );
  INV_X1 U598 ( .A(n391), .ZN(n392) );
  INV_X1 U599 ( .A(n393), .ZN(n394) );
  INV_X1 U600 ( .A(n395), .ZN(n396) );
  INV_X1 U601 ( .A(n14976), .ZN(n14970) );
  INV_X1 U602 ( .A(n14976), .ZN(n14971) );
  INV_X1 U603 ( .A(n14975), .ZN(n14972) );
  BUF_X1 U604 ( .A(n14974), .Z(n14976) );
  BUF_X1 U605 ( .A(n242), .Z(n14602) );
  BUF_X1 U606 ( .A(n504), .Z(n14502) );
  BUF_X1 U607 ( .A(n569), .Z(n14499) );
  BUF_X1 U608 ( .A(n1028), .Z(n14311) );
  BUF_X1 U609 ( .A(n175), .Z(n14605) );
  BUF_X1 U610 ( .A(n634), .Z(n14496) );
  BUF_X1 U611 ( .A(n700), .Z(n14453) );
  BUF_X1 U612 ( .A(n962), .Z(n14354) );
  BUF_X1 U613 ( .A(n242), .Z(n14601) );
  BUF_X1 U614 ( .A(n242), .Z(n14600) );
  BUF_X1 U615 ( .A(n504), .Z(n14501) );
  BUF_X1 U616 ( .A(n504), .Z(n14500) );
  BUF_X1 U617 ( .A(n569), .Z(n14498) );
  BUF_X1 U618 ( .A(n569), .Z(n14497) );
  BUF_X1 U619 ( .A(n1028), .Z(n14310) );
  BUF_X1 U620 ( .A(n1028), .Z(n14309) );
  NAND2_X1 U621 ( .A1(n5757), .A2(n14649), .ZN(n79) );
  NAND2_X1 U622 ( .A1(n5758), .A2(n14649), .ZN(n82) );
  NAND2_X1 U623 ( .A1(n5762), .A2(n14649), .ZN(n85) );
  NAND2_X1 U624 ( .A1(n5754), .A2(n14649), .ZN(n88) );
  NAND2_X1 U625 ( .A1(n5755), .A2(n14649), .ZN(n91) );
  NAND2_X1 U626 ( .A1(n5727), .A2(n14649), .ZN(n67) );
  NAND2_X1 U627 ( .A1(n14596), .A2(n5727), .ZN(n370) );
  NAND2_X1 U628 ( .A1(n14596), .A2(n5757), .ZN(n373) );
  NAND2_X1 U629 ( .A1(n14596), .A2(n5758), .ZN(n375) );
  NAND2_X1 U630 ( .A1(n14596), .A2(n5762), .ZN(n377) );
  NAND2_X1 U631 ( .A1(n14596), .A2(n5754), .ZN(n379) );
  NAND2_X1 U632 ( .A1(n14596), .A2(n5755), .ZN(n381) );
  NAND2_X1 U633 ( .A1(n14551), .A2(n5727), .ZN(n437) );
  NAND2_X1 U634 ( .A1(n14551), .A2(n5757), .ZN(n440) );
  NAND2_X1 U635 ( .A1(n14551), .A2(n5758), .ZN(n442) );
  NAND2_X1 U636 ( .A1(n14551), .A2(n5762), .ZN(n444) );
  NAND2_X1 U637 ( .A1(n14551), .A2(n5754), .ZN(n446) );
  NAND2_X1 U638 ( .A1(n14551), .A2(n5755), .ZN(n448) );
  NAND2_X1 U639 ( .A1(n14403), .A2(n5727), .ZN(n895) );
  NAND2_X1 U640 ( .A1(n14403), .A2(n5757), .ZN(n898) );
  NAND2_X1 U641 ( .A1(n14403), .A2(n5758), .ZN(n900) );
  NAND2_X1 U642 ( .A1(n14403), .A2(n5762), .ZN(n902) );
  NAND2_X1 U643 ( .A1(n14403), .A2(n5754), .ZN(n904) );
  NAND2_X1 U644 ( .A1(n14403), .A2(n5755), .ZN(n906) );
  NAND2_X1 U645 ( .A1(n14605), .A2(n5778), .ZN(n227) );
  NAND2_X1 U646 ( .A1(n14605), .A2(n5766), .ZN(n229) );
  NAND2_X1 U647 ( .A1(n14605), .A2(n5790), .ZN(n231) );
  NAND2_X1 U648 ( .A1(n14605), .A2(n5798), .ZN(n233) );
  NAND2_X1 U649 ( .A1(n14605), .A2(n5782), .ZN(n235) );
  NAND2_X1 U650 ( .A1(n14605), .A2(n5774), .ZN(n237) );
  NAND2_X1 U651 ( .A1(n14599), .A2(n5778), .ZN(n359) );
  NAND2_X1 U652 ( .A1(n14599), .A2(n5766), .ZN(n361) );
  NAND2_X1 U653 ( .A1(n14599), .A2(n5790), .ZN(n363) );
  NAND2_X1 U654 ( .A1(n14599), .A2(n5798), .ZN(n365) );
  NAND2_X1 U655 ( .A1(n14599), .A2(n5782), .ZN(n367) );
  NAND2_X1 U656 ( .A1(n14599), .A2(n5774), .ZN(n369) );
  NAND2_X1 U657 ( .A1(n14496), .A2(n5778), .ZN(n686) );
  NAND2_X1 U658 ( .A1(n14496), .A2(n5766), .ZN(n688) );
  NAND2_X1 U659 ( .A1(n14496), .A2(n5790), .ZN(n690) );
  NAND2_X1 U660 ( .A1(n14496), .A2(n5798), .ZN(n692) );
  NAND2_X1 U661 ( .A1(n14496), .A2(n5782), .ZN(n694) );
  NAND2_X1 U662 ( .A1(n14496), .A2(n5774), .ZN(n696) );
  NAND2_X1 U663 ( .A1(n14453), .A2(n5778), .ZN(n752) );
  NAND2_X1 U664 ( .A1(n14453), .A2(n5766), .ZN(n754) );
  NAND2_X1 U665 ( .A1(n14453), .A2(n5790), .ZN(n756) );
  NAND2_X1 U666 ( .A1(n14453), .A2(n5798), .ZN(n758) );
  NAND2_X1 U667 ( .A1(n14453), .A2(n5782), .ZN(n760) );
  NAND2_X1 U668 ( .A1(n14453), .A2(n5774), .ZN(n762) );
  NAND2_X1 U669 ( .A1(n14410), .A2(n5778), .ZN(n818) );
  NAND2_X1 U670 ( .A1(n14410), .A2(n5766), .ZN(n820) );
  NAND2_X1 U671 ( .A1(n14410), .A2(n5790), .ZN(n822) );
  NAND2_X1 U672 ( .A1(n14410), .A2(n5798), .ZN(n824) );
  NAND2_X1 U673 ( .A1(n14410), .A2(n5782), .ZN(n826) );
  NAND2_X1 U674 ( .A1(n14410), .A2(n5774), .ZN(n828) );
  NAND2_X1 U675 ( .A1(n14407), .A2(n5778), .ZN(n883) );
  NAND2_X1 U676 ( .A1(n14407), .A2(n5766), .ZN(n885) );
  NAND2_X1 U677 ( .A1(n14407), .A2(n5790), .ZN(n887) );
  NAND2_X1 U678 ( .A1(n14407), .A2(n5798), .ZN(n889) );
  NAND2_X1 U679 ( .A1(n14407), .A2(n5782), .ZN(n891) );
  NAND2_X1 U680 ( .A1(n14407), .A2(n5774), .ZN(n893) );
  NAND2_X1 U681 ( .A1(n14354), .A2(n5778), .ZN(n1014) );
  NAND2_X1 U682 ( .A1(n14354), .A2(n5766), .ZN(n1016) );
  NAND2_X1 U683 ( .A1(n14354), .A2(n5790), .ZN(n1018) );
  NAND2_X1 U684 ( .A1(n14354), .A2(n5798), .ZN(n1020) );
  NAND2_X1 U685 ( .A1(n14354), .A2(n5782), .ZN(n1022) );
  NAND2_X1 U686 ( .A1(n14354), .A2(n5774), .ZN(n1024) );
  NAND2_X1 U687 ( .A1(n14308), .A2(n5778), .ZN(n1156) );
  NAND2_X1 U688 ( .A1(n14308), .A2(n5766), .ZN(n1158) );
  NAND2_X1 U689 ( .A1(n14308), .A2(n5790), .ZN(n1160) );
  NAND2_X1 U690 ( .A1(n14308), .A2(n5798), .ZN(n1163) );
  NAND2_X1 U691 ( .A1(n14308), .A2(n5782), .ZN(n1166) );
  NAND2_X1 U692 ( .A1(n14308), .A2(n5774), .ZN(n1168) );
  NAND2_X1 U693 ( .A1(n14602), .A2(n5727), .ZN(n241) );
  NAND2_X1 U694 ( .A1(n14602), .A2(n5757), .ZN(n244) );
  NAND2_X1 U695 ( .A1(n14602), .A2(n5758), .ZN(n246) );
  NAND2_X1 U696 ( .A1(n14602), .A2(n5762), .ZN(n248) );
  NAND2_X1 U697 ( .A1(n14602), .A2(n5754), .ZN(n250) );
  NAND2_X1 U698 ( .A1(n14602), .A2(n5755), .ZN(n252) );
  NAND2_X1 U699 ( .A1(n14502), .A2(n5727), .ZN(n503) );
  NAND2_X1 U700 ( .A1(n14502), .A2(n5757), .ZN(n506) );
  NAND2_X1 U701 ( .A1(n14502), .A2(n5758), .ZN(n508) );
  NAND2_X1 U702 ( .A1(n14502), .A2(n5762), .ZN(n510) );
  NAND2_X1 U703 ( .A1(n14502), .A2(n5754), .ZN(n512) );
  NAND2_X1 U704 ( .A1(n14502), .A2(n5755), .ZN(n514) );
  NAND2_X1 U705 ( .A1(n14499), .A2(n5727), .ZN(n568) );
  NAND2_X1 U706 ( .A1(n14499), .A2(n5757), .ZN(n571) );
  NAND2_X1 U707 ( .A1(n14499), .A2(n5758), .ZN(n573) );
  NAND2_X1 U708 ( .A1(n14499), .A2(n5762), .ZN(n575) );
  NAND2_X1 U709 ( .A1(n14499), .A2(n5754), .ZN(n577) );
  NAND2_X1 U710 ( .A1(n14499), .A2(n5755), .ZN(n579) );
  NAND2_X1 U711 ( .A1(n14311), .A2(n5727), .ZN(n1027) );
  NAND2_X1 U712 ( .A1(n14311), .A2(n5757), .ZN(n1030) );
  NAND2_X1 U713 ( .A1(n14311), .A2(n5758), .ZN(n1032) );
  NAND2_X1 U714 ( .A1(n14311), .A2(n5762), .ZN(n1034) );
  NAND2_X1 U715 ( .A1(n14311), .A2(n5754), .ZN(n1036) );
  NAND2_X1 U716 ( .A1(n14311), .A2(n5755), .ZN(n1038) );
  NAND2_X1 U717 ( .A1(n14595), .A2(n5729), .ZN(n383) );
  NAND2_X1 U718 ( .A1(n14595), .A2(n5730), .ZN(n385) );
  NAND2_X1 U719 ( .A1(n14595), .A2(n5738), .ZN(n387) );
  NAND2_X1 U720 ( .A1(n14595), .A2(n5739), .ZN(n389) );
  NAND2_X1 U721 ( .A1(n14595), .A2(n5741), .ZN(n391) );
  NAND2_X1 U722 ( .A1(n14595), .A2(n5742), .ZN(n393) );
  NAND2_X1 U723 ( .A1(n14595), .A2(n5746), .ZN(n395) );
  NAND2_X1 U724 ( .A1(n5763), .A2(n14647), .ZN(n133) );
  NAND2_X1 U725 ( .A1(n5785), .A2(n14647), .ZN(n136) );
  NAND2_X1 U726 ( .A1(n5793), .A2(n14647), .ZN(n139) );
  NAND2_X1 U727 ( .A1(n5777), .A2(n14647), .ZN(n142) );
  NAND2_X1 U728 ( .A1(n5765), .A2(n14647), .ZN(n145) );
  NAND2_X1 U729 ( .A1(n5786), .A2(n14647), .ZN(n148) );
  NAND2_X1 U730 ( .A1(n5794), .A2(n14647), .ZN(n151) );
  NAND2_X1 U731 ( .A1(n5778), .A2(n14647), .ZN(n154) );
  NAND2_X1 U732 ( .A1(n5766), .A2(n14647), .ZN(n157) );
  NAND2_X1 U733 ( .A1(n5790), .A2(n14647), .ZN(n160) );
  NAND2_X1 U734 ( .A1(n5798), .A2(n14647), .ZN(n163) );
  NAND2_X1 U735 ( .A1(n5782), .A2(n14647), .ZN(n166) );
  NAND2_X1 U736 ( .A1(n5774), .A2(n14647), .ZN(n169) );
  NAND2_X1 U737 ( .A1(n5729), .A2(n14648), .ZN(n94) );
  NAND2_X1 U738 ( .A1(n5730), .A2(n14648), .ZN(n97) );
  NAND2_X1 U739 ( .A1(n5738), .A2(n14648), .ZN(n100) );
  NAND2_X1 U740 ( .A1(n5739), .A2(n14648), .ZN(n103) );
  NAND2_X1 U741 ( .A1(n5741), .A2(n14648), .ZN(n106) );
  NAND2_X1 U742 ( .A1(n5742), .A2(n14648), .ZN(n109) );
  NAND2_X1 U743 ( .A1(n5746), .A2(n14648), .ZN(n112) );
  NAND2_X1 U744 ( .A1(n5747), .A2(n14648), .ZN(n115) );
  NAND2_X1 U745 ( .A1(n5749), .A2(n14648), .ZN(n118) );
  NAND2_X1 U746 ( .A1(n5750), .A2(n14648), .ZN(n121) );
  NAND2_X1 U747 ( .A1(n5783), .A2(n14648), .ZN(n124) );
  NAND2_X1 U748 ( .A1(n5791), .A2(n14648), .ZN(n127) );
  NAND2_X1 U749 ( .A1(n5775), .A2(n14648), .ZN(n130) );
  NAND2_X1 U750 ( .A1(n14603), .A2(n5727), .ZN(n174) );
  NAND2_X1 U751 ( .A1(n14603), .A2(n5757), .ZN(n177) );
  NAND2_X1 U752 ( .A1(n14603), .A2(n5758), .ZN(n179) );
  NAND2_X1 U753 ( .A1(n14603), .A2(n5762), .ZN(n181) );
  NAND2_X1 U754 ( .A1(n14603), .A2(n5754), .ZN(n183) );
  NAND2_X1 U755 ( .A1(n14603), .A2(n5755), .ZN(n185) );
  NAND2_X1 U756 ( .A1(n14603), .A2(n5729), .ZN(n187) );
  NAND2_X1 U757 ( .A1(n14603), .A2(n5730), .ZN(n189) );
  NAND2_X1 U758 ( .A1(n14603), .A2(n5738), .ZN(n191) );
  NAND2_X1 U759 ( .A1(n14603), .A2(n5739), .ZN(n193) );
  NAND2_X1 U760 ( .A1(n14603), .A2(n5741), .ZN(n195) );
  NAND2_X1 U761 ( .A1(n14603), .A2(n5742), .ZN(n197) );
  NAND2_X1 U762 ( .A1(n14603), .A2(n5746), .ZN(n199) );
  NAND2_X1 U763 ( .A1(n14604), .A2(n5747), .ZN(n201) );
  NAND2_X1 U764 ( .A1(n14604), .A2(n5749), .ZN(n203) );
  NAND2_X1 U765 ( .A1(n14604), .A2(n5750), .ZN(n205) );
  NAND2_X1 U766 ( .A1(n14604), .A2(n5783), .ZN(n207) );
  NAND2_X1 U767 ( .A1(n14604), .A2(n5791), .ZN(n209) );
  NAND2_X1 U768 ( .A1(n14604), .A2(n5775), .ZN(n211) );
  NAND2_X1 U769 ( .A1(n14604), .A2(n5763), .ZN(n213) );
  NAND2_X1 U770 ( .A1(n14604), .A2(n5785), .ZN(n215) );
  NAND2_X1 U771 ( .A1(n14604), .A2(n5793), .ZN(n217) );
  NAND2_X1 U772 ( .A1(n14604), .A2(n5777), .ZN(n219) );
  NAND2_X1 U773 ( .A1(n14604), .A2(n5765), .ZN(n221) );
  NAND2_X1 U774 ( .A1(n14604), .A2(n5786), .ZN(n223) );
  NAND2_X1 U775 ( .A1(n14604), .A2(n5794), .ZN(n225) );
  NAND2_X1 U776 ( .A1(n14601), .A2(n5729), .ZN(n254) );
  NAND2_X1 U777 ( .A1(n14601), .A2(n5730), .ZN(n256) );
  NAND2_X1 U778 ( .A1(n14601), .A2(n5738), .ZN(n258) );
  NAND2_X1 U779 ( .A1(n14601), .A2(n5739), .ZN(n260) );
  NAND2_X1 U780 ( .A1(n14601), .A2(n5741), .ZN(n262) );
  NAND2_X1 U781 ( .A1(n14601), .A2(n5742), .ZN(n264) );
  NAND2_X1 U782 ( .A1(n14601), .A2(n5746), .ZN(n266) );
  NAND2_X1 U783 ( .A1(n14601), .A2(n5747), .ZN(n268) );
  NAND2_X1 U784 ( .A1(n14601), .A2(n5749), .ZN(n270) );
  NAND2_X1 U785 ( .A1(n14601), .A2(n5750), .ZN(n272) );
  NAND2_X1 U786 ( .A1(n14601), .A2(n5783), .ZN(n274) );
  NAND2_X1 U787 ( .A1(n14601), .A2(n5791), .ZN(n276) );
  NAND2_X1 U788 ( .A1(n14601), .A2(n5775), .ZN(n278) );
  NAND2_X1 U789 ( .A1(n14600), .A2(n5763), .ZN(n280) );
  NAND2_X1 U790 ( .A1(n14600), .A2(n5785), .ZN(n282) );
  NAND2_X1 U791 ( .A1(n14600), .A2(n5793), .ZN(n284) );
  NAND2_X1 U792 ( .A1(n14600), .A2(n5777), .ZN(n286) );
  NAND2_X1 U793 ( .A1(n14600), .A2(n5765), .ZN(n288) );
  NAND2_X1 U794 ( .A1(n14600), .A2(n5786), .ZN(n290) );
  NAND2_X1 U795 ( .A1(n14600), .A2(n5794), .ZN(n292) );
  NAND2_X1 U796 ( .A1(n14600), .A2(n5778), .ZN(n294) );
  NAND2_X1 U797 ( .A1(n14600), .A2(n5766), .ZN(n296) );
  NAND2_X1 U798 ( .A1(n14600), .A2(n5790), .ZN(n298) );
  NAND2_X1 U799 ( .A1(n14600), .A2(n5798), .ZN(n300) );
  NAND2_X1 U800 ( .A1(n14600), .A2(n5782), .ZN(n302) );
  NAND2_X1 U801 ( .A1(n14600), .A2(n5774), .ZN(n304) );
  NAND2_X1 U802 ( .A1(n14597), .A2(n5727), .ZN(n306) );
  NAND2_X1 U803 ( .A1(n14597), .A2(n5757), .ZN(n309) );
  NAND2_X1 U804 ( .A1(n14597), .A2(n5758), .ZN(n311) );
  NAND2_X1 U805 ( .A1(n14597), .A2(n5762), .ZN(n313) );
  NAND2_X1 U806 ( .A1(n14597), .A2(n5754), .ZN(n315) );
  NAND2_X1 U807 ( .A1(n14597), .A2(n5755), .ZN(n317) );
  NAND2_X1 U808 ( .A1(n14597), .A2(n5729), .ZN(n319) );
  NAND2_X1 U809 ( .A1(n14597), .A2(n5730), .ZN(n321) );
  NAND2_X1 U810 ( .A1(n14597), .A2(n5738), .ZN(n323) );
  NAND2_X1 U811 ( .A1(n14597), .A2(n5739), .ZN(n325) );
  NAND2_X1 U812 ( .A1(n14597), .A2(n5741), .ZN(n327) );
  NAND2_X1 U813 ( .A1(n14597), .A2(n5742), .ZN(n329) );
  NAND2_X1 U814 ( .A1(n14597), .A2(n5746), .ZN(n331) );
  NAND2_X1 U815 ( .A1(n14598), .A2(n5747), .ZN(n333) );
  NAND2_X1 U816 ( .A1(n14598), .A2(n5749), .ZN(n335) );
  NAND2_X1 U817 ( .A1(n14598), .A2(n5750), .ZN(n337) );
  NAND2_X1 U818 ( .A1(n14598), .A2(n5783), .ZN(n339) );
  NAND2_X1 U819 ( .A1(n14598), .A2(n5791), .ZN(n341) );
  NAND2_X1 U820 ( .A1(n14598), .A2(n5775), .ZN(n343) );
  NAND2_X1 U821 ( .A1(n14598), .A2(n5763), .ZN(n345) );
  NAND2_X1 U822 ( .A1(n14598), .A2(n5785), .ZN(n347) );
  NAND2_X1 U823 ( .A1(n14598), .A2(n5793), .ZN(n349) );
  NAND2_X1 U824 ( .A1(n14598), .A2(n5777), .ZN(n351) );
  NAND2_X1 U825 ( .A1(n14598), .A2(n5765), .ZN(n353) );
  NAND2_X1 U826 ( .A1(n14598), .A2(n5786), .ZN(n355) );
  NAND2_X1 U827 ( .A1(n14598), .A2(n5794), .ZN(n357) );
  NAND2_X1 U828 ( .A1(n14595), .A2(n5747), .ZN(n398) );
  NAND2_X1 U829 ( .A1(n14595), .A2(n5749), .ZN(n400) );
  NAND2_X1 U830 ( .A1(n14595), .A2(n5750), .ZN(n402) );
  NAND2_X1 U831 ( .A1(n14595), .A2(n5783), .ZN(n404) );
  NAND2_X1 U832 ( .A1(n14595), .A2(n5791), .ZN(n406) );
  NAND2_X1 U833 ( .A1(n14595), .A2(n5775), .ZN(n408) );
  NAND2_X1 U834 ( .A1(n14594), .A2(n5763), .ZN(n410) );
  NAND2_X1 U835 ( .A1(n14594), .A2(n5785), .ZN(n412) );
  NAND2_X1 U836 ( .A1(n14594), .A2(n5793), .ZN(n414) );
  NAND2_X1 U837 ( .A1(n14594), .A2(n5777), .ZN(n416) );
  NAND2_X1 U838 ( .A1(n14594), .A2(n5765), .ZN(n418) );
  NAND2_X1 U839 ( .A1(n14594), .A2(n5786), .ZN(n420) );
  NAND2_X1 U840 ( .A1(n14594), .A2(n5794), .ZN(n422) );
  NAND2_X1 U841 ( .A1(n14594), .A2(n5778), .ZN(n424) );
  NAND2_X1 U842 ( .A1(n14594), .A2(n5766), .ZN(n426) );
  NAND2_X1 U843 ( .A1(n14594), .A2(n5790), .ZN(n428) );
  NAND2_X1 U844 ( .A1(n14594), .A2(n5798), .ZN(n430) );
  NAND2_X1 U845 ( .A1(n14594), .A2(n5782), .ZN(n432) );
  NAND2_X1 U846 ( .A1(n14594), .A2(n5774), .ZN(n434) );
  NAND2_X1 U847 ( .A1(n14550), .A2(n5729), .ZN(n450) );
  NAND2_X1 U848 ( .A1(n14550), .A2(n5730), .ZN(n452) );
  NAND2_X1 U849 ( .A1(n14550), .A2(n5738), .ZN(n454) );
  NAND2_X1 U850 ( .A1(n14550), .A2(n5739), .ZN(n456) );
  NAND2_X1 U851 ( .A1(n14550), .A2(n5741), .ZN(n458) );
  NAND2_X1 U852 ( .A1(n14550), .A2(n5742), .ZN(n460) );
  NAND2_X1 U853 ( .A1(n14550), .A2(n5746), .ZN(n462) );
  NAND2_X1 U854 ( .A1(n14550), .A2(n5747), .ZN(n464) );
  NAND2_X1 U855 ( .A1(n14550), .A2(n5749), .ZN(n466) );
  NAND2_X1 U856 ( .A1(n14550), .A2(n5750), .ZN(n468) );
  NAND2_X1 U857 ( .A1(n14550), .A2(n5783), .ZN(n470) );
  NAND2_X1 U858 ( .A1(n14550), .A2(n5791), .ZN(n472) );
  NAND2_X1 U859 ( .A1(n14550), .A2(n5775), .ZN(n474) );
  NAND2_X1 U860 ( .A1(n14549), .A2(n5763), .ZN(n476) );
  NAND2_X1 U861 ( .A1(n14549), .A2(n5785), .ZN(n478) );
  NAND2_X1 U862 ( .A1(n14549), .A2(n5793), .ZN(n480) );
  NAND2_X1 U863 ( .A1(n14549), .A2(n5777), .ZN(n482) );
  NAND2_X1 U864 ( .A1(n14549), .A2(n5765), .ZN(n484) );
  NAND2_X1 U865 ( .A1(n14549), .A2(n5786), .ZN(n486) );
  NAND2_X1 U866 ( .A1(n14549), .A2(n5794), .ZN(n488) );
  NAND2_X1 U867 ( .A1(n14549), .A2(n5778), .ZN(n490) );
  NAND2_X1 U868 ( .A1(n14549), .A2(n5766), .ZN(n492) );
  NAND2_X1 U869 ( .A1(n14549), .A2(n5790), .ZN(n494) );
  NAND2_X1 U870 ( .A1(n14549), .A2(n5798), .ZN(n496) );
  NAND2_X1 U871 ( .A1(n14549), .A2(n5782), .ZN(n498) );
  NAND2_X1 U872 ( .A1(n14549), .A2(n5774), .ZN(n500) );
  NAND2_X1 U873 ( .A1(n14501), .A2(n5729), .ZN(n516) );
  NAND2_X1 U874 ( .A1(n14501), .A2(n5730), .ZN(n518) );
  NAND2_X1 U875 ( .A1(n14501), .A2(n5738), .ZN(n520) );
  NAND2_X1 U876 ( .A1(n14501), .A2(n5739), .ZN(n522) );
  NAND2_X1 U877 ( .A1(n14501), .A2(n5741), .ZN(n524) );
  NAND2_X1 U878 ( .A1(n14501), .A2(n5742), .ZN(n526) );
  NAND2_X1 U879 ( .A1(n14501), .A2(n5746), .ZN(n528) );
  NAND2_X1 U880 ( .A1(n14501), .A2(n5747), .ZN(n530) );
  NAND2_X1 U881 ( .A1(n14501), .A2(n5749), .ZN(n532) );
  NAND2_X1 U882 ( .A1(n14501), .A2(n5750), .ZN(n534) );
  NAND2_X1 U883 ( .A1(n14501), .A2(n5783), .ZN(n536) );
  NAND2_X1 U884 ( .A1(n14501), .A2(n5791), .ZN(n538) );
  NAND2_X1 U885 ( .A1(n14501), .A2(n5775), .ZN(n540) );
  NAND2_X1 U886 ( .A1(n14500), .A2(n5763), .ZN(n542) );
  NAND2_X1 U887 ( .A1(n14500), .A2(n5785), .ZN(n544) );
  NAND2_X1 U888 ( .A1(n14500), .A2(n5793), .ZN(n546) );
  NAND2_X1 U889 ( .A1(n14500), .A2(n5777), .ZN(n548) );
  NAND2_X1 U890 ( .A1(n14500), .A2(n5765), .ZN(n550) );
  NAND2_X1 U891 ( .A1(n14500), .A2(n5786), .ZN(n552) );
  NAND2_X1 U892 ( .A1(n14500), .A2(n5794), .ZN(n554) );
  NAND2_X1 U893 ( .A1(n14500), .A2(n5778), .ZN(n556) );
  NAND2_X1 U894 ( .A1(n14500), .A2(n5766), .ZN(n558) );
  NAND2_X1 U895 ( .A1(n14500), .A2(n5790), .ZN(n560) );
  NAND2_X1 U896 ( .A1(n14500), .A2(n5798), .ZN(n562) );
  NAND2_X1 U897 ( .A1(n14500), .A2(n5782), .ZN(n564) );
  NAND2_X1 U898 ( .A1(n14500), .A2(n5774), .ZN(n566) );
  NAND2_X1 U899 ( .A1(n14498), .A2(n5729), .ZN(n581) );
  NAND2_X1 U900 ( .A1(n14498), .A2(n5730), .ZN(n583) );
  NAND2_X1 U901 ( .A1(n14498), .A2(n5738), .ZN(n585) );
  NAND2_X1 U902 ( .A1(n14498), .A2(n5739), .ZN(n587) );
  NAND2_X1 U903 ( .A1(n14498), .A2(n5741), .ZN(n589) );
  NAND2_X1 U904 ( .A1(n14498), .A2(n5742), .ZN(n591) );
  NAND2_X1 U905 ( .A1(n14498), .A2(n5746), .ZN(n593) );
  NAND2_X1 U906 ( .A1(n14498), .A2(n5747), .ZN(n595) );
  NAND2_X1 U907 ( .A1(n14498), .A2(n5749), .ZN(n597) );
  NAND2_X1 U908 ( .A1(n14498), .A2(n5750), .ZN(n599) );
  NAND2_X1 U909 ( .A1(n14498), .A2(n5783), .ZN(n601) );
  NAND2_X1 U910 ( .A1(n14498), .A2(n5791), .ZN(n603) );
  NAND2_X1 U911 ( .A1(n14498), .A2(n5775), .ZN(n605) );
  NAND2_X1 U912 ( .A1(n14497), .A2(n5763), .ZN(n607) );
  NAND2_X1 U913 ( .A1(n14497), .A2(n5785), .ZN(n609) );
  NAND2_X1 U914 ( .A1(n14497), .A2(n5793), .ZN(n611) );
  NAND2_X1 U915 ( .A1(n14497), .A2(n5777), .ZN(n613) );
  NAND2_X1 U916 ( .A1(n14497), .A2(n5765), .ZN(n615) );
  NAND2_X1 U917 ( .A1(n14497), .A2(n5786), .ZN(n617) );
  NAND2_X1 U918 ( .A1(n14497), .A2(n5794), .ZN(n619) );
  NAND2_X1 U919 ( .A1(n14497), .A2(n5778), .ZN(n621) );
  NAND2_X1 U920 ( .A1(n14497), .A2(n5766), .ZN(n623) );
  NAND2_X1 U921 ( .A1(n14497), .A2(n5790), .ZN(n625) );
  NAND2_X1 U922 ( .A1(n14497), .A2(n5798), .ZN(n627) );
  NAND2_X1 U923 ( .A1(n14497), .A2(n5782), .ZN(n629) );
  NAND2_X1 U924 ( .A1(n14497), .A2(n5774), .ZN(n631) );
  NAND2_X1 U925 ( .A1(n14494), .A2(n5727), .ZN(n633) );
  NAND2_X1 U926 ( .A1(n14494), .A2(n5757), .ZN(n636) );
  NAND2_X1 U927 ( .A1(n14494), .A2(n5758), .ZN(n638) );
  NAND2_X1 U928 ( .A1(n14494), .A2(n5762), .ZN(n640) );
  NAND2_X1 U929 ( .A1(n14494), .A2(n5754), .ZN(n642) );
  NAND2_X1 U930 ( .A1(n14494), .A2(n5755), .ZN(n644) );
  NAND2_X1 U931 ( .A1(n14494), .A2(n5729), .ZN(n646) );
  NAND2_X1 U932 ( .A1(n14494), .A2(n5730), .ZN(n648) );
  NAND2_X1 U933 ( .A1(n14494), .A2(n5738), .ZN(n650) );
  NAND2_X1 U934 ( .A1(n14494), .A2(n5739), .ZN(n652) );
  NAND2_X1 U935 ( .A1(n14494), .A2(n5741), .ZN(n654) );
  NAND2_X1 U936 ( .A1(n14494), .A2(n5742), .ZN(n656) );
  NAND2_X1 U937 ( .A1(n14494), .A2(n5746), .ZN(n658) );
  NAND2_X1 U938 ( .A1(n14495), .A2(n5747), .ZN(n660) );
  NAND2_X1 U939 ( .A1(n14495), .A2(n5749), .ZN(n662) );
  NAND2_X1 U940 ( .A1(n14495), .A2(n5750), .ZN(n664) );
  NAND2_X1 U941 ( .A1(n14495), .A2(n5783), .ZN(n666) );
  NAND2_X1 U942 ( .A1(n14495), .A2(n5791), .ZN(n668) );
  NAND2_X1 U943 ( .A1(n14495), .A2(n5775), .ZN(n670) );
  NAND2_X1 U944 ( .A1(n14495), .A2(n5763), .ZN(n672) );
  NAND2_X1 U945 ( .A1(n14495), .A2(n5785), .ZN(n674) );
  NAND2_X1 U946 ( .A1(n14495), .A2(n5793), .ZN(n676) );
  NAND2_X1 U947 ( .A1(n14495), .A2(n5777), .ZN(n678) );
  NAND2_X1 U948 ( .A1(n14495), .A2(n5765), .ZN(n680) );
  NAND2_X1 U949 ( .A1(n14495), .A2(n5786), .ZN(n682) );
  NAND2_X1 U950 ( .A1(n14495), .A2(n5794), .ZN(n684) );
  NAND2_X1 U951 ( .A1(n14451), .A2(n5727), .ZN(n699) );
  NAND2_X1 U952 ( .A1(n14451), .A2(n5757), .ZN(n702) );
  NAND2_X1 U953 ( .A1(n14451), .A2(n5758), .ZN(n704) );
  NAND2_X1 U954 ( .A1(n14451), .A2(n5762), .ZN(n706) );
  NAND2_X1 U955 ( .A1(n14451), .A2(n5754), .ZN(n708) );
  NAND2_X1 U956 ( .A1(n14451), .A2(n5755), .ZN(n710) );
  NAND2_X1 U957 ( .A1(n14451), .A2(n5729), .ZN(n712) );
  NAND2_X1 U958 ( .A1(n14451), .A2(n5730), .ZN(n714) );
  NAND2_X1 U959 ( .A1(n14451), .A2(n5738), .ZN(n716) );
  NAND2_X1 U960 ( .A1(n14451), .A2(n5739), .ZN(n718) );
  NAND2_X1 U961 ( .A1(n14451), .A2(n5741), .ZN(n720) );
  NAND2_X1 U962 ( .A1(n14451), .A2(n5742), .ZN(n722) );
  NAND2_X1 U963 ( .A1(n14451), .A2(n5746), .ZN(n724) );
  NAND2_X1 U964 ( .A1(n14452), .A2(n5747), .ZN(n726) );
  NAND2_X1 U965 ( .A1(n14452), .A2(n5749), .ZN(n728) );
  NAND2_X1 U966 ( .A1(n14452), .A2(n5750), .ZN(n730) );
  NAND2_X1 U967 ( .A1(n14452), .A2(n5783), .ZN(n732) );
  NAND2_X1 U968 ( .A1(n14452), .A2(n5791), .ZN(n734) );
  NAND2_X1 U969 ( .A1(n14452), .A2(n5775), .ZN(n736) );
  NAND2_X1 U970 ( .A1(n14452), .A2(n5763), .ZN(n738) );
  NAND2_X1 U971 ( .A1(n14452), .A2(n5785), .ZN(n740) );
  NAND2_X1 U972 ( .A1(n14452), .A2(n5793), .ZN(n742) );
  NAND2_X1 U973 ( .A1(n14452), .A2(n5777), .ZN(n744) );
  NAND2_X1 U974 ( .A1(n14452), .A2(n5765), .ZN(n746) );
  NAND2_X1 U975 ( .A1(n14452), .A2(n5786), .ZN(n748) );
  NAND2_X1 U976 ( .A1(n14452), .A2(n5794), .ZN(n750) );
  NAND2_X1 U977 ( .A1(n14408), .A2(n5727), .ZN(n765) );
  NAND2_X1 U978 ( .A1(n14408), .A2(n5757), .ZN(n768) );
  NAND2_X1 U979 ( .A1(n14408), .A2(n5758), .ZN(n770) );
  NAND2_X1 U980 ( .A1(n14408), .A2(n5762), .ZN(n772) );
  NAND2_X1 U981 ( .A1(n14408), .A2(n5754), .ZN(n774) );
  NAND2_X1 U982 ( .A1(n14408), .A2(n5755), .ZN(n776) );
  NAND2_X1 U983 ( .A1(n14408), .A2(n5729), .ZN(n778) );
  NAND2_X1 U984 ( .A1(n14408), .A2(n5730), .ZN(n780) );
  NAND2_X1 U985 ( .A1(n14408), .A2(n5738), .ZN(n782) );
  NAND2_X1 U986 ( .A1(n14408), .A2(n5739), .ZN(n784) );
  NAND2_X1 U987 ( .A1(n14408), .A2(n5741), .ZN(n786) );
  NAND2_X1 U988 ( .A1(n14408), .A2(n5742), .ZN(n788) );
  NAND2_X1 U989 ( .A1(n14408), .A2(n5746), .ZN(n790) );
  NAND2_X1 U990 ( .A1(n14409), .A2(n5747), .ZN(n792) );
  NAND2_X1 U991 ( .A1(n14409), .A2(n5749), .ZN(n794) );
  NAND2_X1 U992 ( .A1(n14409), .A2(n5750), .ZN(n796) );
  NAND2_X1 U993 ( .A1(n14409), .A2(n5783), .ZN(n798) );
  NAND2_X1 U994 ( .A1(n14409), .A2(n5791), .ZN(n800) );
  NAND2_X1 U995 ( .A1(n14409), .A2(n5775), .ZN(n802) );
  NAND2_X1 U996 ( .A1(n14409), .A2(n5763), .ZN(n804) );
  NAND2_X1 U997 ( .A1(n14409), .A2(n5785), .ZN(n806) );
  NAND2_X1 U998 ( .A1(n14409), .A2(n5793), .ZN(n808) );
  NAND2_X1 U999 ( .A1(n14409), .A2(n5777), .ZN(n810) );
  NAND2_X1 U1000 ( .A1(n14409), .A2(n5765), .ZN(n812) );
  NAND2_X1 U1001 ( .A1(n14409), .A2(n5786), .ZN(n814) );
  NAND2_X1 U1002 ( .A1(n14409), .A2(n5794), .ZN(n816) );
  NAND2_X1 U1003 ( .A1(n14405), .A2(n5727), .ZN(n830) );
  NAND2_X1 U1004 ( .A1(n14405), .A2(n5757), .ZN(n833) );
  NAND2_X1 U1005 ( .A1(n14405), .A2(n5758), .ZN(n835) );
  NAND2_X1 U1006 ( .A1(n14405), .A2(n5762), .ZN(n837) );
  NAND2_X1 U1007 ( .A1(n14405), .A2(n5754), .ZN(n839) );
  NAND2_X1 U1008 ( .A1(n14405), .A2(n5755), .ZN(n841) );
  NAND2_X1 U1009 ( .A1(n14405), .A2(n5729), .ZN(n843) );
  NAND2_X1 U1010 ( .A1(n14405), .A2(n5730), .ZN(n845) );
  NAND2_X1 U1011 ( .A1(n14405), .A2(n5738), .ZN(n847) );
  NAND2_X1 U1012 ( .A1(n14405), .A2(n5739), .ZN(n849) );
  NAND2_X1 U1013 ( .A1(n14405), .A2(n5741), .ZN(n851) );
  NAND2_X1 U1014 ( .A1(n14405), .A2(n5742), .ZN(n853) );
  NAND2_X1 U1015 ( .A1(n14405), .A2(n5746), .ZN(n855) );
  NAND2_X1 U1016 ( .A1(n14406), .A2(n5747), .ZN(n857) );
  NAND2_X1 U1017 ( .A1(n14406), .A2(n5749), .ZN(n859) );
  NAND2_X1 U1018 ( .A1(n14406), .A2(n5750), .ZN(n861) );
  NAND2_X1 U1019 ( .A1(n14406), .A2(n5783), .ZN(n863) );
  NAND2_X1 U1020 ( .A1(n14406), .A2(n5791), .ZN(n865) );
  NAND2_X1 U1021 ( .A1(n14406), .A2(n5775), .ZN(n867) );
  NAND2_X1 U1022 ( .A1(n14406), .A2(n5763), .ZN(n869) );
  NAND2_X1 U1023 ( .A1(n14406), .A2(n5785), .ZN(n871) );
  NAND2_X1 U1024 ( .A1(n14406), .A2(n5793), .ZN(n873) );
  NAND2_X1 U1025 ( .A1(n14406), .A2(n5777), .ZN(n875) );
  NAND2_X1 U1026 ( .A1(n14406), .A2(n5765), .ZN(n877) );
  NAND2_X1 U1027 ( .A1(n14406), .A2(n5786), .ZN(n879) );
  NAND2_X1 U1028 ( .A1(n14406), .A2(n5794), .ZN(n881) );
  NAND2_X1 U1029 ( .A1(n14402), .A2(n5729), .ZN(n908) );
  NAND2_X1 U1030 ( .A1(n14402), .A2(n5730), .ZN(n910) );
  NAND2_X1 U1031 ( .A1(n14402), .A2(n5738), .ZN(n912) );
  NAND2_X1 U1032 ( .A1(n14402), .A2(n5739), .ZN(n914) );
  NAND2_X1 U1033 ( .A1(n14402), .A2(n5741), .ZN(n916) );
  NAND2_X1 U1034 ( .A1(n14402), .A2(n5742), .ZN(n918) );
  NAND2_X1 U1035 ( .A1(n14402), .A2(n5746), .ZN(n920) );
  NAND2_X1 U1036 ( .A1(n14402), .A2(n5747), .ZN(n922) );
  NAND2_X1 U1037 ( .A1(n14402), .A2(n5749), .ZN(n924) );
  NAND2_X1 U1038 ( .A1(n14402), .A2(n5750), .ZN(n926) );
  NAND2_X1 U1039 ( .A1(n14402), .A2(n5783), .ZN(n928) );
  NAND2_X1 U1040 ( .A1(n14402), .A2(n5791), .ZN(n930) );
  NAND2_X1 U1041 ( .A1(n14402), .A2(n5775), .ZN(n932) );
  NAND2_X1 U1042 ( .A1(n14401), .A2(n5763), .ZN(n934) );
  NAND2_X1 U1043 ( .A1(n14401), .A2(n5785), .ZN(n936) );
  NAND2_X1 U1044 ( .A1(n14401), .A2(n5793), .ZN(n938) );
  NAND2_X1 U1045 ( .A1(n14401), .A2(n5777), .ZN(n940) );
  NAND2_X1 U1046 ( .A1(n14401), .A2(n5765), .ZN(n942) );
  NAND2_X1 U1047 ( .A1(n14401), .A2(n5786), .ZN(n944) );
  NAND2_X1 U1048 ( .A1(n14401), .A2(n5794), .ZN(n946) );
  NAND2_X1 U1049 ( .A1(n14401), .A2(n5778), .ZN(n948) );
  NAND2_X1 U1050 ( .A1(n14401), .A2(n5766), .ZN(n950) );
  NAND2_X1 U1051 ( .A1(n14401), .A2(n5790), .ZN(n952) );
  NAND2_X1 U1052 ( .A1(n14401), .A2(n5798), .ZN(n954) );
  NAND2_X1 U1053 ( .A1(n14401), .A2(n5782), .ZN(n956) );
  NAND2_X1 U1054 ( .A1(n14401), .A2(n5774), .ZN(n958) );
  NAND2_X1 U1055 ( .A1(n14352), .A2(n5727), .ZN(n961) );
  NAND2_X1 U1056 ( .A1(n14352), .A2(n5757), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(n14352), .A2(n5758), .ZN(n966) );
  NAND2_X1 U1058 ( .A1(n14352), .A2(n5762), .ZN(n968) );
  NAND2_X1 U1059 ( .A1(n14352), .A2(n5754), .ZN(n970) );
  NAND2_X1 U1060 ( .A1(n14352), .A2(n5755), .ZN(n972) );
  NAND2_X1 U1061 ( .A1(n14352), .A2(n5729), .ZN(n974) );
  NAND2_X1 U1062 ( .A1(n14352), .A2(n5730), .ZN(n976) );
  NAND2_X1 U1063 ( .A1(n14352), .A2(n5738), .ZN(n978) );
  NAND2_X1 U1064 ( .A1(n14352), .A2(n5739), .ZN(n980) );
  NAND2_X1 U1065 ( .A1(n14352), .A2(n5741), .ZN(n982) );
  NAND2_X1 U1066 ( .A1(n14352), .A2(n5742), .ZN(n984) );
  NAND2_X1 U1067 ( .A1(n14352), .A2(n5746), .ZN(n986) );
  NAND2_X1 U1068 ( .A1(n14353), .A2(n5747), .ZN(n988) );
  NAND2_X1 U1069 ( .A1(n14353), .A2(n5749), .ZN(n990) );
  NAND2_X1 U1070 ( .A1(n14353), .A2(n5750), .ZN(n992) );
  NAND2_X1 U1071 ( .A1(n14353), .A2(n5783), .ZN(n994) );
  NAND2_X1 U1072 ( .A1(n14353), .A2(n5791), .ZN(n996) );
  NAND2_X1 U1073 ( .A1(n14353), .A2(n5775), .ZN(n998) );
  NAND2_X1 U1074 ( .A1(n14353), .A2(n5763), .ZN(n1000) );
  NAND2_X1 U1075 ( .A1(n14353), .A2(n5785), .ZN(n1002) );
  NAND2_X1 U1076 ( .A1(n14353), .A2(n5793), .ZN(n1004) );
  NAND2_X1 U1077 ( .A1(n14353), .A2(n5777), .ZN(n1006) );
  NAND2_X1 U1078 ( .A1(n14353), .A2(n5765), .ZN(n1008) );
  NAND2_X1 U1079 ( .A1(n14353), .A2(n5786), .ZN(n1010) );
  NAND2_X1 U1080 ( .A1(n14353), .A2(n5794), .ZN(n1012) );
  NAND2_X1 U1081 ( .A1(n14310), .A2(n5729), .ZN(n1040) );
  NAND2_X1 U1082 ( .A1(n14310), .A2(n5730), .ZN(n1042) );
  NAND2_X1 U1083 ( .A1(n14310), .A2(n5738), .ZN(n1044) );
  NAND2_X1 U1084 ( .A1(n14310), .A2(n5739), .ZN(n1046) );
  NAND2_X1 U1085 ( .A1(n14310), .A2(n5741), .ZN(n1048) );
  NAND2_X1 U1086 ( .A1(n14310), .A2(n5742), .ZN(n1050) );
  NAND2_X1 U1087 ( .A1(n14310), .A2(n5746), .ZN(n1052) );
  NAND2_X1 U1088 ( .A1(n14310), .A2(n5747), .ZN(n1054) );
  NAND2_X1 U1089 ( .A1(n14310), .A2(n5749), .ZN(n1056) );
  NAND2_X1 U1090 ( .A1(n14310), .A2(n5750), .ZN(n1058) );
  NAND2_X1 U1091 ( .A1(n14310), .A2(n5783), .ZN(n1060) );
  NAND2_X1 U1092 ( .A1(n14310), .A2(n5791), .ZN(n1062) );
  NAND2_X1 U1093 ( .A1(n14310), .A2(n5775), .ZN(n1064) );
  NAND2_X1 U1094 ( .A1(n14309), .A2(n5763), .ZN(n1066) );
  NAND2_X1 U1095 ( .A1(n14309), .A2(n5785), .ZN(n1068) );
  NAND2_X1 U1096 ( .A1(n14309), .A2(n5793), .ZN(n1070) );
  NAND2_X1 U1097 ( .A1(n14309), .A2(n5777), .ZN(n1072) );
  NAND2_X1 U1098 ( .A1(n14309), .A2(n5765), .ZN(n1074) );
  NAND2_X1 U1099 ( .A1(n14309), .A2(n5786), .ZN(n1076) );
  NAND2_X1 U1100 ( .A1(n14309), .A2(n5794), .ZN(n1078) );
  NAND2_X1 U1101 ( .A1(n14309), .A2(n5778), .ZN(n1080) );
  NAND2_X1 U1102 ( .A1(n14309), .A2(n5766), .ZN(n1082) );
  NAND2_X1 U1103 ( .A1(n14309), .A2(n5790), .ZN(n1084) );
  NAND2_X1 U1104 ( .A1(n14309), .A2(n5798), .ZN(n1086) );
  NAND2_X1 U1105 ( .A1(n14309), .A2(n5782), .ZN(n1088) );
  NAND2_X1 U1106 ( .A1(n14309), .A2(n5774), .ZN(n1090) );
  NAND2_X1 U1107 ( .A1(n14306), .A2(n5727), .ZN(n1092) );
  NAND2_X1 U1108 ( .A1(n14306), .A2(n5757), .ZN(n1097) );
  NAND2_X1 U1109 ( .A1(n14306), .A2(n5758), .ZN(n1100) );
  NAND2_X1 U1110 ( .A1(n14306), .A2(n5762), .ZN(n1103) );
  NAND2_X1 U1111 ( .A1(n14306), .A2(n5754), .ZN(n1106) );
  NAND2_X1 U1112 ( .A1(n14306), .A2(n5755), .ZN(n1109) );
  NAND2_X1 U1113 ( .A1(n14306), .A2(n5729), .ZN(n1111) );
  NAND2_X1 U1114 ( .A1(n14306), .A2(n5730), .ZN(n1113) );
  NAND2_X1 U1115 ( .A1(n14306), .A2(n5738), .ZN(n1115) );
  NAND2_X1 U1116 ( .A1(n14306), .A2(n5739), .ZN(n1118) );
  NAND2_X1 U1117 ( .A1(n14306), .A2(n5741), .ZN(n1120) );
  NAND2_X1 U1118 ( .A1(n14306), .A2(n5742), .ZN(n1122) );
  NAND2_X1 U1119 ( .A1(n14306), .A2(n5746), .ZN(n1124) );
  NAND2_X1 U1120 ( .A1(n14307), .A2(n5747), .ZN(n1127) );
  NAND2_X1 U1121 ( .A1(n14307), .A2(n5749), .ZN(n1129) );
  NAND2_X1 U1122 ( .A1(n14307), .A2(n5750), .ZN(n1131) );
  NAND2_X1 U1123 ( .A1(n14307), .A2(n5783), .ZN(n1133) );
  NAND2_X1 U1124 ( .A1(n14307), .A2(n5791), .ZN(n1136) );
  NAND2_X1 U1125 ( .A1(n14307), .A2(n5775), .ZN(n1138) );
  NAND2_X1 U1126 ( .A1(n14307), .A2(n5763), .ZN(n1140) );
  NAND2_X1 U1127 ( .A1(n14307), .A2(n5785), .ZN(n1142) );
  NAND2_X1 U1128 ( .A1(n14307), .A2(n5793), .ZN(n1145) );
  NAND2_X1 U1129 ( .A1(n14307), .A2(n5777), .ZN(n1147) );
  NAND2_X1 U1130 ( .A1(n14307), .A2(n5765), .ZN(n1149) );
  NAND2_X1 U1131 ( .A1(n14307), .A2(n5786), .ZN(n1151) );
  NAND2_X1 U1132 ( .A1(n14307), .A2(n5794), .ZN(n1154) );
  BUF_X1 U1133 ( .A(n14981), .Z(n14975) );
  BUF_X1 U1134 ( .A(n14355), .Z(n14361) );
  BUF_X1 U1135 ( .A(n14981), .Z(n14973) );
  BUF_X1 U1136 ( .A(n14981), .Z(n14974) );
  BUF_X1 U1137 ( .A(n1207), .Z(n14296) );
  BUF_X1 U1138 ( .A(n1180), .Z(n14305) );
  BUF_X1 U1139 ( .A(n1189), .Z(n14302) );
  BUF_X1 U1140 ( .A(n1198), .Z(n14299) );
  BUF_X1 U1141 ( .A(n1220), .Z(n14293) );
  BUF_X1 U1142 ( .A(n1229), .Z(n14290) );
  BUF_X1 U1143 ( .A(n1238), .Z(n14287) );
  BUF_X1 U1144 ( .A(n1247), .Z(n14284) );
  BUF_X1 U1145 ( .A(n5898), .Z(n14447) );
  BUF_X1 U1146 ( .A(n5898), .Z(n14444) );
  BUF_X1 U1147 ( .A(n5898), .Z(n14441) );
  BUF_X1 U1148 ( .A(n5898), .Z(n14438) );
  BUF_X1 U1149 ( .A(n5898), .Z(n14435) );
  BUF_X1 U1150 ( .A(n5898), .Z(n14432) );
  BUF_X1 U1151 ( .A(n5898), .Z(n14429) );
  BUF_X1 U1152 ( .A(n5898), .Z(n14426) );
  BUF_X1 U1153 ( .A(n5898), .Z(n14423) );
  BUF_X1 U1154 ( .A(n5898), .Z(n14420) );
  BUF_X1 U1155 ( .A(n5898), .Z(n14417) );
  BUF_X1 U1156 ( .A(n5898), .Z(n14414) );
  BUF_X1 U1157 ( .A(n5898), .Z(n14411) );
  BUF_X1 U1158 ( .A(n5900), .Z(n14449) );
  BUF_X1 U1159 ( .A(n763), .Z(n14448) );
  BUF_X1 U1160 ( .A(n5900), .Z(n14446) );
  BUF_X1 U1161 ( .A(n763), .Z(n14445) );
  BUF_X1 U1162 ( .A(n5900), .Z(n14443) );
  BUF_X1 U1163 ( .A(n763), .Z(n14442) );
  BUF_X1 U1164 ( .A(n5900), .Z(n14440) );
  BUF_X1 U1165 ( .A(n763), .Z(n14439) );
  BUF_X1 U1166 ( .A(n5900), .Z(n14437) );
  BUF_X1 U1167 ( .A(n763), .Z(n14436) );
  BUF_X1 U1168 ( .A(n5900), .Z(n14434) );
  BUF_X1 U1169 ( .A(n763), .Z(n14433) );
  BUF_X1 U1170 ( .A(n5900), .Z(n14431) );
  BUF_X1 U1171 ( .A(n763), .Z(n14430) );
  BUF_X1 U1172 ( .A(n5900), .Z(n14428) );
  BUF_X1 U1173 ( .A(n763), .Z(n14427) );
  BUF_X1 U1174 ( .A(n5900), .Z(n14425) );
  BUF_X1 U1175 ( .A(n763), .Z(n14424) );
  BUF_X1 U1176 ( .A(n5900), .Z(n14422) );
  BUF_X1 U1177 ( .A(n763), .Z(n14421) );
  BUF_X1 U1178 ( .A(n5900), .Z(n14419) );
  BUF_X1 U1179 ( .A(n763), .Z(n14418) );
  BUF_X1 U1180 ( .A(n5900), .Z(n14416) );
  BUF_X1 U1181 ( .A(n763), .Z(n14415) );
  BUF_X1 U1182 ( .A(n5900), .Z(n14413) );
  BUF_X1 U1183 ( .A(n763), .Z(n14412) );
  BUF_X1 U1184 ( .A(n14355), .Z(n14362) );
  BUF_X1 U1185 ( .A(n14355), .Z(n14363) );
  BUF_X1 U1186 ( .A(n14355), .Z(n14364) );
  BUF_X1 U1187 ( .A(n14355), .Z(n14365) );
  BUF_X1 U1188 ( .A(n14355), .Z(n14366) );
  BUF_X1 U1189 ( .A(n14355), .Z(n14367) );
  BUF_X1 U1190 ( .A(n14356), .Z(n14368) );
  BUF_X1 U1191 ( .A(n14356), .Z(n14369) );
  BUF_X1 U1192 ( .A(n14356), .Z(n14370) );
  BUF_X1 U1193 ( .A(n14356), .Z(n14371) );
  BUF_X1 U1194 ( .A(n14356), .Z(n14372) );
  BUF_X1 U1195 ( .A(n14356), .Z(n14373) );
  BUF_X1 U1196 ( .A(n14356), .Z(n14374) );
  BUF_X1 U1197 ( .A(n14357), .Z(n14375) );
  BUF_X1 U1198 ( .A(n14357), .Z(n14376) );
  BUF_X1 U1199 ( .A(n14357), .Z(n14377) );
  BUF_X1 U1200 ( .A(n14357), .Z(n14378) );
  BUF_X1 U1201 ( .A(n14357), .Z(n14379) );
  BUF_X1 U1202 ( .A(n14357), .Z(n14380) );
  BUF_X1 U1203 ( .A(n14357), .Z(n14381) );
  BUF_X1 U1204 ( .A(n14358), .Z(n14382) );
  BUF_X1 U1205 ( .A(n14358), .Z(n14383) );
  BUF_X1 U1206 ( .A(n14358), .Z(n14384) );
  BUF_X1 U1207 ( .A(n14358), .Z(n14385) );
  BUF_X1 U1208 ( .A(n14358), .Z(n14386) );
  BUF_X1 U1209 ( .A(n14358), .Z(n14387) );
  BUF_X1 U1210 ( .A(n14358), .Z(n14388) );
  BUF_X1 U1211 ( .A(n14359), .Z(n14389) );
  BUF_X1 U1212 ( .A(n14359), .Z(n14390) );
  BUF_X1 U1213 ( .A(n14359), .Z(n14391) );
  BUF_X1 U1214 ( .A(n14359), .Z(n14392) );
  BUF_X1 U1215 ( .A(n14359), .Z(n14393) );
  BUF_X1 U1216 ( .A(n14359), .Z(n14394) );
  BUF_X1 U1217 ( .A(n14359), .Z(n14395) );
  BUF_X1 U1218 ( .A(n14360), .Z(n14396) );
  BUF_X1 U1219 ( .A(n14360), .Z(n14397) );
  BUF_X1 U1220 ( .A(n14360), .Z(n14398) );
  BUF_X1 U1221 ( .A(n14360), .Z(n14399) );
  BUF_X1 U1222 ( .A(n1180), .Z(n14303) );
  BUF_X1 U1223 ( .A(n1189), .Z(n14300) );
  BUF_X1 U1224 ( .A(n1198), .Z(n14297) );
  BUF_X1 U1225 ( .A(n1207), .Z(n14294) );
  BUF_X1 U1226 ( .A(n1220), .Z(n14291) );
  BUF_X1 U1227 ( .A(n1229), .Z(n14288) );
  BUF_X1 U1228 ( .A(n1238), .Z(n14285) );
  BUF_X1 U1229 ( .A(n1247), .Z(n14282) );
  BUF_X1 U1230 ( .A(n1180), .Z(n14304) );
  BUF_X1 U1231 ( .A(n1189), .Z(n14301) );
  BUF_X1 U1232 ( .A(n1198), .Z(n14298) );
  BUF_X1 U1233 ( .A(n1207), .Z(n14295) );
  BUF_X1 U1234 ( .A(n1220), .Z(n14292) );
  BUF_X1 U1235 ( .A(n1229), .Z(n14289) );
  BUF_X1 U1236 ( .A(n1238), .Z(n14286) );
  BUF_X1 U1237 ( .A(n1247), .Z(n14283) );
  BUF_X1 U1238 ( .A(n14976), .Z(n14977) );
  BUF_X1 U1239 ( .A(n14976), .Z(n14978) );
  BUF_X1 U1240 ( .A(n14976), .Z(n14979) );
  BUF_X1 U1241 ( .A(n14976), .Z(n14980) );
  NOR3_X1 U1242 ( .A1(n14974), .A2(n14606), .A3(n14987), .ZN(n242) );
  NOR3_X1 U1243 ( .A1(n14987), .A2(n14974), .A3(n14553), .ZN(n504) );
  NOR3_X1 U1244 ( .A1(n14987), .A2(n14973), .A3(n14509), .ZN(n569) );
  NOR3_X1 U1245 ( .A1(n14987), .A2(n14973), .A3(n14361), .ZN(n1028) );
  BUF_X1 U1246 ( .A(n959), .Z(n14355) );
  AND3_X1 U1247 ( .A1(n14972), .A2(n14987), .A3(n14450), .ZN(n700) );
  AND3_X1 U1248 ( .A1(n14972), .A2(n14987), .A3(n14351), .ZN(n962) );
  AND3_X1 U1249 ( .A1(n14972), .A2(n14987), .A3(n14493), .ZN(n634) );
  AND3_X1 U1250 ( .A1(n14972), .A2(n14987), .A3(n5897), .ZN(n175) );
  BUF_X1 U1251 ( .A(n14646), .Z(n14649) );
  BUF_X1 U1252 ( .A(n307), .Z(n14599) );
  BUF_X1 U1253 ( .A(n766), .Z(n14410) );
  BUF_X1 U1254 ( .A(n831), .Z(n14407) );
  BUF_X1 U1255 ( .A(n1093), .Z(n14308) );
  BUF_X1 U1256 ( .A(n14593), .Z(n14596) );
  BUF_X1 U1257 ( .A(n14552), .Z(n14551) );
  BUF_X1 U1258 ( .A(n14404), .Z(n14403) );
  BUF_X1 U1259 ( .A(n14503), .Z(n14509) );
  BUF_X1 U1260 ( .A(n435), .Z(n14553) );
  INV_X1 U1261 ( .A(WE), .ZN(n14981) );
  BUF_X1 U1262 ( .A(n959), .Z(n14356) );
  BUF_X1 U1263 ( .A(n959), .Z(n14357) );
  BUF_X1 U1264 ( .A(n959), .Z(n14358) );
  BUF_X1 U1265 ( .A(n959), .Z(n14359) );
  BUF_X1 U1266 ( .A(n959), .Z(n14360) );
  BUF_X1 U1267 ( .A(n1260), .Z(n14281) );
  BUF_X1 U1268 ( .A(n1269), .Z(n5956) );
  BUF_X1 U1269 ( .A(n1300), .Z(n5937) );
  BUF_X1 U1270 ( .A(n1309), .Z(n5933) );
  BUF_X1 U1271 ( .A(n1278), .Z(n5950) );
  BUF_X1 U1272 ( .A(n1287), .Z(n5944) );
  BUF_X1 U1273 ( .A(n1318), .Z(n5926) );
  BUF_X1 U1274 ( .A(n1327), .Z(n5916) );
  BUF_X1 U1275 ( .A(n435), .Z(n14591) );
  BUF_X1 U1276 ( .A(n5905), .Z(n14590) );
  BUF_X1 U1277 ( .A(n5908), .Z(n14348) );
  BUF_X1 U1278 ( .A(n5908), .Z(n14345) );
  BUF_X1 U1279 ( .A(n5908), .Z(n14342) );
  BUF_X1 U1280 ( .A(n5908), .Z(n14339) );
  BUF_X1 U1281 ( .A(n5908), .Z(n14336) );
  BUF_X1 U1282 ( .A(n5908), .Z(n14333) );
  BUF_X1 U1283 ( .A(n5908), .Z(n14330) );
  BUF_X1 U1284 ( .A(n5908), .Z(n14327) );
  BUF_X1 U1285 ( .A(n5908), .Z(n14324) );
  BUF_X1 U1286 ( .A(n5908), .Z(n14321) );
  BUF_X1 U1287 ( .A(n5908), .Z(n14318) );
  BUF_X1 U1288 ( .A(n5908), .Z(n14315) );
  BUF_X1 U1289 ( .A(n5908), .Z(n14312) );
  BUF_X1 U1290 ( .A(n5909), .Z(n14350) );
  BUF_X1 U1291 ( .A(n1025), .Z(n14349) );
  BUF_X1 U1292 ( .A(n5909), .Z(n14347) );
  BUF_X1 U1293 ( .A(n1025), .Z(n14346) );
  BUF_X1 U1294 ( .A(n5909), .Z(n14344) );
  BUF_X1 U1295 ( .A(n1025), .Z(n14343) );
  BUF_X1 U1296 ( .A(n5909), .Z(n14341) );
  BUF_X1 U1297 ( .A(n1025), .Z(n14340) );
  BUF_X1 U1298 ( .A(n5909), .Z(n14338) );
  BUF_X1 U1299 ( .A(n1025), .Z(n14337) );
  BUF_X1 U1300 ( .A(n5909), .Z(n14335) );
  BUF_X1 U1301 ( .A(n1025), .Z(n14334) );
  BUF_X1 U1302 ( .A(n5909), .Z(n14332) );
  BUF_X1 U1303 ( .A(n1025), .Z(n14331) );
  BUF_X1 U1304 ( .A(n5909), .Z(n14329) );
  BUF_X1 U1305 ( .A(n1025), .Z(n14328) );
  BUF_X1 U1306 ( .A(n5909), .Z(n14326) );
  BUF_X1 U1307 ( .A(n1025), .Z(n14325) );
  BUF_X1 U1308 ( .A(n5909), .Z(n14323) );
  BUF_X1 U1309 ( .A(n1025), .Z(n14322) );
  BUF_X1 U1310 ( .A(n5909), .Z(n14320) );
  BUF_X1 U1311 ( .A(n1025), .Z(n14319) );
  BUF_X1 U1312 ( .A(n5909), .Z(n14317) );
  BUF_X1 U1313 ( .A(n1025), .Z(n14316) );
  BUF_X1 U1314 ( .A(n5909), .Z(n14314) );
  BUF_X1 U1315 ( .A(n1025), .Z(n14313) );
  BUF_X1 U1316 ( .A(n14503), .Z(n14510) );
  BUF_X1 U1317 ( .A(n14503), .Z(n14511) );
  BUF_X1 U1318 ( .A(n14503), .Z(n14512) );
  BUF_X1 U1319 ( .A(n14503), .Z(n14513) );
  BUF_X1 U1320 ( .A(n14503), .Z(n14514) );
  BUF_X1 U1321 ( .A(n14503), .Z(n14515) );
  BUF_X1 U1322 ( .A(n14504), .Z(n14516) );
  BUF_X1 U1323 ( .A(n14504), .Z(n14517) );
  BUF_X1 U1324 ( .A(n14504), .Z(n14518) );
  BUF_X1 U1325 ( .A(n14504), .Z(n14519) );
  BUF_X1 U1326 ( .A(n14504), .Z(n14520) );
  BUF_X1 U1327 ( .A(n14504), .Z(n14521) );
  BUF_X1 U1328 ( .A(n14504), .Z(n14522) );
  BUF_X1 U1329 ( .A(n14505), .Z(n14523) );
  BUF_X1 U1330 ( .A(n14505), .Z(n14524) );
  BUF_X1 U1331 ( .A(n14505), .Z(n14525) );
  BUF_X1 U1332 ( .A(n14505), .Z(n14526) );
  BUF_X1 U1333 ( .A(n14505), .Z(n14527) );
  BUF_X1 U1334 ( .A(n14505), .Z(n14528) );
  BUF_X1 U1335 ( .A(n14505), .Z(n14529) );
  BUF_X1 U1336 ( .A(n14506), .Z(n14530) );
  BUF_X1 U1337 ( .A(n14506), .Z(n14531) );
  BUF_X1 U1338 ( .A(n14506), .Z(n14532) );
  BUF_X1 U1339 ( .A(n14506), .Z(n14533) );
  BUF_X1 U1340 ( .A(n14506), .Z(n14534) );
  BUF_X1 U1341 ( .A(n14506), .Z(n14535) );
  BUF_X1 U1342 ( .A(n14506), .Z(n14536) );
  BUF_X1 U1343 ( .A(n14507), .Z(n14537) );
  BUF_X1 U1344 ( .A(n14507), .Z(n14538) );
  BUF_X1 U1345 ( .A(n14507), .Z(n14539) );
  BUF_X1 U1346 ( .A(n14507), .Z(n14540) );
  BUF_X1 U1347 ( .A(n14507), .Z(n14541) );
  BUF_X1 U1348 ( .A(n14507), .Z(n14542) );
  BUF_X1 U1349 ( .A(n14507), .Z(n14543) );
  BUF_X1 U1350 ( .A(n14508), .Z(n14544) );
  BUF_X1 U1351 ( .A(n14508), .Z(n14545) );
  BUF_X1 U1352 ( .A(n14508), .Z(n14546) );
  BUF_X1 U1353 ( .A(n14508), .Z(n14547) );
  BUF_X1 U1354 ( .A(n1260), .Z(n5957) );
  BUF_X1 U1355 ( .A(n1269), .Z(n5954) );
  BUF_X1 U1356 ( .A(n1300), .Z(n5934) );
  BUF_X1 U1357 ( .A(n1309), .Z(n5928) );
  BUF_X1 U1358 ( .A(n1260), .Z(n14280) );
  BUF_X1 U1359 ( .A(n1269), .Z(n5955) );
  BUF_X1 U1360 ( .A(n1300), .Z(n5936) );
  BUF_X1 U1361 ( .A(n1309), .Z(n5929) );
  BUF_X1 U1362 ( .A(n1278), .Z(n5945) );
  BUF_X1 U1363 ( .A(n1287), .Z(n5941) );
  BUF_X1 U1364 ( .A(n1318), .Z(n5917) );
  BUF_X1 U1365 ( .A(n1327), .Z(n5913) );
  BUF_X1 U1366 ( .A(n1278), .Z(n5949) );
  BUF_X1 U1367 ( .A(n1287), .Z(n5942) );
  BUF_X1 U1368 ( .A(n1318), .Z(n5925) );
  BUF_X1 U1369 ( .A(n1327), .Z(n5914) );
  BUF_X1 U1370 ( .A(n435), .Z(n14555) );
  BUF_X1 U1371 ( .A(n435), .Z(n14557) );
  BUF_X1 U1372 ( .A(n435), .Z(n14559) );
  BUF_X1 U1373 ( .A(n435), .Z(n14561) );
  BUF_X1 U1374 ( .A(n435), .Z(n14563) );
  BUF_X1 U1375 ( .A(n435), .Z(n14565) );
  BUF_X1 U1376 ( .A(n435), .Z(n14567) );
  BUF_X1 U1377 ( .A(n435), .Z(n14569) );
  BUF_X1 U1378 ( .A(n435), .Z(n14571) );
  BUF_X1 U1379 ( .A(n435), .Z(n14573) );
  BUF_X1 U1380 ( .A(n435), .Z(n14575) );
  BUF_X1 U1381 ( .A(n435), .Z(n14577) );
  BUF_X1 U1382 ( .A(n435), .Z(n14579) );
  BUF_X1 U1383 ( .A(n435), .Z(n14581) );
  BUF_X1 U1384 ( .A(n435), .Z(n14583) );
  BUF_X1 U1385 ( .A(n435), .Z(n14585) );
  BUF_X1 U1386 ( .A(n435), .Z(n14587) );
  BUF_X1 U1387 ( .A(n435), .Z(n14589) );
  BUF_X1 U1388 ( .A(n697), .Z(n14492) );
  BUF_X1 U1389 ( .A(n697), .Z(n14490) );
  BUF_X1 U1390 ( .A(n697), .Z(n14488) );
  BUF_X1 U1391 ( .A(n697), .Z(n14486) );
  BUF_X1 U1392 ( .A(n697), .Z(n14484) );
  BUF_X1 U1393 ( .A(n697), .Z(n14482) );
  BUF_X1 U1394 ( .A(n697), .Z(n14480) );
  BUF_X1 U1395 ( .A(n697), .Z(n14478) );
  BUF_X1 U1396 ( .A(n697), .Z(n14476) );
  BUF_X1 U1397 ( .A(n697), .Z(n14474) );
  BUF_X1 U1398 ( .A(n697), .Z(n14472) );
  BUF_X1 U1399 ( .A(n697), .Z(n14470) );
  BUF_X1 U1400 ( .A(n697), .Z(n14468) );
  BUF_X1 U1401 ( .A(n697), .Z(n14466) );
  BUF_X1 U1402 ( .A(n697), .Z(n14464) );
  BUF_X1 U1403 ( .A(n697), .Z(n14462) );
  BUF_X1 U1404 ( .A(n697), .Z(n14460) );
  BUF_X1 U1405 ( .A(n697), .Z(n14458) );
  BUF_X1 U1406 ( .A(n697), .Z(n14456) );
  BUF_X1 U1407 ( .A(n697), .Z(n14454) );
  BUF_X1 U1408 ( .A(n5905), .Z(n14554) );
  BUF_X1 U1409 ( .A(n5905), .Z(n14556) );
  BUF_X1 U1410 ( .A(n5905), .Z(n14558) );
  BUF_X1 U1411 ( .A(n5905), .Z(n14560) );
  BUF_X1 U1412 ( .A(n5905), .Z(n14562) );
  BUF_X1 U1413 ( .A(n5905), .Z(n14564) );
  BUF_X1 U1414 ( .A(n5905), .Z(n14566) );
  BUF_X1 U1415 ( .A(n5905), .Z(n14568) );
  BUF_X1 U1416 ( .A(n5905), .Z(n14570) );
  BUF_X1 U1417 ( .A(n5905), .Z(n14572) );
  BUF_X1 U1418 ( .A(n5905), .Z(n14574) );
  BUF_X1 U1419 ( .A(n5905), .Z(n14576) );
  BUF_X1 U1420 ( .A(n5905), .Z(n14578) );
  BUF_X1 U1421 ( .A(n5905), .Z(n14580) );
  BUF_X1 U1422 ( .A(n5905), .Z(n14582) );
  BUF_X1 U1423 ( .A(n5905), .Z(n14584) );
  BUF_X1 U1424 ( .A(n5905), .Z(n14586) );
  BUF_X1 U1425 ( .A(n5905), .Z(n14588) );
  BUF_X1 U1426 ( .A(n5901), .Z(n14491) );
  BUF_X1 U1427 ( .A(n5901), .Z(n14489) );
  BUF_X1 U1428 ( .A(n5901), .Z(n14487) );
  BUF_X1 U1429 ( .A(n5901), .Z(n14485) );
  BUF_X1 U1430 ( .A(n5901), .Z(n14483) );
  BUF_X1 U1431 ( .A(n5901), .Z(n14481) );
  BUF_X1 U1432 ( .A(n5901), .Z(n14479) );
  BUF_X1 U1433 ( .A(n5901), .Z(n14477) );
  BUF_X1 U1434 ( .A(n5901), .Z(n14475) );
  BUF_X1 U1435 ( .A(n5901), .Z(n14473) );
  BUF_X1 U1436 ( .A(n5901), .Z(n14471) );
  BUF_X1 U1437 ( .A(n5901), .Z(n14469) );
  BUF_X1 U1438 ( .A(n5901), .Z(n14467) );
  BUF_X1 U1439 ( .A(n5901), .Z(n14465) );
  BUF_X1 U1440 ( .A(n5901), .Z(n14463) );
  BUF_X1 U1441 ( .A(n5901), .Z(n14461) );
  BUF_X1 U1442 ( .A(n5901), .Z(n14459) );
  BUF_X1 U1443 ( .A(n5901), .Z(n14457) );
  BUF_X1 U1444 ( .A(n5901), .Z(n14455) );
  OR2_X1 U1445 ( .A1(n1169), .A2(n14972), .ZN(n14184) );
  OR2_X1 U1446 ( .A1(n1334), .A2(n14972), .ZN(n14187) );
  OR2_X1 U1447 ( .A1(n1483), .A2(n14972), .ZN(n14190) );
  OR2_X1 U1448 ( .A1(n1632), .A2(n14972), .ZN(n14193) );
  OR2_X1 U1449 ( .A1(n1781), .A2(n14972), .ZN(n14196) );
  OR2_X1 U1450 ( .A1(n1930), .A2(n14972), .ZN(n14199) );
  OR2_X1 U1451 ( .A1(n2079), .A2(n14972), .ZN(n14202) );
  OR2_X1 U1452 ( .A1(n2228), .A2(n14972), .ZN(n14205) );
  OR2_X1 U1453 ( .A1(n2377), .A2(n14972), .ZN(n14208) );
  OR2_X1 U1454 ( .A1(n2526), .A2(n14972), .ZN(n14211) );
  OR2_X1 U1455 ( .A1(n2675), .A2(n14972), .ZN(n14214) );
  OR2_X1 U1456 ( .A1(n2824), .A2(n14972), .ZN(n14217) );
  OR2_X1 U1457 ( .A1(n2973), .A2(n14972), .ZN(n14220) );
  OR2_X1 U1458 ( .A1(n3122), .A2(n14972), .ZN(n14223) );
  OR2_X1 U1459 ( .A1(n3271), .A2(n14972), .ZN(n14226) );
  OR2_X1 U1460 ( .A1(n3420), .A2(n14972), .ZN(n14229) );
  OR2_X1 U1461 ( .A1(n3569), .A2(n14972), .ZN(n14232) );
  OR2_X1 U1462 ( .A1(n3718), .A2(n14972), .ZN(n14235) );
  OR2_X1 U1463 ( .A1(n3867), .A2(n14972), .ZN(n14238) );
  OR2_X1 U1464 ( .A1(n4016), .A2(n14971), .ZN(n14241) );
  OR2_X1 U1465 ( .A1(n4165), .A2(n14970), .ZN(n14244) );
  OR2_X1 U1466 ( .A1(n4314), .A2(n14970), .ZN(n14247) );
  OR2_X1 U1467 ( .A1(n4463), .A2(n14971), .ZN(n14250) );
  OR2_X1 U1468 ( .A1(n4612), .A2(n14970), .ZN(n14253) );
  OR2_X1 U1469 ( .A1(n4761), .A2(n14971), .ZN(n14256) );
  OR2_X1 U1470 ( .A1(n4910), .A2(n14970), .ZN(n14259) );
  OR2_X1 U1471 ( .A1(n5059), .A2(n14971), .ZN(n14262) );
  OR2_X1 U1472 ( .A1(n5208), .A2(n14970), .ZN(n14265) );
  OR2_X1 U1473 ( .A1(n5357), .A2(n14971), .ZN(n14268) );
  OR2_X1 U1474 ( .A1(n5506), .A2(n14972), .ZN(n14271) );
  OR2_X1 U1475 ( .A1(n5655), .A2(n14970), .ZN(n14274) );
  OR2_X1 U1476 ( .A1(n5804), .A2(n14971), .ZN(n14277) );
  BUF_X1 U1477 ( .A(n501), .Z(n14503) );
  AND2_X1 U1478 ( .A1(OFFSET[1]), .A2(n1164), .ZN(n1101) );
  AND2_X1 U1479 ( .A1(OFFSET[1]), .A2(OFFSET[0]), .ZN(n1104) );
  AND3_X1 U1480 ( .A1(n5897), .A2(n14972), .A3(n14984), .ZN(n307) );
  AND3_X1 U1481 ( .A1(n14984), .A2(n14972), .A3(n14450), .ZN(n831) );
  AND3_X1 U1482 ( .A1(n14985), .A2(n14972), .A3(n14351), .ZN(n1093) );
  AND3_X1 U1483 ( .A1(n14984), .A2(n14972), .A3(n14493), .ZN(n766) );
  AND3_X1 U1484 ( .A1(n5887), .A2(n5888), .A3(OFFSET[4]), .ZN(n1134) );
  AND3_X1 U1485 ( .A1(OFFSET[2]), .A2(n5888), .A3(OFFSET[4]), .ZN(n1143) );
  AND3_X1 U1486 ( .A1(OFFSET[3]), .A2(n5887), .A3(OFFSET[4]), .ZN(n1152) );
  AND3_X1 U1487 ( .A1(OFFSET[3]), .A2(OFFSET[2]), .A3(OFFSET[4]), .ZN(n1161)
         );
  AND2_X1 U1488 ( .A1(n5952), .A2(n14988), .ZN(n239) );
  NOR2_X1 U1489 ( .A1(n14982), .A2(ADDR[3]), .ZN(n5952) );
  BUF_X1 U1490 ( .A(n896), .Z(n14404) );
  NOR3_X1 U1491 ( .A1(n14975), .A2(n14984), .A3(n14361), .ZN(n896) );
  BUF_X1 U1492 ( .A(n372), .Z(n14593) );
  NOR3_X1 U1493 ( .A1(n14975), .A2(n14983), .A3(n14553), .ZN(n372) );
  BUF_X1 U1494 ( .A(n77), .Z(n14646) );
  NOR3_X1 U1495 ( .A1(n14606), .A2(n14983), .A3(n14973), .ZN(n77) );
  BUF_X1 U1496 ( .A(n438), .Z(n14552) );
  NOR3_X1 U1497 ( .A1(n14974), .A2(n14983), .A3(n14509), .ZN(n438) );
  AND2_X1 U1498 ( .A1(ADDR[3]), .A2(n14988), .ZN(n5959) );
  INV_X1 U1499 ( .A(OFFSET[3]), .ZN(n5888) );
  INV_X1 U1500 ( .A(OFFSET[2]), .ZN(n5887) );
  BUF_X1 U1501 ( .A(n171), .Z(n14606) );
  INV_X1 U1502 ( .A(n14984), .ZN(n14987) );
  INV_X1 U1503 ( .A(OFFSET[0]), .ZN(n1164) );
  BUF_X1 U1504 ( .A(n68), .Z(n14930) );
  BUF_X1 U1505 ( .A(n69), .Z(n14890) );
  BUF_X1 U1506 ( .A(n70), .Z(n14850) );
  BUF_X1 U1507 ( .A(n71), .Z(n14810) );
  BUF_X1 U1508 ( .A(n72), .Z(n14770) );
  BUF_X1 U1509 ( .A(n73), .Z(n14730) );
  BUF_X1 U1510 ( .A(n74), .Z(n14690) );
  BUF_X1 U1511 ( .A(n75), .Z(n14650) );
  BUF_X1 U1512 ( .A(n68), .Z(n14958) );
  BUF_X1 U1513 ( .A(n69), .Z(n14891) );
  BUF_X1 U1514 ( .A(n70), .Z(n14851) );
  BUF_X1 U1515 ( .A(n71), .Z(n14811) );
  BUF_X1 U1516 ( .A(n72), .Z(n14771) );
  BUF_X1 U1517 ( .A(n73), .Z(n14731) );
  BUF_X1 U1518 ( .A(n74), .Z(n14691) );
  BUF_X1 U1519 ( .A(n75), .Z(n14651) );
  BUF_X1 U1520 ( .A(n68), .Z(n14957) );
  BUF_X1 U1521 ( .A(n69), .Z(n14892) );
  BUF_X1 U1522 ( .A(n70), .Z(n14852) );
  BUF_X1 U1523 ( .A(n71), .Z(n14812) );
  BUF_X1 U1524 ( .A(n72), .Z(n14772) );
  BUF_X1 U1525 ( .A(n73), .Z(n14732) );
  BUF_X1 U1526 ( .A(n74), .Z(n14692) );
  BUF_X1 U1527 ( .A(n75), .Z(n14652) );
  BUF_X1 U1528 ( .A(n68), .Z(n14956) );
  BUF_X1 U1529 ( .A(n69), .Z(n14893) );
  BUF_X1 U1530 ( .A(n70), .Z(n14853) );
  BUF_X1 U1531 ( .A(n71), .Z(n14813) );
  BUF_X1 U1532 ( .A(n72), .Z(n14773) );
  BUF_X1 U1533 ( .A(n73), .Z(n14733) );
  BUF_X1 U1534 ( .A(n74), .Z(n14693) );
  BUF_X1 U1535 ( .A(n75), .Z(n14653) );
  BUF_X1 U1536 ( .A(n68), .Z(n14955) );
  BUF_X1 U1537 ( .A(n69), .Z(n14894) );
  BUF_X1 U1538 ( .A(n70), .Z(n14854) );
  BUF_X1 U1539 ( .A(n71), .Z(n14814) );
  BUF_X1 U1540 ( .A(n72), .Z(n14774) );
  BUF_X1 U1541 ( .A(n73), .Z(n14734) );
  BUF_X1 U1542 ( .A(n74), .Z(n14694) );
  BUF_X1 U1543 ( .A(n75), .Z(n14654) );
  BUF_X1 U1544 ( .A(n69), .Z(n14895) );
  BUF_X1 U1545 ( .A(n70), .Z(n14855) );
  BUF_X1 U1546 ( .A(n71), .Z(n14815) );
  BUF_X1 U1547 ( .A(n72), .Z(n14775) );
  BUF_X1 U1548 ( .A(n73), .Z(n14735) );
  BUF_X1 U1549 ( .A(n74), .Z(n14695) );
  BUF_X1 U1550 ( .A(n75), .Z(n14655) );
  BUF_X1 U1551 ( .A(n68), .Z(n14953) );
  BUF_X1 U1552 ( .A(n69), .Z(n14896) );
  BUF_X1 U1553 ( .A(n70), .Z(n14856) );
  BUF_X1 U1554 ( .A(n71), .Z(n14816) );
  BUF_X1 U1555 ( .A(n72), .Z(n14776) );
  BUF_X1 U1556 ( .A(n73), .Z(n14736) );
  BUF_X1 U1557 ( .A(n74), .Z(n14696) );
  BUF_X1 U1558 ( .A(n75), .Z(n14656) );
  BUF_X1 U1559 ( .A(n68), .Z(n14952) );
  BUF_X1 U1560 ( .A(n69), .Z(n14897) );
  BUF_X1 U1561 ( .A(n70), .Z(n14857) );
  BUF_X1 U1562 ( .A(n71), .Z(n14817) );
  BUF_X1 U1563 ( .A(n72), .Z(n14777) );
  BUF_X1 U1564 ( .A(n73), .Z(n14737) );
  BUF_X1 U1565 ( .A(n74), .Z(n14697) );
  BUF_X1 U1566 ( .A(n75), .Z(n14657) );
  BUF_X1 U1567 ( .A(n68), .Z(n14951) );
  BUF_X1 U1568 ( .A(n69), .Z(n14898) );
  BUF_X1 U1569 ( .A(n70), .Z(n14858) );
  BUF_X1 U1570 ( .A(n71), .Z(n14818) );
  BUF_X1 U1571 ( .A(n72), .Z(n14778) );
  BUF_X1 U1572 ( .A(n73), .Z(n14738) );
  BUF_X1 U1573 ( .A(n74), .Z(n14698) );
  BUF_X1 U1574 ( .A(n75), .Z(n14658) );
  BUF_X1 U1575 ( .A(n68), .Z(n14950) );
  BUF_X1 U1576 ( .A(n68), .Z(n14954) );
  BUF_X1 U1577 ( .A(n69), .Z(n14899) );
  BUF_X1 U1578 ( .A(n70), .Z(n14859) );
  BUF_X1 U1579 ( .A(n71), .Z(n14819) );
  BUF_X1 U1580 ( .A(n72), .Z(n14779) );
  BUF_X1 U1581 ( .A(n73), .Z(n14739) );
  BUF_X1 U1582 ( .A(n74), .Z(n14699) );
  BUF_X1 U1583 ( .A(n75), .Z(n14659) );
  BUF_X1 U1584 ( .A(n69), .Z(n14900) );
  BUF_X1 U1585 ( .A(n70), .Z(n14860) );
  BUF_X1 U1586 ( .A(n71), .Z(n14820) );
  BUF_X1 U1587 ( .A(n72), .Z(n14780) );
  BUF_X1 U1588 ( .A(n73), .Z(n14740) );
  BUF_X1 U1589 ( .A(n74), .Z(n14700) );
  BUF_X1 U1590 ( .A(n75), .Z(n14660) );
  BUF_X1 U1591 ( .A(n69), .Z(n14901) );
  BUF_X1 U1592 ( .A(n70), .Z(n14861) );
  BUF_X1 U1593 ( .A(n71), .Z(n14821) );
  BUF_X1 U1594 ( .A(n72), .Z(n14781) );
  BUF_X1 U1595 ( .A(n73), .Z(n14741) );
  BUF_X1 U1596 ( .A(n74), .Z(n14701) );
  BUF_X1 U1597 ( .A(n75), .Z(n14661) );
  BUF_X1 U1598 ( .A(n68), .Z(n14967) );
  BUF_X1 U1599 ( .A(n69), .Z(n14902) );
  BUF_X1 U1600 ( .A(n70), .Z(n14862) );
  BUF_X1 U1601 ( .A(n71), .Z(n14822) );
  BUF_X1 U1602 ( .A(n72), .Z(n14782) );
  BUF_X1 U1603 ( .A(n73), .Z(n14742) );
  BUF_X1 U1604 ( .A(n74), .Z(n14702) );
  BUF_X1 U1605 ( .A(n75), .Z(n14662) );
  BUF_X1 U1606 ( .A(n68), .Z(n14966) );
  BUF_X1 U1607 ( .A(n69), .Z(n14903) );
  BUF_X1 U1608 ( .A(n70), .Z(n14863) );
  BUF_X1 U1609 ( .A(n71), .Z(n14823) );
  BUF_X1 U1610 ( .A(n72), .Z(n14783) );
  BUF_X1 U1611 ( .A(n73), .Z(n14743) );
  BUF_X1 U1612 ( .A(n74), .Z(n14703) );
  BUF_X1 U1613 ( .A(n75), .Z(n14663) );
  BUF_X1 U1614 ( .A(n68), .Z(n14965) );
  BUF_X1 U1615 ( .A(n69), .Z(n14904) );
  BUF_X1 U1616 ( .A(n70), .Z(n14864) );
  BUF_X1 U1617 ( .A(n71), .Z(n14824) );
  BUF_X1 U1618 ( .A(n72), .Z(n14784) );
  BUF_X1 U1619 ( .A(n73), .Z(n14744) );
  BUF_X1 U1620 ( .A(n74), .Z(n14704) );
  BUF_X1 U1621 ( .A(n75), .Z(n14664) );
  BUF_X1 U1622 ( .A(n69), .Z(n14905) );
  BUF_X1 U1623 ( .A(n70), .Z(n14865) );
  BUF_X1 U1624 ( .A(n71), .Z(n14825) );
  BUF_X1 U1625 ( .A(n72), .Z(n14785) );
  BUF_X1 U1626 ( .A(n73), .Z(n14745) );
  BUF_X1 U1627 ( .A(n74), .Z(n14705) );
  BUF_X1 U1628 ( .A(n75), .Z(n14665) );
  BUF_X1 U1629 ( .A(n68), .Z(n14963) );
  BUF_X1 U1630 ( .A(n69), .Z(n14906) );
  BUF_X1 U1631 ( .A(n70), .Z(n14866) );
  BUF_X1 U1632 ( .A(n71), .Z(n14826) );
  BUF_X1 U1633 ( .A(n72), .Z(n14786) );
  BUF_X1 U1634 ( .A(n73), .Z(n14746) );
  BUF_X1 U1635 ( .A(n74), .Z(n14706) );
  BUF_X1 U1636 ( .A(n75), .Z(n14666) );
  BUF_X1 U1637 ( .A(n68), .Z(n14962) );
  BUF_X1 U1638 ( .A(n69), .Z(n14907) );
  BUF_X1 U1639 ( .A(n70), .Z(n14867) );
  BUF_X1 U1640 ( .A(n71), .Z(n14827) );
  BUF_X1 U1641 ( .A(n72), .Z(n14787) );
  BUF_X1 U1642 ( .A(n73), .Z(n14747) );
  BUF_X1 U1643 ( .A(n74), .Z(n14707) );
  BUF_X1 U1644 ( .A(n75), .Z(n14667) );
  BUF_X1 U1645 ( .A(n68), .Z(n14961) );
  BUF_X1 U1646 ( .A(n69), .Z(n14908) );
  BUF_X1 U1647 ( .A(n70), .Z(n14868) );
  BUF_X1 U1648 ( .A(n71), .Z(n14828) );
  BUF_X1 U1649 ( .A(n72), .Z(n14788) );
  BUF_X1 U1650 ( .A(n73), .Z(n14748) );
  BUF_X1 U1651 ( .A(n74), .Z(n14708) );
  BUF_X1 U1652 ( .A(n75), .Z(n14668) );
  BUF_X1 U1653 ( .A(n68), .Z(n14960) );
  BUF_X1 U1654 ( .A(n68), .Z(n14959) );
  BUF_X1 U1655 ( .A(n68), .Z(n14964) );
  BUF_X1 U1656 ( .A(n69), .Z(n14909) );
  BUF_X1 U1657 ( .A(n70), .Z(n14869) );
  BUF_X1 U1658 ( .A(n71), .Z(n14829) );
  BUF_X1 U1659 ( .A(n72), .Z(n14789) );
  BUF_X1 U1660 ( .A(n73), .Z(n14749) );
  BUF_X1 U1661 ( .A(n74), .Z(n14709) );
  BUF_X1 U1662 ( .A(n75), .Z(n14669) );
  BUF_X1 U1663 ( .A(n69), .Z(n14910) );
  BUF_X1 U1664 ( .A(n70), .Z(n14870) );
  BUF_X1 U1665 ( .A(n71), .Z(n14830) );
  BUF_X1 U1666 ( .A(n72), .Z(n14790) );
  BUF_X1 U1667 ( .A(n73), .Z(n14750) );
  BUF_X1 U1668 ( .A(n74), .Z(n14710) );
  BUF_X1 U1669 ( .A(n75), .Z(n14670) );
  BUF_X1 U1670 ( .A(n68), .Z(n14938) );
  BUF_X1 U1671 ( .A(n69), .Z(n14911) );
  BUF_X1 U1672 ( .A(n70), .Z(n14871) );
  BUF_X1 U1673 ( .A(n71), .Z(n14831) );
  BUF_X1 U1674 ( .A(n72), .Z(n14791) );
  BUF_X1 U1675 ( .A(n73), .Z(n14751) );
  BUF_X1 U1676 ( .A(n74), .Z(n14711) );
  BUF_X1 U1677 ( .A(n75), .Z(n14671) );
  BUF_X1 U1678 ( .A(n68), .Z(n14937) );
  BUF_X1 U1679 ( .A(n69), .Z(n14912) );
  BUF_X1 U1680 ( .A(n70), .Z(n14872) );
  BUF_X1 U1681 ( .A(n71), .Z(n14832) );
  BUF_X1 U1682 ( .A(n72), .Z(n14792) );
  BUF_X1 U1683 ( .A(n73), .Z(n14752) );
  BUF_X1 U1684 ( .A(n74), .Z(n14712) );
  BUF_X1 U1685 ( .A(n75), .Z(n14672) );
  BUF_X1 U1686 ( .A(n68), .Z(n14936) );
  BUF_X1 U1687 ( .A(n69), .Z(n14913) );
  BUF_X1 U1688 ( .A(n70), .Z(n14873) );
  BUF_X1 U1689 ( .A(n71), .Z(n14833) );
  BUF_X1 U1690 ( .A(n72), .Z(n14793) );
  BUF_X1 U1691 ( .A(n73), .Z(n14753) );
  BUF_X1 U1692 ( .A(n74), .Z(n14713) );
  BUF_X1 U1693 ( .A(n75), .Z(n14673) );
  BUF_X1 U1694 ( .A(n68), .Z(n14935) );
  BUF_X1 U1695 ( .A(n69), .Z(n14914) );
  BUF_X1 U1696 ( .A(n70), .Z(n14874) );
  BUF_X1 U1697 ( .A(n71), .Z(n14834) );
  BUF_X1 U1698 ( .A(n72), .Z(n14794) );
  BUF_X1 U1699 ( .A(n73), .Z(n14754) );
  BUF_X1 U1700 ( .A(n74), .Z(n14714) );
  BUF_X1 U1701 ( .A(n75), .Z(n14674) );
  BUF_X1 U1702 ( .A(n69), .Z(n14915) );
  BUF_X1 U1703 ( .A(n70), .Z(n14875) );
  BUF_X1 U1704 ( .A(n71), .Z(n14835) );
  BUF_X1 U1705 ( .A(n72), .Z(n14795) );
  BUF_X1 U1706 ( .A(n73), .Z(n14755) );
  BUF_X1 U1707 ( .A(n74), .Z(n14715) );
  BUF_X1 U1708 ( .A(n75), .Z(n14675) );
  BUF_X1 U1709 ( .A(n68), .Z(n14933) );
  BUF_X1 U1710 ( .A(n69), .Z(n14916) );
  BUF_X1 U1711 ( .A(n70), .Z(n14876) );
  BUF_X1 U1712 ( .A(n71), .Z(n14836) );
  BUF_X1 U1713 ( .A(n72), .Z(n14796) );
  BUF_X1 U1714 ( .A(n73), .Z(n14756) );
  BUF_X1 U1715 ( .A(n74), .Z(n14716) );
  BUF_X1 U1716 ( .A(n75), .Z(n14676) );
  BUF_X1 U1717 ( .A(n68), .Z(n14932) );
  BUF_X1 U1718 ( .A(n69), .Z(n14917) );
  BUF_X1 U1719 ( .A(n70), .Z(n14877) );
  BUF_X1 U1720 ( .A(n71), .Z(n14837) );
  BUF_X1 U1721 ( .A(n72), .Z(n14797) );
  BUF_X1 U1722 ( .A(n73), .Z(n14757) );
  BUF_X1 U1723 ( .A(n74), .Z(n14717) );
  BUF_X1 U1724 ( .A(n75), .Z(n14677) );
  BUF_X1 U1725 ( .A(n68), .Z(n14931) );
  BUF_X1 U1726 ( .A(n69), .Z(n14918) );
  BUF_X1 U1727 ( .A(n70), .Z(n14878) );
  BUF_X1 U1728 ( .A(n71), .Z(n14838) );
  BUF_X1 U1729 ( .A(n72), .Z(n14798) );
  BUF_X1 U1730 ( .A(n73), .Z(n14758) );
  BUF_X1 U1731 ( .A(n74), .Z(n14718) );
  BUF_X1 U1732 ( .A(n75), .Z(n14678) );
  BUF_X1 U1733 ( .A(n68), .Z(n14934) );
  BUF_X1 U1734 ( .A(n69), .Z(n14919) );
  BUF_X1 U1735 ( .A(n70), .Z(n14879) );
  BUF_X1 U1736 ( .A(n71), .Z(n14839) );
  BUF_X1 U1737 ( .A(n72), .Z(n14799) );
  BUF_X1 U1738 ( .A(n73), .Z(n14759) );
  BUF_X1 U1739 ( .A(n74), .Z(n14719) );
  BUF_X1 U1740 ( .A(n75), .Z(n14679) );
  BUF_X1 U1741 ( .A(n69), .Z(n14920) );
  BUF_X1 U1742 ( .A(n70), .Z(n14880) );
  BUF_X1 U1743 ( .A(n71), .Z(n14840) );
  BUF_X1 U1744 ( .A(n72), .Z(n14800) );
  BUF_X1 U1745 ( .A(n73), .Z(n14760) );
  BUF_X1 U1746 ( .A(n74), .Z(n14720) );
  BUF_X1 U1747 ( .A(n75), .Z(n14680) );
  BUF_X1 U1748 ( .A(n68), .Z(n14948) );
  BUF_X1 U1749 ( .A(n69), .Z(n14921) );
  BUF_X1 U1750 ( .A(n70), .Z(n14881) );
  BUF_X1 U1751 ( .A(n71), .Z(n14841) );
  BUF_X1 U1752 ( .A(n72), .Z(n14801) );
  BUF_X1 U1753 ( .A(n73), .Z(n14761) );
  BUF_X1 U1754 ( .A(n74), .Z(n14721) );
  BUF_X1 U1755 ( .A(n75), .Z(n14681) );
  BUF_X1 U1756 ( .A(n68), .Z(n14947) );
  BUF_X1 U1757 ( .A(n69), .Z(n14922) );
  BUF_X1 U1758 ( .A(n70), .Z(n14882) );
  BUF_X1 U1759 ( .A(n71), .Z(n14842) );
  BUF_X1 U1760 ( .A(n72), .Z(n14802) );
  BUF_X1 U1761 ( .A(n73), .Z(n14762) );
  BUF_X1 U1762 ( .A(n74), .Z(n14722) );
  BUF_X1 U1763 ( .A(n75), .Z(n14682) );
  BUF_X1 U1764 ( .A(n68), .Z(n14946) );
  BUF_X1 U1765 ( .A(n69), .Z(n14923) );
  BUF_X1 U1766 ( .A(n70), .Z(n14883) );
  BUF_X1 U1767 ( .A(n71), .Z(n14843) );
  BUF_X1 U1768 ( .A(n72), .Z(n14803) );
  BUF_X1 U1769 ( .A(n73), .Z(n14763) );
  BUF_X1 U1770 ( .A(n74), .Z(n14723) );
  BUF_X1 U1771 ( .A(n75), .Z(n14683) );
  BUF_X1 U1772 ( .A(n68), .Z(n14945) );
  BUF_X1 U1773 ( .A(n69), .Z(n14924) );
  BUF_X1 U1774 ( .A(n70), .Z(n14884) );
  BUF_X1 U1775 ( .A(n71), .Z(n14844) );
  BUF_X1 U1776 ( .A(n72), .Z(n14804) );
  BUF_X1 U1777 ( .A(n73), .Z(n14764) );
  BUF_X1 U1778 ( .A(n74), .Z(n14724) );
  BUF_X1 U1779 ( .A(n75), .Z(n14684) );
  BUF_X1 U1780 ( .A(n69), .Z(n14925) );
  BUF_X1 U1781 ( .A(n70), .Z(n14885) );
  BUF_X1 U1782 ( .A(n71), .Z(n14845) );
  BUF_X1 U1783 ( .A(n72), .Z(n14805) );
  BUF_X1 U1784 ( .A(n73), .Z(n14765) );
  BUF_X1 U1785 ( .A(n74), .Z(n14725) );
  BUF_X1 U1786 ( .A(n75), .Z(n14685) );
  BUF_X1 U1787 ( .A(n68), .Z(n14943) );
  BUF_X1 U1788 ( .A(n69), .Z(n14926) );
  BUF_X1 U1789 ( .A(n70), .Z(n14886) );
  BUF_X1 U1790 ( .A(n71), .Z(n14846) );
  BUF_X1 U1791 ( .A(n72), .Z(n14806) );
  BUF_X1 U1792 ( .A(n73), .Z(n14766) );
  BUF_X1 U1793 ( .A(n74), .Z(n14726) );
  BUF_X1 U1794 ( .A(n75), .Z(n14686) );
  BUF_X1 U1795 ( .A(n68), .Z(n14942) );
  BUF_X1 U1796 ( .A(n69), .Z(n14927) );
  BUF_X1 U1797 ( .A(n70), .Z(n14887) );
  BUF_X1 U1798 ( .A(n71), .Z(n14847) );
  BUF_X1 U1799 ( .A(n72), .Z(n14807) );
  BUF_X1 U1800 ( .A(n73), .Z(n14767) );
  BUF_X1 U1801 ( .A(n74), .Z(n14727) );
  BUF_X1 U1802 ( .A(n75), .Z(n14687) );
  BUF_X1 U1803 ( .A(n68), .Z(n14941) );
  BUF_X1 U1804 ( .A(n69), .Z(n14928) );
  BUF_X1 U1805 ( .A(n70), .Z(n14888) );
  BUF_X1 U1806 ( .A(n71), .Z(n14848) );
  BUF_X1 U1807 ( .A(n72), .Z(n14808) );
  BUF_X1 U1808 ( .A(n73), .Z(n14768) );
  BUF_X1 U1809 ( .A(n74), .Z(n14728) );
  BUF_X1 U1810 ( .A(n75), .Z(n14688) );
  BUF_X1 U1811 ( .A(n68), .Z(n14940) );
  BUF_X1 U1812 ( .A(n68), .Z(n14939) );
  BUF_X1 U1813 ( .A(n68), .Z(n14944) );
  BUF_X1 U1814 ( .A(n68), .Z(n14949) );
  BUF_X1 U1815 ( .A(n68), .Z(n14968) );
  NOR4_X1 U1816 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1173)
         );
  AOI21_X1 U1817 ( .B1(n1205), .B2(n1206), .A(n14294), .ZN(n1174) );
  AOI21_X1 U1818 ( .B1(n1196), .B2(n1197), .A(n14297), .ZN(n1175) );
  AOI21_X1 U1819 ( .B1(n1187), .B2(n1188), .A(n14300), .ZN(n1176) );
  NOR4_X1 U1820 ( .A1(n1339), .A2(n1340), .A3(n1341), .A4(n1342), .ZN(n1338)
         );
  AOI21_X1 U1821 ( .B1(n1367), .B2(n1368), .A(n14294), .ZN(n1339) );
  AOI21_X1 U1822 ( .B1(n1359), .B2(n1360), .A(n14297), .ZN(n1340) );
  AOI21_X1 U1823 ( .B1(n1351), .B2(n1352), .A(n14300), .ZN(n1341) );
  NOR4_X1 U1824 ( .A1(n1488), .A2(n1489), .A3(n1490), .A4(n1491), .ZN(n1487)
         );
  AOI21_X1 U1825 ( .B1(n1516), .B2(n1517), .A(n14294), .ZN(n1488) );
  AOI21_X1 U1826 ( .B1(n1508), .B2(n1509), .A(n14297), .ZN(n1489) );
  AOI21_X1 U1827 ( .B1(n1500), .B2(n1501), .A(n14300), .ZN(n1490) );
  NOR4_X1 U1828 ( .A1(n1637), .A2(n1638), .A3(n1639), .A4(n1640), .ZN(n1636)
         );
  AOI21_X1 U1829 ( .B1(n1665), .B2(n1666), .A(n14294), .ZN(n1637) );
  AOI21_X1 U1830 ( .B1(n1657), .B2(n1658), .A(n14297), .ZN(n1638) );
  AOI21_X1 U1831 ( .B1(n1649), .B2(n1650), .A(n14300), .ZN(n1639) );
  NOR4_X1 U1832 ( .A1(n1786), .A2(n1787), .A3(n1788), .A4(n1789), .ZN(n1785)
         );
  AOI21_X1 U1833 ( .B1(n1814), .B2(n1815), .A(n14294), .ZN(n1786) );
  AOI21_X1 U1834 ( .B1(n1806), .B2(n1807), .A(n14297), .ZN(n1787) );
  AOI21_X1 U1835 ( .B1(n1798), .B2(n1799), .A(n14300), .ZN(n1788) );
  NOR4_X1 U1836 ( .A1(n1935), .A2(n1936), .A3(n1937), .A4(n1938), .ZN(n1934)
         );
  AOI21_X1 U1837 ( .B1(n1963), .B2(n1964), .A(n14294), .ZN(n1935) );
  AOI21_X1 U1838 ( .B1(n1955), .B2(n1956), .A(n14297), .ZN(n1936) );
  AOI21_X1 U1839 ( .B1(n1947), .B2(n1948), .A(n14300), .ZN(n1937) );
  NOR4_X1 U1840 ( .A1(n2084), .A2(n2085), .A3(n2086), .A4(n2087), .ZN(n2083)
         );
  AOI21_X1 U1841 ( .B1(n2112), .B2(n2113), .A(n14294), .ZN(n2084) );
  AOI21_X1 U1842 ( .B1(n2104), .B2(n2105), .A(n14297), .ZN(n2085) );
  AOI21_X1 U1843 ( .B1(n2096), .B2(n2097), .A(n14300), .ZN(n2086) );
  NOR4_X1 U1844 ( .A1(n2233), .A2(n2234), .A3(n2235), .A4(n2236), .ZN(n2232)
         );
  AOI21_X1 U1845 ( .B1(n2261), .B2(n2262), .A(n14294), .ZN(n2233) );
  AOI21_X1 U1846 ( .B1(n2253), .B2(n2254), .A(n14297), .ZN(n2234) );
  AOI21_X1 U1847 ( .B1(n2245), .B2(n2246), .A(n14300), .ZN(n2235) );
  NOR4_X1 U1848 ( .A1(n2382), .A2(n2383), .A3(n2384), .A4(n2385), .ZN(n2381)
         );
  AOI21_X1 U1849 ( .B1(n2410), .B2(n2411), .A(n14294), .ZN(n2382) );
  AOI21_X1 U1850 ( .B1(n2402), .B2(n2403), .A(n14297), .ZN(n2383) );
  AOI21_X1 U1851 ( .B1(n2394), .B2(n2395), .A(n14300), .ZN(n2384) );
  NOR4_X1 U1852 ( .A1(n2531), .A2(n2532), .A3(n2533), .A4(n2534), .ZN(n2530)
         );
  AOI21_X1 U1853 ( .B1(n2559), .B2(n2560), .A(n14294), .ZN(n2531) );
  AOI21_X1 U1854 ( .B1(n2551), .B2(n2552), .A(n14297), .ZN(n2532) );
  AOI21_X1 U1855 ( .B1(n2543), .B2(n2544), .A(n14300), .ZN(n2533) );
  NOR4_X1 U1856 ( .A1(n2680), .A2(n2681), .A3(n2682), .A4(n2683), .ZN(n2679)
         );
  AOI21_X1 U1857 ( .B1(n2708), .B2(n2709), .A(n14294), .ZN(n2680) );
  AOI21_X1 U1858 ( .B1(n2700), .B2(n2701), .A(n14297), .ZN(n2681) );
  AOI21_X1 U1859 ( .B1(n2692), .B2(n2693), .A(n14300), .ZN(n2682) );
  NOR4_X1 U1860 ( .A1(n2829), .A2(n2830), .A3(n2831), .A4(n2832), .ZN(n2828)
         );
  AOI21_X1 U1861 ( .B1(n2857), .B2(n2858), .A(n14294), .ZN(n2829) );
  AOI21_X1 U1862 ( .B1(n2849), .B2(n2850), .A(n14297), .ZN(n2830) );
  AOI21_X1 U1863 ( .B1(n2841), .B2(n2842), .A(n14300), .ZN(n2831) );
  NOR4_X1 U1864 ( .A1(n2978), .A2(n2979), .A3(n2980), .A4(n2981), .ZN(n2977)
         );
  AOI21_X1 U1865 ( .B1(n3006), .B2(n3007), .A(n14294), .ZN(n2978) );
  AOI21_X1 U1866 ( .B1(n2998), .B2(n2999), .A(n14297), .ZN(n2979) );
  AOI21_X1 U1867 ( .B1(n2990), .B2(n2991), .A(n14300), .ZN(n2980) );
  NOR4_X1 U1868 ( .A1(n3127), .A2(n3128), .A3(n3129), .A4(n3130), .ZN(n3126)
         );
  AOI21_X1 U1869 ( .B1(n3155), .B2(n3156), .A(n14295), .ZN(n3127) );
  AOI21_X1 U1870 ( .B1(n3147), .B2(n3148), .A(n14298), .ZN(n3128) );
  AOI21_X1 U1871 ( .B1(n3139), .B2(n3140), .A(n14301), .ZN(n3129) );
  NOR4_X1 U1872 ( .A1(n3276), .A2(n3277), .A3(n3278), .A4(n3279), .ZN(n3275)
         );
  AOI21_X1 U1873 ( .B1(n3304), .B2(n3305), .A(n14295), .ZN(n3276) );
  AOI21_X1 U1874 ( .B1(n3296), .B2(n3297), .A(n14298), .ZN(n3277) );
  AOI21_X1 U1875 ( .B1(n3288), .B2(n3289), .A(n14301), .ZN(n3278) );
  NOR4_X1 U1876 ( .A1(n3425), .A2(n3426), .A3(n3427), .A4(n3428), .ZN(n3424)
         );
  AOI21_X1 U1877 ( .B1(n3453), .B2(n3454), .A(n14295), .ZN(n3425) );
  AOI21_X1 U1878 ( .B1(n3445), .B2(n3446), .A(n14298), .ZN(n3426) );
  AOI21_X1 U1879 ( .B1(n3437), .B2(n3438), .A(n14301), .ZN(n3427) );
  NOR4_X1 U1880 ( .A1(n3574), .A2(n3575), .A3(n3576), .A4(n3577), .ZN(n3573)
         );
  AOI21_X1 U1881 ( .B1(n3602), .B2(n3603), .A(n14295), .ZN(n3574) );
  AOI21_X1 U1882 ( .B1(n3594), .B2(n3595), .A(n14298), .ZN(n3575) );
  AOI21_X1 U1883 ( .B1(n3586), .B2(n3587), .A(n14301), .ZN(n3576) );
  NOR4_X1 U1884 ( .A1(n3723), .A2(n3724), .A3(n3725), .A4(n3726), .ZN(n3722)
         );
  AOI21_X1 U1885 ( .B1(n3751), .B2(n3752), .A(n14295), .ZN(n3723) );
  AOI21_X1 U1886 ( .B1(n3743), .B2(n3744), .A(n14298), .ZN(n3724) );
  AOI21_X1 U1887 ( .B1(n3735), .B2(n3736), .A(n14301), .ZN(n3725) );
  NOR4_X1 U1888 ( .A1(n3872), .A2(n3873), .A3(n3874), .A4(n3875), .ZN(n3871)
         );
  AOI21_X1 U1889 ( .B1(n3900), .B2(n3901), .A(n14295), .ZN(n3872) );
  AOI21_X1 U1890 ( .B1(n3892), .B2(n3893), .A(n14298), .ZN(n3873) );
  AOI21_X1 U1891 ( .B1(n3884), .B2(n3885), .A(n14301), .ZN(n3874) );
  NOR4_X1 U1892 ( .A1(n4021), .A2(n4022), .A3(n4023), .A4(n4024), .ZN(n4020)
         );
  AOI21_X1 U1893 ( .B1(n4049), .B2(n4050), .A(n14295), .ZN(n4021) );
  AOI21_X1 U1894 ( .B1(n4041), .B2(n4042), .A(n14298), .ZN(n4022) );
  AOI21_X1 U1895 ( .B1(n4033), .B2(n4034), .A(n14301), .ZN(n4023) );
  NOR4_X1 U1896 ( .A1(n4170), .A2(n4171), .A3(n4172), .A4(n4173), .ZN(n4169)
         );
  AOI21_X1 U1897 ( .B1(n4198), .B2(n4199), .A(n14295), .ZN(n4170) );
  AOI21_X1 U1898 ( .B1(n4190), .B2(n4191), .A(n14298), .ZN(n4171) );
  AOI21_X1 U1899 ( .B1(n4182), .B2(n4183), .A(n14301), .ZN(n4172) );
  NOR4_X1 U1900 ( .A1(n4319), .A2(n4320), .A3(n4321), .A4(n4322), .ZN(n4318)
         );
  AOI21_X1 U1901 ( .B1(n4347), .B2(n4348), .A(n14295), .ZN(n4319) );
  AOI21_X1 U1902 ( .B1(n4339), .B2(n4340), .A(n14298), .ZN(n4320) );
  AOI21_X1 U1903 ( .B1(n4331), .B2(n4332), .A(n14301), .ZN(n4321) );
  NOR4_X1 U1904 ( .A1(n4468), .A2(n4469), .A3(n4470), .A4(n4471), .ZN(n4467)
         );
  AOI21_X1 U1905 ( .B1(n4496), .B2(n4497), .A(n14295), .ZN(n4468) );
  AOI21_X1 U1906 ( .B1(n4488), .B2(n4489), .A(n14298), .ZN(n4469) );
  AOI21_X1 U1907 ( .B1(n4480), .B2(n4481), .A(n14301), .ZN(n4470) );
  NOR4_X1 U1908 ( .A1(n4617), .A2(n4618), .A3(n4619), .A4(n4620), .ZN(n4616)
         );
  AOI21_X1 U1909 ( .B1(n4645), .B2(n4646), .A(n14295), .ZN(n4617) );
  AOI21_X1 U1910 ( .B1(n4637), .B2(n4638), .A(n14298), .ZN(n4618) );
  AOI21_X1 U1911 ( .B1(n4629), .B2(n4630), .A(n14301), .ZN(n4619) );
  NOR4_X1 U1912 ( .A1(n4766), .A2(n4767), .A3(n4768), .A4(n4769), .ZN(n4765)
         );
  AOI21_X1 U1913 ( .B1(n4794), .B2(n4795), .A(n14295), .ZN(n4766) );
  AOI21_X1 U1914 ( .B1(n4786), .B2(n4787), .A(n14298), .ZN(n4767) );
  AOI21_X1 U1915 ( .B1(n4778), .B2(n4779), .A(n14301), .ZN(n4768) );
  NOR4_X1 U1916 ( .A1(n4915), .A2(n4916), .A3(n4917), .A4(n4918), .ZN(n4914)
         );
  AOI21_X1 U1917 ( .B1(n4943), .B2(n4944), .A(n14295), .ZN(n4915) );
  AOI21_X1 U1918 ( .B1(n4935), .B2(n4936), .A(n14298), .ZN(n4916) );
  AOI21_X1 U1919 ( .B1(n4927), .B2(n4928), .A(n14301), .ZN(n4917) );
  NOR4_X1 U1920 ( .A1(n5064), .A2(n5065), .A3(n5066), .A4(n5067), .ZN(n5063)
         );
  AOI21_X1 U1921 ( .B1(n5092), .B2(n5093), .A(n14296), .ZN(n5064) );
  AOI21_X1 U1922 ( .B1(n5084), .B2(n5085), .A(n14299), .ZN(n5065) );
  AOI21_X1 U1923 ( .B1(n5076), .B2(n5077), .A(n14302), .ZN(n5066) );
  NOR4_X1 U1924 ( .A1(n5213), .A2(n5214), .A3(n5215), .A4(n5216), .ZN(n5212)
         );
  AOI21_X1 U1925 ( .B1(n5241), .B2(n5242), .A(n14296), .ZN(n5213) );
  AOI21_X1 U1926 ( .B1(n5233), .B2(n5234), .A(n14299), .ZN(n5214) );
  AOI21_X1 U1927 ( .B1(n5225), .B2(n5226), .A(n14302), .ZN(n5215) );
  NOR4_X1 U1928 ( .A1(n5362), .A2(n5363), .A3(n5364), .A4(n5365), .ZN(n5361)
         );
  AOI21_X1 U1929 ( .B1(n5390), .B2(n5391), .A(n14296), .ZN(n5362) );
  AOI21_X1 U1930 ( .B1(n5382), .B2(n5383), .A(n14299), .ZN(n5363) );
  AOI21_X1 U1931 ( .B1(n5374), .B2(n5375), .A(n14302), .ZN(n5364) );
  NOR4_X1 U1932 ( .A1(n5511), .A2(n5512), .A3(n5513), .A4(n5514), .ZN(n5510)
         );
  AOI21_X1 U1933 ( .B1(n5539), .B2(n5540), .A(n14296), .ZN(n5511) );
  AOI21_X1 U1934 ( .B1(n5531), .B2(n5532), .A(n14299), .ZN(n5512) );
  AOI21_X1 U1935 ( .B1(n5523), .B2(n5524), .A(n14302), .ZN(n5513) );
  NOR4_X1 U1936 ( .A1(n5660), .A2(n5661), .A3(n5662), .A4(n5663), .ZN(n5659)
         );
  AOI21_X1 U1937 ( .B1(n5688), .B2(n5689), .A(n14296), .ZN(n5660) );
  AOI21_X1 U1938 ( .B1(n5680), .B2(n5681), .A(n14299), .ZN(n5661) );
  AOI21_X1 U1939 ( .B1(n5672), .B2(n5673), .A(n14302), .ZN(n5662) );
  NOR4_X1 U1940 ( .A1(n5809), .A2(n5810), .A3(n5811), .A4(n5812), .ZN(n5808)
         );
  AOI21_X1 U1941 ( .B1(n5829), .B2(n5830), .A(n14299), .ZN(n5810) );
  AOI21_X1 U1942 ( .B1(n5821), .B2(n5822), .A(n14302), .ZN(n5811) );
  AOI21_X1 U1943 ( .B1(n5813), .B2(n5814), .A(n14305), .ZN(n5812) );
  BUF_X1 U1944 ( .A(n501), .Z(n14504) );
  BUF_X1 U1945 ( .A(n501), .Z(n14505) );
  BUF_X1 U1946 ( .A(n501), .Z(n14506) );
  BUF_X1 U1947 ( .A(n501), .Z(n14507) );
  BUF_X1 U1948 ( .A(n501), .Z(n14508) );
  NAND4_X1 U1949 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1169)
         );
  NOR4_X1 U1950 ( .A1(n1294), .A2(n1295), .A3(n1296), .A4(n1297), .ZN(n1170)
         );
  NOR4_X1 U1951 ( .A1(n1254), .A2(n1255), .A3(n1256), .A4(n1257), .ZN(n1171)
         );
  NOR4_X1 U1952 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n1172)
         );
  NAND4_X1 U1953 ( .A1(n1335), .A2(n1336), .A3(n1337), .A4(n1338), .ZN(n1334)
         );
  NOR4_X1 U1954 ( .A1(n1447), .A2(n1448), .A3(n1449), .A4(n1450), .ZN(n1335)
         );
  NOR4_X1 U1955 ( .A1(n1411), .A2(n1412), .A3(n1413), .A4(n1414), .ZN(n1336)
         );
  NOR4_X1 U1956 ( .A1(n1375), .A2(n1376), .A3(n1377), .A4(n1378), .ZN(n1337)
         );
  NAND4_X1 U1957 ( .A1(n1484), .A2(n1485), .A3(n1486), .A4(n1487), .ZN(n1483)
         );
  NOR4_X1 U1958 ( .A1(n1596), .A2(n1597), .A3(n1598), .A4(n1599), .ZN(n1484)
         );
  NOR4_X1 U1959 ( .A1(n1560), .A2(n1561), .A3(n1562), .A4(n1563), .ZN(n1485)
         );
  NOR4_X1 U1960 ( .A1(n1524), .A2(n1525), .A3(n1526), .A4(n1527), .ZN(n1486)
         );
  NAND4_X1 U1961 ( .A1(n1633), .A2(n1634), .A3(n1635), .A4(n1636), .ZN(n1632)
         );
  NOR4_X1 U1962 ( .A1(n1745), .A2(n1746), .A3(n1747), .A4(n1748), .ZN(n1633)
         );
  NOR4_X1 U1963 ( .A1(n1709), .A2(n1710), .A3(n1711), .A4(n1712), .ZN(n1634)
         );
  NOR4_X1 U1964 ( .A1(n1673), .A2(n1674), .A3(n1675), .A4(n1676), .ZN(n1635)
         );
  NAND4_X1 U1965 ( .A1(n1782), .A2(n1783), .A3(n1784), .A4(n1785), .ZN(n1781)
         );
  NOR4_X1 U1966 ( .A1(n1894), .A2(n1895), .A3(n1896), .A4(n1897), .ZN(n1782)
         );
  NOR4_X1 U1967 ( .A1(n1858), .A2(n1859), .A3(n1860), .A4(n1861), .ZN(n1783)
         );
  NOR4_X1 U1968 ( .A1(n1822), .A2(n1823), .A3(n1824), .A4(n1825), .ZN(n1784)
         );
  NAND4_X1 U1969 ( .A1(n1931), .A2(n1932), .A3(n1933), .A4(n1934), .ZN(n1930)
         );
  NOR4_X1 U1970 ( .A1(n2043), .A2(n2044), .A3(n2045), .A4(n2046), .ZN(n1931)
         );
  NOR4_X1 U1971 ( .A1(n2007), .A2(n2008), .A3(n2009), .A4(n2010), .ZN(n1932)
         );
  NOR4_X1 U1972 ( .A1(n1971), .A2(n1972), .A3(n1973), .A4(n1974), .ZN(n1933)
         );
  NAND4_X1 U1973 ( .A1(n2080), .A2(n2081), .A3(n2082), .A4(n2083), .ZN(n2079)
         );
  NOR4_X1 U1974 ( .A1(n2192), .A2(n2193), .A3(n2194), .A4(n2195), .ZN(n2080)
         );
  NOR4_X1 U1975 ( .A1(n2156), .A2(n2157), .A3(n2158), .A4(n2159), .ZN(n2081)
         );
  NOR4_X1 U1976 ( .A1(n2120), .A2(n2121), .A3(n2122), .A4(n2123), .ZN(n2082)
         );
  NAND4_X1 U1977 ( .A1(n2229), .A2(n2230), .A3(n2231), .A4(n2232), .ZN(n2228)
         );
  NOR4_X1 U1978 ( .A1(n2341), .A2(n2342), .A3(n2343), .A4(n2344), .ZN(n2229)
         );
  NOR4_X1 U1979 ( .A1(n2305), .A2(n2306), .A3(n2307), .A4(n2308), .ZN(n2230)
         );
  NOR4_X1 U1980 ( .A1(n2269), .A2(n2270), .A3(n2271), .A4(n2272), .ZN(n2231)
         );
  NAND4_X1 U1981 ( .A1(n2378), .A2(n2379), .A3(n2380), .A4(n2381), .ZN(n2377)
         );
  NOR4_X1 U1982 ( .A1(n2490), .A2(n2491), .A3(n2492), .A4(n2493), .ZN(n2378)
         );
  NOR4_X1 U1983 ( .A1(n2454), .A2(n2455), .A3(n2456), .A4(n2457), .ZN(n2379)
         );
  NOR4_X1 U1984 ( .A1(n2418), .A2(n2419), .A3(n2420), .A4(n2421), .ZN(n2380)
         );
  NAND4_X1 U1985 ( .A1(n2527), .A2(n2528), .A3(n2529), .A4(n2530), .ZN(n2526)
         );
  NOR4_X1 U1986 ( .A1(n2639), .A2(n2640), .A3(n2641), .A4(n2642), .ZN(n2527)
         );
  NOR4_X1 U1987 ( .A1(n2603), .A2(n2604), .A3(n2605), .A4(n2606), .ZN(n2528)
         );
  NOR4_X1 U1988 ( .A1(n2567), .A2(n2568), .A3(n2569), .A4(n2570), .ZN(n2529)
         );
  NAND4_X1 U1989 ( .A1(n2676), .A2(n2677), .A3(n2678), .A4(n2679), .ZN(n2675)
         );
  NOR4_X1 U1990 ( .A1(n2788), .A2(n2789), .A3(n2790), .A4(n2791), .ZN(n2676)
         );
  NOR4_X1 U1991 ( .A1(n2752), .A2(n2753), .A3(n2754), .A4(n2755), .ZN(n2677)
         );
  NOR4_X1 U1992 ( .A1(n2716), .A2(n2717), .A3(n2718), .A4(n2719), .ZN(n2678)
         );
  NAND4_X1 U1993 ( .A1(n2825), .A2(n2826), .A3(n2827), .A4(n2828), .ZN(n2824)
         );
  NOR4_X1 U1994 ( .A1(n2937), .A2(n2938), .A3(n2939), .A4(n2940), .ZN(n2825)
         );
  NOR4_X1 U1995 ( .A1(n2901), .A2(n2902), .A3(n2903), .A4(n2904), .ZN(n2826)
         );
  NOR4_X1 U1996 ( .A1(n2865), .A2(n2866), .A3(n2867), .A4(n2868), .ZN(n2827)
         );
  NAND4_X1 U1997 ( .A1(n2974), .A2(n2975), .A3(n2976), .A4(n2977), .ZN(n2973)
         );
  NOR4_X1 U1998 ( .A1(n3086), .A2(n3087), .A3(n3088), .A4(n3089), .ZN(n2974)
         );
  NOR4_X1 U1999 ( .A1(n3050), .A2(n3051), .A3(n3052), .A4(n3053), .ZN(n2975)
         );
  NOR4_X1 U2000 ( .A1(n3014), .A2(n3015), .A3(n3016), .A4(n3017), .ZN(n2976)
         );
  NAND4_X1 U2001 ( .A1(n3123), .A2(n3124), .A3(n3125), .A4(n3126), .ZN(n3122)
         );
  NOR4_X1 U2002 ( .A1(n3235), .A2(n3236), .A3(n3237), .A4(n3238), .ZN(n3123)
         );
  NOR4_X1 U2003 ( .A1(n3199), .A2(n3200), .A3(n3201), .A4(n3202), .ZN(n3124)
         );
  NOR4_X1 U2004 ( .A1(n3163), .A2(n3164), .A3(n3165), .A4(n3166), .ZN(n3125)
         );
  NAND4_X1 U2005 ( .A1(n3272), .A2(n3273), .A3(n3274), .A4(n3275), .ZN(n3271)
         );
  NOR4_X1 U2006 ( .A1(n3384), .A2(n3385), .A3(n3386), .A4(n3387), .ZN(n3272)
         );
  NOR4_X1 U2007 ( .A1(n3348), .A2(n3349), .A3(n3350), .A4(n3351), .ZN(n3273)
         );
  NOR4_X1 U2008 ( .A1(n3312), .A2(n3313), .A3(n3314), .A4(n3315), .ZN(n3274)
         );
  NAND4_X1 U2009 ( .A1(n3421), .A2(n3422), .A3(n3423), .A4(n3424), .ZN(n3420)
         );
  NOR4_X1 U2010 ( .A1(n3533), .A2(n3534), .A3(n3535), .A4(n3536), .ZN(n3421)
         );
  NOR4_X1 U2011 ( .A1(n3497), .A2(n3498), .A3(n3499), .A4(n3500), .ZN(n3422)
         );
  NOR4_X1 U2012 ( .A1(n3461), .A2(n3462), .A3(n3463), .A4(n3464), .ZN(n3423)
         );
  NAND4_X1 U2013 ( .A1(n3570), .A2(n3571), .A3(n3572), .A4(n3573), .ZN(n3569)
         );
  NOR4_X1 U2014 ( .A1(n3682), .A2(n3683), .A3(n3684), .A4(n3685), .ZN(n3570)
         );
  NOR4_X1 U2015 ( .A1(n3646), .A2(n3647), .A3(n3648), .A4(n3649), .ZN(n3571)
         );
  NOR4_X1 U2016 ( .A1(n3610), .A2(n3611), .A3(n3612), .A4(n3613), .ZN(n3572)
         );
  NAND4_X1 U2017 ( .A1(n3719), .A2(n3720), .A3(n3721), .A4(n3722), .ZN(n3718)
         );
  NOR4_X1 U2018 ( .A1(n3831), .A2(n3832), .A3(n3833), .A4(n3834), .ZN(n3719)
         );
  NOR4_X1 U2019 ( .A1(n3795), .A2(n3796), .A3(n3797), .A4(n3798), .ZN(n3720)
         );
  NOR4_X1 U2020 ( .A1(n3759), .A2(n3760), .A3(n3761), .A4(n3762), .ZN(n3721)
         );
  NAND4_X1 U2021 ( .A1(n3868), .A2(n3869), .A3(n3870), .A4(n3871), .ZN(n3867)
         );
  NOR4_X1 U2022 ( .A1(n3980), .A2(n3981), .A3(n3982), .A4(n3983), .ZN(n3868)
         );
  NOR4_X1 U2023 ( .A1(n3944), .A2(n3945), .A3(n3946), .A4(n3947), .ZN(n3869)
         );
  NOR4_X1 U2024 ( .A1(n3908), .A2(n3909), .A3(n3910), .A4(n3911), .ZN(n3870)
         );
  NAND4_X1 U2025 ( .A1(n4017), .A2(n4018), .A3(n4019), .A4(n4020), .ZN(n4016)
         );
  NOR4_X1 U2026 ( .A1(n4129), .A2(n4130), .A3(n4131), .A4(n4132), .ZN(n4017)
         );
  NOR4_X1 U2027 ( .A1(n4093), .A2(n4094), .A3(n4095), .A4(n4096), .ZN(n4018)
         );
  NOR4_X1 U2028 ( .A1(n4057), .A2(n4058), .A3(n4059), .A4(n4060), .ZN(n4019)
         );
  NAND4_X1 U2029 ( .A1(n4166), .A2(n4167), .A3(n4168), .A4(n4169), .ZN(n4165)
         );
  NOR4_X1 U2030 ( .A1(n4278), .A2(n4279), .A3(n4280), .A4(n4281), .ZN(n4166)
         );
  NOR4_X1 U2031 ( .A1(n4242), .A2(n4243), .A3(n4244), .A4(n4245), .ZN(n4167)
         );
  NOR4_X1 U2032 ( .A1(n4206), .A2(n4207), .A3(n4208), .A4(n4209), .ZN(n4168)
         );
  NAND4_X1 U2033 ( .A1(n4315), .A2(n4316), .A3(n4317), .A4(n4318), .ZN(n4314)
         );
  NOR4_X1 U2034 ( .A1(n4427), .A2(n4428), .A3(n4429), .A4(n4430), .ZN(n4315)
         );
  NOR4_X1 U2035 ( .A1(n4391), .A2(n4392), .A3(n4393), .A4(n4394), .ZN(n4316)
         );
  NOR4_X1 U2036 ( .A1(n4355), .A2(n4356), .A3(n4357), .A4(n4358), .ZN(n4317)
         );
  NAND4_X1 U2037 ( .A1(n4464), .A2(n4465), .A3(n4466), .A4(n4467), .ZN(n4463)
         );
  NOR4_X1 U2038 ( .A1(n4576), .A2(n4577), .A3(n4578), .A4(n4579), .ZN(n4464)
         );
  NOR4_X1 U2039 ( .A1(n4540), .A2(n4541), .A3(n4542), .A4(n4543), .ZN(n4465)
         );
  NOR4_X1 U2040 ( .A1(n4504), .A2(n4505), .A3(n4506), .A4(n4507), .ZN(n4466)
         );
  NAND4_X1 U2041 ( .A1(n4613), .A2(n4614), .A3(n4615), .A4(n4616), .ZN(n4612)
         );
  NOR4_X1 U2042 ( .A1(n4725), .A2(n4726), .A3(n4727), .A4(n4728), .ZN(n4613)
         );
  NOR4_X1 U2043 ( .A1(n4689), .A2(n4690), .A3(n4691), .A4(n4692), .ZN(n4614)
         );
  NOR4_X1 U2044 ( .A1(n4653), .A2(n4654), .A3(n4655), .A4(n4656), .ZN(n4615)
         );
  NAND4_X1 U2045 ( .A1(n4762), .A2(n4763), .A3(n4764), .A4(n4765), .ZN(n4761)
         );
  NOR4_X1 U2046 ( .A1(n4874), .A2(n4875), .A3(n4876), .A4(n4877), .ZN(n4762)
         );
  NOR4_X1 U2047 ( .A1(n4838), .A2(n4839), .A3(n4840), .A4(n4841), .ZN(n4763)
         );
  NOR4_X1 U2048 ( .A1(n4802), .A2(n4803), .A3(n4804), .A4(n4805), .ZN(n4764)
         );
  NAND4_X1 U2049 ( .A1(n4911), .A2(n4912), .A3(n4913), .A4(n4914), .ZN(n4910)
         );
  NOR4_X1 U2050 ( .A1(n5023), .A2(n5024), .A3(n5025), .A4(n5026), .ZN(n4911)
         );
  NOR4_X1 U2051 ( .A1(n4987), .A2(n4988), .A3(n4989), .A4(n4990), .ZN(n4912)
         );
  NOR4_X1 U2052 ( .A1(n4951), .A2(n4952), .A3(n4953), .A4(n4954), .ZN(n4913)
         );
  NAND4_X1 U2053 ( .A1(n5060), .A2(n5061), .A3(n5062), .A4(n5063), .ZN(n5059)
         );
  NOR4_X1 U2054 ( .A1(n5172), .A2(n5173), .A3(n5174), .A4(n5175), .ZN(n5060)
         );
  NOR4_X1 U2055 ( .A1(n5136), .A2(n5137), .A3(n5138), .A4(n5139), .ZN(n5061)
         );
  NOR4_X1 U2056 ( .A1(n5100), .A2(n5101), .A3(n5102), .A4(n5103), .ZN(n5062)
         );
  NAND4_X1 U2057 ( .A1(n5209), .A2(n5210), .A3(n5211), .A4(n5212), .ZN(n5208)
         );
  NOR4_X1 U2058 ( .A1(n5321), .A2(n5322), .A3(n5323), .A4(n5324), .ZN(n5209)
         );
  NOR4_X1 U2059 ( .A1(n5285), .A2(n5286), .A3(n5287), .A4(n5288), .ZN(n5210)
         );
  NOR4_X1 U2060 ( .A1(n5249), .A2(n5250), .A3(n5251), .A4(n5252), .ZN(n5211)
         );
  NAND4_X1 U2061 ( .A1(n5358), .A2(n5359), .A3(n5360), .A4(n5361), .ZN(n5357)
         );
  NOR4_X1 U2062 ( .A1(n5470), .A2(n5471), .A3(n5472), .A4(n5473), .ZN(n5358)
         );
  NOR4_X1 U2063 ( .A1(n5434), .A2(n5435), .A3(n5436), .A4(n5437), .ZN(n5359)
         );
  NOR4_X1 U2064 ( .A1(n5398), .A2(n5399), .A3(n5400), .A4(n5401), .ZN(n5360)
         );
  NAND4_X1 U2065 ( .A1(n5507), .A2(n5508), .A3(n5509), .A4(n5510), .ZN(n5506)
         );
  NOR4_X1 U2066 ( .A1(n5619), .A2(n5620), .A3(n5621), .A4(n5622), .ZN(n5507)
         );
  NOR4_X1 U2067 ( .A1(n5583), .A2(n5584), .A3(n5585), .A4(n5586), .ZN(n5508)
         );
  NOR4_X1 U2068 ( .A1(n5547), .A2(n5548), .A3(n5549), .A4(n5550), .ZN(n5509)
         );
  NAND4_X1 U2069 ( .A1(n5656), .A2(n5657), .A3(n5658), .A4(n5659), .ZN(n5655)
         );
  NOR4_X1 U2070 ( .A1(n5768), .A2(n5769), .A3(n5770), .A4(n5771), .ZN(n5656)
         );
  NOR4_X1 U2071 ( .A1(n5732), .A2(n5733), .A3(n5734), .A4(n5735), .ZN(n5657)
         );
  NOR4_X1 U2072 ( .A1(n5696), .A2(n5697), .A3(n5698), .A4(n5699), .ZN(n5658)
         );
  NAND4_X1 U2073 ( .A1(n5805), .A2(n5806), .A3(n5807), .A4(n5808), .ZN(n5804)
         );
  NOR4_X1 U2074 ( .A1(n5919), .A2(n5920), .A3(n5921), .A4(n5922), .ZN(n5805)
         );
  NOR4_X1 U2075 ( .A1(n5881), .A2(n5882), .A3(n5883), .A4(n5884), .ZN(n5806)
         );
  NOR4_X1 U2076 ( .A1(n5845), .A2(n5846), .A3(n5847), .A4(n5848), .ZN(n5807)
         );
  BUF_X1 U2077 ( .A(n171), .Z(n14644) );
  BUF_X1 U2078 ( .A(n5906), .Z(n14643) );
  BUF_X1 U2079 ( .A(n171), .Z(n14634) );
  BUF_X1 U2080 ( .A(n171), .Z(n14632) );
  BUF_X1 U2081 ( .A(n171), .Z(n14628) );
  BUF_X1 U2082 ( .A(n171), .Z(n14626) );
  BUF_X1 U2083 ( .A(n171), .Z(n14630) );
  BUF_X1 U2084 ( .A(n171), .Z(n14642) );
  BUF_X1 U2085 ( .A(n171), .Z(n14638) );
  BUF_X1 U2086 ( .A(n171), .Z(n14636) );
  BUF_X1 U2087 ( .A(n171), .Z(n14640) );
  BUF_X1 U2088 ( .A(n171), .Z(n14614) );
  BUF_X1 U2089 ( .A(n171), .Z(n14612) );
  BUF_X1 U2090 ( .A(n171), .Z(n14610) );
  BUF_X1 U2091 ( .A(n171), .Z(n14608) );
  BUF_X1 U2092 ( .A(n171), .Z(n14624) );
  BUF_X1 U2093 ( .A(n171), .Z(n14622) );
  BUF_X1 U2094 ( .A(n171), .Z(n14618) );
  BUF_X1 U2095 ( .A(n171), .Z(n14616) );
  BUF_X1 U2096 ( .A(n171), .Z(n14620) );
  BUF_X1 U2097 ( .A(n5906), .Z(n14633) );
  BUF_X1 U2098 ( .A(n5906), .Z(n14631) );
  BUF_X1 U2099 ( .A(n5906), .Z(n14629) );
  BUF_X1 U2100 ( .A(n5906), .Z(n14627) );
  BUF_X1 U2101 ( .A(n5906), .Z(n14641) );
  BUF_X1 U2102 ( .A(n5906), .Z(n14639) );
  BUF_X1 U2103 ( .A(n5906), .Z(n14637) );
  BUF_X1 U2104 ( .A(n5906), .Z(n14635) );
  BUF_X1 U2105 ( .A(n5906), .Z(n14615) );
  BUF_X1 U2106 ( .A(n5906), .Z(n14613) );
  BUF_X1 U2107 ( .A(n5906), .Z(n14609) );
  BUF_X1 U2108 ( .A(n5906), .Z(n14607) );
  BUF_X1 U2109 ( .A(n5906), .Z(n14611) );
  BUF_X1 U2110 ( .A(n5906), .Z(n14623) );
  BUF_X1 U2111 ( .A(n5906), .Z(n14621) );
  BUF_X1 U2112 ( .A(n5906), .Z(n14619) );
  BUF_X1 U2113 ( .A(n5906), .Z(n14617) );
  BUF_X1 U2114 ( .A(n5906), .Z(n14625) );
  OAI22_X1 U2115 ( .A1(n6614), .A2(n1157), .B1(n14929), .B2(n1158), .ZN(n14145) );
  OAI22_X1 U2116 ( .A1(n6598), .A2(n1157), .B1(n14889), .B2(n1158), .ZN(n14146) );
  OAI22_X1 U2117 ( .A1(n6582), .A2(n1157), .B1(n14849), .B2(n1158), .ZN(n14147) );
  OAI22_X1 U2118 ( .A1(n6566), .A2(n1157), .B1(n14809), .B2(n1158), .ZN(n14148) );
  OAI22_X1 U2119 ( .A1(n6550), .A2(n1157), .B1(n14769), .B2(n1158), .ZN(n14149) );
  OAI22_X1 U2120 ( .A1(n6534), .A2(n1157), .B1(n14729), .B2(n1158), .ZN(n14150) );
  OAI22_X1 U2121 ( .A1(n6518), .A2(n1157), .B1(n14689), .B2(n1158), .ZN(n14151) );
  OAI22_X1 U2122 ( .A1(n6486), .A2(n1159), .B1(n14929), .B2(n1160), .ZN(n14153) );
  OAI22_X1 U2123 ( .A1(n6470), .A2(n1159), .B1(n14889), .B2(n1160), .ZN(n14154) );
  OAI22_X1 U2124 ( .A1(n6454), .A2(n1159), .B1(n14849), .B2(n1160), .ZN(n14155) );
  OAI22_X1 U2125 ( .A1(n6438), .A2(n1159), .B1(n14809), .B2(n1160), .ZN(n14156) );
  OAI22_X1 U2126 ( .A1(n6422), .A2(n1159), .B1(n14769), .B2(n1160), .ZN(n14157) );
  OAI22_X1 U2127 ( .A1(n6406), .A2(n1159), .B1(n14729), .B2(n1160), .ZN(n14158) );
  OAI22_X1 U2128 ( .A1(n6390), .A2(n1159), .B1(n14689), .B2(n1160), .ZN(n14159) );
  OAI22_X1 U2129 ( .A1(n6358), .A2(n1162), .B1(n14929), .B2(n1163), .ZN(n14161) );
  OAI22_X1 U2130 ( .A1(n6342), .A2(n1162), .B1(n14889), .B2(n1163), .ZN(n14162) );
  OAI22_X1 U2131 ( .A1(n6326), .A2(n1162), .B1(n14849), .B2(n1163), .ZN(n14163) );
  OAI22_X1 U2132 ( .A1(n6310), .A2(n1162), .B1(n14809), .B2(n1163), .ZN(n14164) );
  OAI22_X1 U2133 ( .A1(n6294), .A2(n1162), .B1(n14769), .B2(n1163), .ZN(n14165) );
  OAI22_X1 U2134 ( .A1(n6278), .A2(n1162), .B1(n14729), .B2(n1163), .ZN(n14166) );
  OAI22_X1 U2135 ( .A1(n6262), .A2(n1162), .B1(n14689), .B2(n1163), .ZN(n14167) );
  OAI22_X1 U2136 ( .A1(n6230), .A2(n1165), .B1(n14929), .B2(n1166), .ZN(n14169) );
  OAI22_X1 U2137 ( .A1(n6214), .A2(n1165), .B1(n14889), .B2(n1166), .ZN(n14170) );
  OAI22_X1 U2138 ( .A1(n6198), .A2(n1165), .B1(n14849), .B2(n1166), .ZN(n14171) );
  OAI22_X1 U2139 ( .A1(n6182), .A2(n1165), .B1(n14809), .B2(n1166), .ZN(n14172) );
  OAI22_X1 U2140 ( .A1(n6166), .A2(n1165), .B1(n14769), .B2(n1166), .ZN(n14173) );
  OAI22_X1 U2141 ( .A1(n6150), .A2(n1165), .B1(n14729), .B2(n1166), .ZN(n14174) );
  OAI22_X1 U2142 ( .A1(n6134), .A2(n1165), .B1(n14689), .B2(n1166), .ZN(n14175) );
  OAI22_X1 U2143 ( .A1(n6102), .A2(n1167), .B1(n14929), .B2(n1168), .ZN(n14177) );
  OAI22_X1 U2144 ( .A1(n6086), .A2(n1167), .B1(n14889), .B2(n1168), .ZN(n14178) );
  OAI22_X1 U2145 ( .A1(n6070), .A2(n1167), .B1(n14849), .B2(n1168), .ZN(n14179) );
  OAI22_X1 U2146 ( .A1(n6054), .A2(n1167), .B1(n14809), .B2(n1168), .ZN(n14180) );
  OAI22_X1 U2147 ( .A1(n6038), .A2(n1167), .B1(n14769), .B2(n1168), .ZN(n14181) );
  OAI22_X1 U2148 ( .A1(n6022), .A2(n1167), .B1(n14729), .B2(n1168), .ZN(n14182) );
  OAI22_X1 U2149 ( .A1(n6006), .A2(n1167), .B1(n14689), .B2(n1168), .ZN(n14183) );
  OAI22_X1 U2150 ( .A1(n14969), .A2(n370), .B1(n10075), .B2(n371), .ZN(n11112)
         );
  OAI22_X1 U2151 ( .A1(n14969), .A2(n373), .B1(n9947), .B2(n374), .ZN(n11120)
         );
  OAI22_X1 U2152 ( .A1(n14969), .A2(n375), .B1(n9819), .B2(n376), .ZN(n11128)
         );
  OAI22_X1 U2153 ( .A1(n14969), .A2(n377), .B1(n9691), .B2(n378), .ZN(n11136)
         );
  OAI22_X1 U2154 ( .A1(n14969), .A2(n379), .B1(n9563), .B2(n380), .ZN(n11144)
         );
  OAI22_X1 U2155 ( .A1(n10081), .A2(n240), .B1(n14954), .B2(n241), .ZN(n10600)
         );
  OAI22_X1 U2156 ( .A1(n10065), .A2(n240), .B1(n14894), .B2(n241), .ZN(n10601)
         );
  OAI22_X1 U2157 ( .A1(n10049), .A2(n240), .B1(n14854), .B2(n241), .ZN(n10602)
         );
  OAI22_X1 U2158 ( .A1(n10033), .A2(n240), .B1(n14814), .B2(n241), .ZN(n10603)
         );
  OAI22_X1 U2159 ( .A1(n10017), .A2(n240), .B1(n14774), .B2(n241), .ZN(n10604)
         );
  OAI22_X1 U2160 ( .A1(n10001), .A2(n240), .B1(n14734), .B2(n241), .ZN(n10605)
         );
  OAI22_X1 U2161 ( .A1(n9985), .A2(n240), .B1(n14694), .B2(n241), .ZN(n10606)
         );
  OAI22_X1 U2162 ( .A1(n9969), .A2(n240), .B1(n14654), .B2(n241), .ZN(n10607)
         );
  OAI22_X1 U2163 ( .A1(n9953), .A2(n243), .B1(n14954), .B2(n244), .ZN(n10608)
         );
  OAI22_X1 U2164 ( .A1(n9937), .A2(n243), .B1(n14895), .B2(n244), .ZN(n10609)
         );
  OAI22_X1 U2165 ( .A1(n9921), .A2(n243), .B1(n14855), .B2(n244), .ZN(n10610)
         );
  OAI22_X1 U2166 ( .A1(n9905), .A2(n243), .B1(n14815), .B2(n244), .ZN(n10611)
         );
  OAI22_X1 U2167 ( .A1(n9889), .A2(n243), .B1(n14775), .B2(n244), .ZN(n10612)
         );
  OAI22_X1 U2168 ( .A1(n9873), .A2(n243), .B1(n14735), .B2(n244), .ZN(n10613)
         );
  OAI22_X1 U2169 ( .A1(n9857), .A2(n243), .B1(n14695), .B2(n244), .ZN(n10614)
         );
  OAI22_X1 U2170 ( .A1(n9841), .A2(n243), .B1(n14655), .B2(n244), .ZN(n10615)
         );
  OAI22_X1 U2171 ( .A1(n9825), .A2(n245), .B1(n14954), .B2(n246), .ZN(n10616)
         );
  OAI22_X1 U2172 ( .A1(n9809), .A2(n245), .B1(n14895), .B2(n246), .ZN(n10617)
         );
  OAI22_X1 U2173 ( .A1(n9793), .A2(n245), .B1(n14855), .B2(n246), .ZN(n10618)
         );
  OAI22_X1 U2174 ( .A1(n9777), .A2(n245), .B1(n14815), .B2(n246), .ZN(n10619)
         );
  OAI22_X1 U2175 ( .A1(n9761), .A2(n245), .B1(n14775), .B2(n246), .ZN(n10620)
         );
  OAI22_X1 U2176 ( .A1(n9745), .A2(n245), .B1(n14735), .B2(n246), .ZN(n10621)
         );
  OAI22_X1 U2177 ( .A1(n9729), .A2(n245), .B1(n14695), .B2(n246), .ZN(n10622)
         );
  OAI22_X1 U2178 ( .A1(n9713), .A2(n245), .B1(n14655), .B2(n246), .ZN(n10623)
         );
  OAI22_X1 U2179 ( .A1(n9697), .A2(n247), .B1(n14954), .B2(n248), .ZN(n10624)
         );
  OAI22_X1 U2180 ( .A1(n9681), .A2(n247), .B1(n14895), .B2(n248), .ZN(n10625)
         );
  OAI22_X1 U2181 ( .A1(n9665), .A2(n247), .B1(n14855), .B2(n248), .ZN(n10626)
         );
  OAI22_X1 U2182 ( .A1(n9649), .A2(n247), .B1(n14815), .B2(n248), .ZN(n10627)
         );
  OAI22_X1 U2183 ( .A1(n9633), .A2(n247), .B1(n14775), .B2(n248), .ZN(n10628)
         );
  OAI22_X1 U2184 ( .A1(n9617), .A2(n247), .B1(n14735), .B2(n248), .ZN(n10629)
         );
  OAI22_X1 U2185 ( .A1(n9601), .A2(n247), .B1(n14695), .B2(n248), .ZN(n10630)
         );
  OAI22_X1 U2186 ( .A1(n9585), .A2(n247), .B1(n14655), .B2(n248), .ZN(n10631)
         );
  OAI22_X1 U2187 ( .A1(n9569), .A2(n249), .B1(n14954), .B2(n250), .ZN(n10632)
         );
  OAI22_X1 U2188 ( .A1(n9553), .A2(n249), .B1(n14895), .B2(n250), .ZN(n10633)
         );
  OAI22_X1 U2189 ( .A1(n9537), .A2(n249), .B1(n14855), .B2(n250), .ZN(n10634)
         );
  OAI22_X1 U2190 ( .A1(n9521), .A2(n249), .B1(n14815), .B2(n250), .ZN(n10635)
         );
  OAI22_X1 U2191 ( .A1(n9505), .A2(n249), .B1(n14775), .B2(n250), .ZN(n10636)
         );
  OAI22_X1 U2192 ( .A1(n9489), .A2(n249), .B1(n14735), .B2(n250), .ZN(n10637)
         );
  OAI22_X1 U2193 ( .A1(n9473), .A2(n249), .B1(n14695), .B2(n250), .ZN(n10638)
         );
  OAI22_X1 U2194 ( .A1(n9457), .A2(n249), .B1(n14655), .B2(n250), .ZN(n10639)
         );
  OAI22_X1 U2195 ( .A1(n9441), .A2(n251), .B1(n14954), .B2(n252), .ZN(n10640)
         );
  OAI22_X1 U2196 ( .A1(n9425), .A2(n251), .B1(n14895), .B2(n252), .ZN(n10641)
         );
  OAI22_X1 U2197 ( .A1(n9409), .A2(n251), .B1(n14855), .B2(n252), .ZN(n10642)
         );
  OAI22_X1 U2198 ( .A1(n9393), .A2(n251), .B1(n14815), .B2(n252), .ZN(n10643)
         );
  OAI22_X1 U2199 ( .A1(n9377), .A2(n251), .B1(n14775), .B2(n252), .ZN(n10644)
         );
  OAI22_X1 U2200 ( .A1(n9361), .A2(n251), .B1(n14735), .B2(n252), .ZN(n10645)
         );
  OAI22_X1 U2201 ( .A1(n9345), .A2(n251), .B1(n14695), .B2(n252), .ZN(n10646)
         );
  OAI22_X1 U2202 ( .A1(n9329), .A2(n251), .B1(n14655), .B2(n252), .ZN(n10647)
         );
  OAI22_X1 U2203 ( .A1(n10083), .A2(n502), .B1(n14964), .B2(n503), .ZN(n11624)
         );
  OAI22_X1 U2204 ( .A1(n10067), .A2(n502), .B1(n14904), .B2(n503), .ZN(n11625)
         );
  OAI22_X1 U2205 ( .A1(n10051), .A2(n502), .B1(n14864), .B2(n503), .ZN(n11626)
         );
  OAI22_X1 U2206 ( .A1(n10035), .A2(n502), .B1(n14824), .B2(n503), .ZN(n11627)
         );
  OAI22_X1 U2207 ( .A1(n10019), .A2(n502), .B1(n14784), .B2(n503), .ZN(n11628)
         );
  OAI22_X1 U2208 ( .A1(n10003), .A2(n502), .B1(n14744), .B2(n503), .ZN(n11629)
         );
  OAI22_X1 U2209 ( .A1(n9987), .A2(n502), .B1(n14704), .B2(n503), .ZN(n11630)
         );
  OAI22_X1 U2210 ( .A1(n9971), .A2(n502), .B1(n14664), .B2(n503), .ZN(n11631)
         );
  OAI22_X1 U2211 ( .A1(n9955), .A2(n505), .B1(n14964), .B2(n506), .ZN(n11632)
         );
  OAI22_X1 U2212 ( .A1(n9939), .A2(n505), .B1(n14904), .B2(n506), .ZN(n11633)
         );
  OAI22_X1 U2213 ( .A1(n9923), .A2(n505), .B1(n14864), .B2(n506), .ZN(n11634)
         );
  OAI22_X1 U2214 ( .A1(n9907), .A2(n505), .B1(n14824), .B2(n506), .ZN(n11635)
         );
  OAI22_X1 U2215 ( .A1(n9891), .A2(n505), .B1(n14784), .B2(n506), .ZN(n11636)
         );
  OAI22_X1 U2216 ( .A1(n9875), .A2(n505), .B1(n14744), .B2(n506), .ZN(n11637)
         );
  OAI22_X1 U2217 ( .A1(n9859), .A2(n505), .B1(n14704), .B2(n506), .ZN(n11638)
         );
  OAI22_X1 U2218 ( .A1(n9843), .A2(n505), .B1(n14664), .B2(n506), .ZN(n11639)
         );
  OAI22_X1 U2219 ( .A1(n9827), .A2(n507), .B1(n14964), .B2(n508), .ZN(n11640)
         );
  OAI22_X1 U2220 ( .A1(n9811), .A2(n507), .B1(n14904), .B2(n508), .ZN(n11641)
         );
  OAI22_X1 U2221 ( .A1(n9795), .A2(n507), .B1(n14864), .B2(n508), .ZN(n11642)
         );
  OAI22_X1 U2222 ( .A1(n9779), .A2(n507), .B1(n14824), .B2(n508), .ZN(n11643)
         );
  OAI22_X1 U2223 ( .A1(n9763), .A2(n507), .B1(n14784), .B2(n508), .ZN(n11644)
         );
  OAI22_X1 U2224 ( .A1(n9747), .A2(n507), .B1(n14744), .B2(n508), .ZN(n11645)
         );
  OAI22_X1 U2225 ( .A1(n9731), .A2(n507), .B1(n14704), .B2(n508), .ZN(n11646)
         );
  OAI22_X1 U2226 ( .A1(n9715), .A2(n507), .B1(n14664), .B2(n508), .ZN(n11647)
         );
  OAI22_X1 U2227 ( .A1(n9699), .A2(n509), .B1(n14964), .B2(n510), .ZN(n11648)
         );
  OAI22_X1 U2228 ( .A1(n9683), .A2(n509), .B1(n14905), .B2(n510), .ZN(n11649)
         );
  OAI22_X1 U2229 ( .A1(n9667), .A2(n509), .B1(n14865), .B2(n510), .ZN(n11650)
         );
  OAI22_X1 U2230 ( .A1(n9651), .A2(n509), .B1(n14825), .B2(n510), .ZN(n11651)
         );
  OAI22_X1 U2231 ( .A1(n9635), .A2(n509), .B1(n14785), .B2(n510), .ZN(n11652)
         );
  OAI22_X1 U2232 ( .A1(n9619), .A2(n509), .B1(n14745), .B2(n510), .ZN(n11653)
         );
  OAI22_X1 U2233 ( .A1(n9603), .A2(n509), .B1(n14705), .B2(n510), .ZN(n11654)
         );
  OAI22_X1 U2234 ( .A1(n9587), .A2(n509), .B1(n14665), .B2(n510), .ZN(n11655)
         );
  OAI22_X1 U2235 ( .A1(n9571), .A2(n511), .B1(n14964), .B2(n512), .ZN(n11656)
         );
  OAI22_X1 U2236 ( .A1(n9555), .A2(n511), .B1(n14905), .B2(n512), .ZN(n11657)
         );
  OAI22_X1 U2237 ( .A1(n9539), .A2(n511), .B1(n14865), .B2(n512), .ZN(n11658)
         );
  OAI22_X1 U2238 ( .A1(n9523), .A2(n511), .B1(n14825), .B2(n512), .ZN(n11659)
         );
  OAI22_X1 U2239 ( .A1(n9507), .A2(n511), .B1(n14785), .B2(n512), .ZN(n11660)
         );
  OAI22_X1 U2240 ( .A1(n9491), .A2(n511), .B1(n14745), .B2(n512), .ZN(n11661)
         );
  OAI22_X1 U2241 ( .A1(n9475), .A2(n511), .B1(n14705), .B2(n512), .ZN(n11662)
         );
  OAI22_X1 U2242 ( .A1(n9459), .A2(n511), .B1(n14665), .B2(n512), .ZN(n11663)
         );
  OAI22_X1 U2243 ( .A1(n9443), .A2(n513), .B1(n14963), .B2(n514), .ZN(n11664)
         );
  OAI22_X1 U2244 ( .A1(n9427), .A2(n513), .B1(n14905), .B2(n514), .ZN(n11665)
         );
  OAI22_X1 U2245 ( .A1(n9411), .A2(n513), .B1(n14865), .B2(n514), .ZN(n11666)
         );
  OAI22_X1 U2246 ( .A1(n9395), .A2(n513), .B1(n14825), .B2(n514), .ZN(n11667)
         );
  OAI22_X1 U2247 ( .A1(n9379), .A2(n513), .B1(n14785), .B2(n514), .ZN(n11668)
         );
  OAI22_X1 U2248 ( .A1(n9363), .A2(n513), .B1(n14745), .B2(n514), .ZN(n11669)
         );
  OAI22_X1 U2249 ( .A1(n9347), .A2(n513), .B1(n14705), .B2(n514), .ZN(n11670)
         );
  OAI22_X1 U2250 ( .A1(n9331), .A2(n513), .B1(n14665), .B2(n514), .ZN(n11671)
         );
  OAI22_X1 U2251 ( .A1(n10087), .A2(n567), .B1(n14961), .B2(n568), .ZN(n11880)
         );
  OAI22_X1 U2252 ( .A1(n10071), .A2(n567), .B1(n14907), .B2(n568), .ZN(n11881)
         );
  OAI22_X1 U2253 ( .A1(n10055), .A2(n567), .B1(n14867), .B2(n568), .ZN(n11882)
         );
  OAI22_X1 U2254 ( .A1(n10039), .A2(n567), .B1(n14827), .B2(n568), .ZN(n11883)
         );
  OAI22_X1 U2255 ( .A1(n10023), .A2(n567), .B1(n14787), .B2(n568), .ZN(n11884)
         );
  OAI22_X1 U2256 ( .A1(n10007), .A2(n567), .B1(n14747), .B2(n568), .ZN(n11885)
         );
  OAI22_X1 U2257 ( .A1(n9991), .A2(n567), .B1(n14707), .B2(n568), .ZN(n11886)
         );
  OAI22_X1 U2258 ( .A1(n9975), .A2(n567), .B1(n14667), .B2(n568), .ZN(n11887)
         );
  OAI22_X1 U2259 ( .A1(n9959), .A2(n570), .B1(n14961), .B2(n571), .ZN(n11888)
         );
  OAI22_X1 U2260 ( .A1(n9943), .A2(n570), .B1(n14907), .B2(n571), .ZN(n11889)
         );
  OAI22_X1 U2261 ( .A1(n9927), .A2(n570), .B1(n14867), .B2(n571), .ZN(n11890)
         );
  OAI22_X1 U2262 ( .A1(n9911), .A2(n570), .B1(n14827), .B2(n571), .ZN(n11891)
         );
  OAI22_X1 U2263 ( .A1(n9895), .A2(n570), .B1(n14787), .B2(n571), .ZN(n11892)
         );
  OAI22_X1 U2264 ( .A1(n9879), .A2(n570), .B1(n14747), .B2(n571), .ZN(n11893)
         );
  OAI22_X1 U2265 ( .A1(n9863), .A2(n570), .B1(n14707), .B2(n571), .ZN(n11894)
         );
  OAI22_X1 U2266 ( .A1(n9847), .A2(n570), .B1(n14667), .B2(n571), .ZN(n11895)
         );
  OAI22_X1 U2267 ( .A1(n9831), .A2(n572), .B1(n14961), .B2(n573), .ZN(n11896)
         );
  OAI22_X1 U2268 ( .A1(n9815), .A2(n572), .B1(n14907), .B2(n573), .ZN(n11897)
         );
  OAI22_X1 U2269 ( .A1(n9799), .A2(n572), .B1(n14867), .B2(n573), .ZN(n11898)
         );
  OAI22_X1 U2270 ( .A1(n9783), .A2(n572), .B1(n14827), .B2(n573), .ZN(n11899)
         );
  OAI22_X1 U2271 ( .A1(n9767), .A2(n572), .B1(n14787), .B2(n573), .ZN(n11900)
         );
  OAI22_X1 U2272 ( .A1(n9751), .A2(n572), .B1(n14747), .B2(n573), .ZN(n11901)
         );
  OAI22_X1 U2273 ( .A1(n9735), .A2(n572), .B1(n14707), .B2(n573), .ZN(n11902)
         );
  OAI22_X1 U2274 ( .A1(n9719), .A2(n572), .B1(n14667), .B2(n573), .ZN(n11903)
         );
  OAI22_X1 U2275 ( .A1(n9703), .A2(n574), .B1(n14961), .B2(n575), .ZN(n11904)
         );
  OAI22_X1 U2276 ( .A1(n9687), .A2(n574), .B1(n14907), .B2(n575), .ZN(n11905)
         );
  OAI22_X1 U2277 ( .A1(n9671), .A2(n574), .B1(n14867), .B2(n575), .ZN(n11906)
         );
  OAI22_X1 U2278 ( .A1(n9655), .A2(n574), .B1(n14827), .B2(n575), .ZN(n11907)
         );
  OAI22_X1 U2279 ( .A1(n9639), .A2(n574), .B1(n14787), .B2(n575), .ZN(n11908)
         );
  OAI22_X1 U2280 ( .A1(n9623), .A2(n574), .B1(n14747), .B2(n575), .ZN(n11909)
         );
  OAI22_X1 U2281 ( .A1(n9607), .A2(n574), .B1(n14707), .B2(n575), .ZN(n11910)
         );
  OAI22_X1 U2282 ( .A1(n9591), .A2(n574), .B1(n14667), .B2(n575), .ZN(n11911)
         );
  OAI22_X1 U2283 ( .A1(n9575), .A2(n576), .B1(n14961), .B2(n577), .ZN(n11912)
         );
  OAI22_X1 U2284 ( .A1(n9559), .A2(n576), .B1(n14907), .B2(n577), .ZN(n11913)
         );
  OAI22_X1 U2285 ( .A1(n9543), .A2(n576), .B1(n14867), .B2(n577), .ZN(n11914)
         );
  OAI22_X1 U2286 ( .A1(n9527), .A2(n576), .B1(n14827), .B2(n577), .ZN(n11915)
         );
  OAI22_X1 U2287 ( .A1(n9511), .A2(n576), .B1(n14787), .B2(n577), .ZN(n11916)
         );
  OAI22_X1 U2288 ( .A1(n9495), .A2(n576), .B1(n14747), .B2(n577), .ZN(n11917)
         );
  OAI22_X1 U2289 ( .A1(n9479), .A2(n576), .B1(n14707), .B2(n577), .ZN(n11918)
         );
  OAI22_X1 U2290 ( .A1(n9463), .A2(n576), .B1(n14667), .B2(n577), .ZN(n11919)
         );
  OAI22_X1 U2291 ( .A1(n9447), .A2(n578), .B1(n14961), .B2(n579), .ZN(n11920)
         );
  OAI22_X1 U2292 ( .A1(n9431), .A2(n578), .B1(n14907), .B2(n579), .ZN(n11921)
         );
  OAI22_X1 U2293 ( .A1(n9415), .A2(n578), .B1(n14867), .B2(n579), .ZN(n11922)
         );
  OAI22_X1 U2294 ( .A1(n9399), .A2(n578), .B1(n14827), .B2(n579), .ZN(n11923)
         );
  OAI22_X1 U2295 ( .A1(n9383), .A2(n578), .B1(n14787), .B2(n579), .ZN(n11924)
         );
  OAI22_X1 U2296 ( .A1(n9367), .A2(n578), .B1(n14747), .B2(n579), .ZN(n11925)
         );
  OAI22_X1 U2297 ( .A1(n9351), .A2(n578), .B1(n14707), .B2(n579), .ZN(n11926)
         );
  OAI22_X1 U2298 ( .A1(n9335), .A2(n578), .B1(n14667), .B2(n579), .ZN(n11927)
         );
  OAI22_X1 U2299 ( .A1(n10082), .A2(n1026), .B1(n14944), .B2(n1027), .ZN(
        n13672) );
  OAI22_X1 U2300 ( .A1(n10066), .A2(n1026), .B1(n14924), .B2(n1027), .ZN(
        n13673) );
  OAI22_X1 U2301 ( .A1(n10050), .A2(n1026), .B1(n14884), .B2(n1027), .ZN(
        n13674) );
  OAI22_X1 U2302 ( .A1(n10034), .A2(n1026), .B1(n14844), .B2(n1027), .ZN(
        n13675) );
  OAI22_X1 U2303 ( .A1(n10018), .A2(n1026), .B1(n14804), .B2(n1027), .ZN(
        n13676) );
  OAI22_X1 U2304 ( .A1(n10002), .A2(n1026), .B1(n14764), .B2(n1027), .ZN(
        n13677) );
  OAI22_X1 U2305 ( .A1(n9986), .A2(n1026), .B1(n14724), .B2(n1027), .ZN(n13678) );
  OAI22_X1 U2306 ( .A1(n9970), .A2(n1026), .B1(n14684), .B2(n1027), .ZN(n13679) );
  OAI22_X1 U2307 ( .A1(n9954), .A2(n1029), .B1(n14944), .B2(n1030), .ZN(n13680) );
  OAI22_X1 U2308 ( .A1(n9938), .A2(n1029), .B1(n14924), .B2(n1030), .ZN(n13681) );
  OAI22_X1 U2309 ( .A1(n9922), .A2(n1029), .B1(n14884), .B2(n1030), .ZN(n13682) );
  OAI22_X1 U2310 ( .A1(n9906), .A2(n1029), .B1(n14844), .B2(n1030), .ZN(n13683) );
  OAI22_X1 U2311 ( .A1(n9890), .A2(n1029), .B1(n14804), .B2(n1030), .ZN(n13684) );
  OAI22_X1 U2312 ( .A1(n9874), .A2(n1029), .B1(n14764), .B2(n1030), .ZN(n13685) );
  OAI22_X1 U2313 ( .A1(n9858), .A2(n1029), .B1(n14724), .B2(n1030), .ZN(n13686) );
  OAI22_X1 U2314 ( .A1(n9842), .A2(n1029), .B1(n14684), .B2(n1030), .ZN(n13687) );
  OAI22_X1 U2315 ( .A1(n9826), .A2(n1031), .B1(n14944), .B2(n1032), .ZN(n13688) );
  OAI22_X1 U2316 ( .A1(n9810), .A2(n1031), .B1(n14924), .B2(n1032), .ZN(n13689) );
  OAI22_X1 U2317 ( .A1(n9794), .A2(n1031), .B1(n14884), .B2(n1032), .ZN(n13690) );
  OAI22_X1 U2318 ( .A1(n9778), .A2(n1031), .B1(n14844), .B2(n1032), .ZN(n13691) );
  OAI22_X1 U2319 ( .A1(n9762), .A2(n1031), .B1(n14804), .B2(n1032), .ZN(n13692) );
  OAI22_X1 U2320 ( .A1(n9746), .A2(n1031), .B1(n14764), .B2(n1032), .ZN(n13693) );
  OAI22_X1 U2321 ( .A1(n9730), .A2(n1031), .B1(n14724), .B2(n1032), .ZN(n13694) );
  OAI22_X1 U2322 ( .A1(n9714), .A2(n1031), .B1(n14684), .B2(n1032), .ZN(n13695) );
  OAI22_X1 U2323 ( .A1(n9698), .A2(n1033), .B1(n14944), .B2(n1034), .ZN(n13696) );
  OAI22_X1 U2324 ( .A1(n9682), .A2(n1033), .B1(n14924), .B2(n1034), .ZN(n13697) );
  OAI22_X1 U2325 ( .A1(n9666), .A2(n1033), .B1(n14884), .B2(n1034), .ZN(n13698) );
  OAI22_X1 U2326 ( .A1(n9650), .A2(n1033), .B1(n14844), .B2(n1034), .ZN(n13699) );
  OAI22_X1 U2327 ( .A1(n9634), .A2(n1033), .B1(n14804), .B2(n1034), .ZN(n13700) );
  OAI22_X1 U2328 ( .A1(n9618), .A2(n1033), .B1(n14764), .B2(n1034), .ZN(n13701) );
  OAI22_X1 U2329 ( .A1(n9602), .A2(n1033), .B1(n14724), .B2(n1034), .ZN(n13702) );
  OAI22_X1 U2330 ( .A1(n9586), .A2(n1033), .B1(n14684), .B2(n1034), .ZN(n13703) );
  OAI22_X1 U2331 ( .A1(n9570), .A2(n1035), .B1(n14944), .B2(n1036), .ZN(n13704) );
  OAI22_X1 U2332 ( .A1(n9554), .A2(n1035), .B1(n14924), .B2(n1036), .ZN(n13705) );
  OAI22_X1 U2333 ( .A1(n9538), .A2(n1035), .B1(n14884), .B2(n1036), .ZN(n13706) );
  OAI22_X1 U2334 ( .A1(n9522), .A2(n1035), .B1(n14844), .B2(n1036), .ZN(n13707) );
  OAI22_X1 U2335 ( .A1(n9506), .A2(n1035), .B1(n14804), .B2(n1036), .ZN(n13708) );
  OAI22_X1 U2336 ( .A1(n9490), .A2(n1035), .B1(n14764), .B2(n1036), .ZN(n13709) );
  OAI22_X1 U2337 ( .A1(n9474), .A2(n1035), .B1(n14724), .B2(n1036), .ZN(n13710) );
  OAI22_X1 U2338 ( .A1(n9458), .A2(n1035), .B1(n14684), .B2(n1036), .ZN(n13711) );
  OAI22_X1 U2339 ( .A1(n9442), .A2(n1037), .B1(n14944), .B2(n1038), .ZN(n13712) );
  OAI22_X1 U2340 ( .A1(n9426), .A2(n1037), .B1(n14924), .B2(n1038), .ZN(n13713) );
  OAI22_X1 U2341 ( .A1(n9410), .A2(n1037), .B1(n14884), .B2(n1038), .ZN(n13714) );
  OAI22_X1 U2342 ( .A1(n9394), .A2(n1037), .B1(n14844), .B2(n1038), .ZN(n13715) );
  OAI22_X1 U2343 ( .A1(n9378), .A2(n1037), .B1(n14804), .B2(n1038), .ZN(n13716) );
  OAI22_X1 U2344 ( .A1(n9362), .A2(n1037), .B1(n14764), .B2(n1038), .ZN(n13717) );
  OAI22_X1 U2345 ( .A1(n9346), .A2(n1037), .B1(n14724), .B2(n1038), .ZN(n13718) );
  OAI22_X1 U2346 ( .A1(n9330), .A2(n1037), .B1(n14684), .B2(n1038), .ZN(n13719) );
  OAI22_X1 U2347 ( .A1(n6749), .A2(n226), .B1(n14955), .B2(n227), .ZN(n10552)
         );
  OAI22_X1 U2348 ( .A1(n6733), .A2(n226), .B1(n14894), .B2(n227), .ZN(n10553)
         );
  OAI22_X1 U2349 ( .A1(n6717), .A2(n226), .B1(n14854), .B2(n227), .ZN(n10554)
         );
  OAI22_X1 U2350 ( .A1(n6701), .A2(n226), .B1(n14814), .B2(n227), .ZN(n10555)
         );
  OAI22_X1 U2351 ( .A1(n6685), .A2(n226), .B1(n14774), .B2(n227), .ZN(n10556)
         );
  OAI22_X1 U2352 ( .A1(n6669), .A2(n226), .B1(n14734), .B2(n227), .ZN(n10557)
         );
  OAI22_X1 U2353 ( .A1(n6653), .A2(n226), .B1(n14694), .B2(n227), .ZN(n10558)
         );
  OAI22_X1 U2354 ( .A1(n6637), .A2(n226), .B1(n14654), .B2(n227), .ZN(n10559)
         );
  OAI22_X1 U2355 ( .A1(n6621), .A2(n228), .B1(n14955), .B2(n229), .ZN(n10560)
         );
  OAI22_X1 U2356 ( .A1(n6605), .A2(n228), .B1(n14894), .B2(n229), .ZN(n10561)
         );
  OAI22_X1 U2357 ( .A1(n6589), .A2(n228), .B1(n14854), .B2(n229), .ZN(n10562)
         );
  OAI22_X1 U2358 ( .A1(n6573), .A2(n228), .B1(n14814), .B2(n229), .ZN(n10563)
         );
  OAI22_X1 U2359 ( .A1(n6557), .A2(n228), .B1(n14774), .B2(n229), .ZN(n10564)
         );
  OAI22_X1 U2360 ( .A1(n6541), .A2(n228), .B1(n14734), .B2(n229), .ZN(n10565)
         );
  OAI22_X1 U2361 ( .A1(n6525), .A2(n228), .B1(n14694), .B2(n229), .ZN(n10566)
         );
  OAI22_X1 U2362 ( .A1(n6509), .A2(n228), .B1(n14654), .B2(n229), .ZN(n10567)
         );
  OAI22_X1 U2363 ( .A1(n6493), .A2(n230), .B1(n14954), .B2(n231), .ZN(n10568)
         );
  OAI22_X1 U2364 ( .A1(n6477), .A2(n230), .B1(n14894), .B2(n231), .ZN(n10569)
         );
  OAI22_X1 U2365 ( .A1(n6461), .A2(n230), .B1(n14854), .B2(n231), .ZN(n10570)
         );
  OAI22_X1 U2366 ( .A1(n6445), .A2(n230), .B1(n14814), .B2(n231), .ZN(n10571)
         );
  OAI22_X1 U2367 ( .A1(n6429), .A2(n230), .B1(n14774), .B2(n231), .ZN(n10572)
         );
  OAI22_X1 U2368 ( .A1(n6413), .A2(n230), .B1(n14734), .B2(n231), .ZN(n10573)
         );
  OAI22_X1 U2369 ( .A1(n6397), .A2(n230), .B1(n14694), .B2(n231), .ZN(n10574)
         );
  OAI22_X1 U2370 ( .A1(n6381), .A2(n230), .B1(n14654), .B2(n231), .ZN(n10575)
         );
  OAI22_X1 U2371 ( .A1(n6365), .A2(n232), .B1(n14954), .B2(n233), .ZN(n10576)
         );
  OAI22_X1 U2372 ( .A1(n6349), .A2(n232), .B1(n14894), .B2(n233), .ZN(n10577)
         );
  OAI22_X1 U2373 ( .A1(n6333), .A2(n232), .B1(n14854), .B2(n233), .ZN(n10578)
         );
  OAI22_X1 U2374 ( .A1(n6317), .A2(n232), .B1(n14814), .B2(n233), .ZN(n10579)
         );
  OAI22_X1 U2375 ( .A1(n6301), .A2(n232), .B1(n14774), .B2(n233), .ZN(n10580)
         );
  OAI22_X1 U2376 ( .A1(n6285), .A2(n232), .B1(n14734), .B2(n233), .ZN(n10581)
         );
  OAI22_X1 U2377 ( .A1(n6269), .A2(n232), .B1(n14694), .B2(n233), .ZN(n10582)
         );
  OAI22_X1 U2378 ( .A1(n6253), .A2(n232), .B1(n14654), .B2(n233), .ZN(n10583)
         );
  OAI22_X1 U2379 ( .A1(n6237), .A2(n234), .B1(n14954), .B2(n235), .ZN(n10584)
         );
  OAI22_X1 U2380 ( .A1(n6221), .A2(n234), .B1(n14894), .B2(n235), .ZN(n10585)
         );
  OAI22_X1 U2381 ( .A1(n6205), .A2(n234), .B1(n14854), .B2(n235), .ZN(n10586)
         );
  OAI22_X1 U2382 ( .A1(n6189), .A2(n234), .B1(n14814), .B2(n235), .ZN(n10587)
         );
  OAI22_X1 U2383 ( .A1(n6173), .A2(n234), .B1(n14774), .B2(n235), .ZN(n10588)
         );
  OAI22_X1 U2384 ( .A1(n6157), .A2(n234), .B1(n14734), .B2(n235), .ZN(n10589)
         );
  OAI22_X1 U2385 ( .A1(n6141), .A2(n234), .B1(n14694), .B2(n235), .ZN(n10590)
         );
  OAI22_X1 U2386 ( .A1(n6125), .A2(n234), .B1(n14654), .B2(n235), .ZN(n10591)
         );
  OAI22_X1 U2387 ( .A1(n6109), .A2(n236), .B1(n14954), .B2(n237), .ZN(n10592)
         );
  OAI22_X1 U2388 ( .A1(n6093), .A2(n236), .B1(n14894), .B2(n237), .ZN(n10593)
         );
  OAI22_X1 U2389 ( .A1(n6077), .A2(n236), .B1(n14854), .B2(n237), .ZN(n10594)
         );
  OAI22_X1 U2390 ( .A1(n6061), .A2(n236), .B1(n14814), .B2(n237), .ZN(n10595)
         );
  OAI22_X1 U2391 ( .A1(n6045), .A2(n236), .B1(n14774), .B2(n237), .ZN(n10596)
         );
  OAI22_X1 U2392 ( .A1(n6029), .A2(n236), .B1(n14734), .B2(n237), .ZN(n10597)
         );
  OAI22_X1 U2393 ( .A1(n6013), .A2(n236), .B1(n14694), .B2(n237), .ZN(n10598)
         );
  OAI22_X1 U2394 ( .A1(n5997), .A2(n236), .B1(n14654), .B2(n237), .ZN(n10599)
         );
  OAI22_X1 U2395 ( .A1(n6757), .A2(n358), .B1(n14950), .B2(n359), .ZN(n11064)
         );
  OAI22_X1 U2396 ( .A1(n6741), .A2(n358), .B1(n14899), .B2(n359), .ZN(n11065)
         );
  OAI22_X1 U2397 ( .A1(n6725), .A2(n358), .B1(n14859), .B2(n359), .ZN(n11066)
         );
  OAI22_X1 U2398 ( .A1(n6709), .A2(n358), .B1(n14819), .B2(n359), .ZN(n11067)
         );
  OAI22_X1 U2399 ( .A1(n6693), .A2(n358), .B1(n14779), .B2(n359), .ZN(n11068)
         );
  OAI22_X1 U2400 ( .A1(n6677), .A2(n358), .B1(n14739), .B2(n359), .ZN(n11069)
         );
  OAI22_X1 U2401 ( .A1(n6661), .A2(n358), .B1(n14699), .B2(n359), .ZN(n11070)
         );
  OAI22_X1 U2402 ( .A1(n6645), .A2(n358), .B1(n14659), .B2(n359), .ZN(n11071)
         );
  OAI22_X1 U2403 ( .A1(n6629), .A2(n360), .B1(n14950), .B2(n361), .ZN(n11072)
         );
  OAI22_X1 U2404 ( .A1(n6613), .A2(n360), .B1(n14899), .B2(n361), .ZN(n11073)
         );
  OAI22_X1 U2405 ( .A1(n6597), .A2(n360), .B1(n14859), .B2(n361), .ZN(n11074)
         );
  OAI22_X1 U2406 ( .A1(n6581), .A2(n360), .B1(n14819), .B2(n361), .ZN(n11075)
         );
  OAI22_X1 U2407 ( .A1(n6565), .A2(n360), .B1(n14779), .B2(n361), .ZN(n11076)
         );
  OAI22_X1 U2408 ( .A1(n6549), .A2(n360), .B1(n14739), .B2(n361), .ZN(n11077)
         );
  OAI22_X1 U2409 ( .A1(n6533), .A2(n360), .B1(n14699), .B2(n361), .ZN(n11078)
         );
  OAI22_X1 U2410 ( .A1(n6517), .A2(n360), .B1(n14659), .B2(n361), .ZN(n11079)
         );
  OAI22_X1 U2411 ( .A1(n6501), .A2(n362), .B1(n14949), .B2(n363), .ZN(n11080)
         );
  OAI22_X1 U2412 ( .A1(n6485), .A2(n362), .B1(n14899), .B2(n363), .ZN(n11081)
         );
  OAI22_X1 U2413 ( .A1(n6469), .A2(n362), .B1(n14859), .B2(n363), .ZN(n11082)
         );
  OAI22_X1 U2414 ( .A1(n6453), .A2(n362), .B1(n14819), .B2(n363), .ZN(n11083)
         );
  OAI22_X1 U2415 ( .A1(n6437), .A2(n362), .B1(n14779), .B2(n363), .ZN(n11084)
         );
  OAI22_X1 U2416 ( .A1(n6421), .A2(n362), .B1(n14739), .B2(n363), .ZN(n11085)
         );
  OAI22_X1 U2417 ( .A1(n6405), .A2(n362), .B1(n14699), .B2(n363), .ZN(n11086)
         );
  OAI22_X1 U2418 ( .A1(n6389), .A2(n362), .B1(n14659), .B2(n363), .ZN(n11087)
         );
  OAI22_X1 U2419 ( .A1(n6373), .A2(n364), .B1(n14949), .B2(n365), .ZN(n11088)
         );
  OAI22_X1 U2420 ( .A1(n6357), .A2(n364), .B1(n14899), .B2(n365), .ZN(n11089)
         );
  OAI22_X1 U2421 ( .A1(n6341), .A2(n364), .B1(n14859), .B2(n365), .ZN(n11090)
         );
  OAI22_X1 U2422 ( .A1(n6325), .A2(n364), .B1(n14819), .B2(n365), .ZN(n11091)
         );
  OAI22_X1 U2423 ( .A1(n6309), .A2(n364), .B1(n14779), .B2(n365), .ZN(n11092)
         );
  OAI22_X1 U2424 ( .A1(n6293), .A2(n364), .B1(n14739), .B2(n365), .ZN(n11093)
         );
  OAI22_X1 U2425 ( .A1(n6277), .A2(n364), .B1(n14699), .B2(n365), .ZN(n11094)
         );
  OAI22_X1 U2426 ( .A1(n6261), .A2(n364), .B1(n14659), .B2(n365), .ZN(n11095)
         );
  OAI22_X1 U2427 ( .A1(n6245), .A2(n366), .B1(n14949), .B2(n367), .ZN(n11096)
         );
  OAI22_X1 U2428 ( .A1(n6229), .A2(n366), .B1(n14899), .B2(n367), .ZN(n11097)
         );
  OAI22_X1 U2429 ( .A1(n6213), .A2(n366), .B1(n14859), .B2(n367), .ZN(n11098)
         );
  OAI22_X1 U2430 ( .A1(n6197), .A2(n366), .B1(n14819), .B2(n367), .ZN(n11099)
         );
  OAI22_X1 U2431 ( .A1(n6181), .A2(n366), .B1(n14779), .B2(n367), .ZN(n11100)
         );
  OAI22_X1 U2432 ( .A1(n6165), .A2(n366), .B1(n14739), .B2(n367), .ZN(n11101)
         );
  OAI22_X1 U2433 ( .A1(n6149), .A2(n366), .B1(n14699), .B2(n367), .ZN(n11102)
         );
  OAI22_X1 U2434 ( .A1(n6133), .A2(n366), .B1(n14659), .B2(n367), .ZN(n11103)
         );
  OAI22_X1 U2435 ( .A1(n6117), .A2(n368), .B1(n14954), .B2(n369), .ZN(n11104)
         );
  OAI22_X1 U2436 ( .A1(n6101), .A2(n368), .B1(n14899), .B2(n369), .ZN(n11105)
         );
  OAI22_X1 U2437 ( .A1(n6085), .A2(n368), .B1(n14859), .B2(n369), .ZN(n11106)
         );
  OAI22_X1 U2438 ( .A1(n6069), .A2(n368), .B1(n14819), .B2(n369), .ZN(n11107)
         );
  OAI22_X1 U2439 ( .A1(n6053), .A2(n368), .B1(n14779), .B2(n369), .ZN(n11108)
         );
  OAI22_X1 U2440 ( .A1(n6037), .A2(n368), .B1(n14739), .B2(n369), .ZN(n11109)
         );
  OAI22_X1 U2441 ( .A1(n6021), .A2(n368), .B1(n14699), .B2(n369), .ZN(n11110)
         );
  OAI22_X1 U2442 ( .A1(n6005), .A2(n368), .B1(n14659), .B2(n369), .ZN(n11111)
         );
  OAI22_X1 U2443 ( .A1(n10059), .A2(n371), .B1(n14899), .B2(n370), .ZN(n11113)
         );
  OAI22_X1 U2444 ( .A1(n10043), .A2(n371), .B1(n14859), .B2(n370), .ZN(n11114)
         );
  OAI22_X1 U2445 ( .A1(n10027), .A2(n371), .B1(n14819), .B2(n370), .ZN(n11115)
         );
  OAI22_X1 U2446 ( .A1(n10011), .A2(n371), .B1(n14779), .B2(n370), .ZN(n11116)
         );
  OAI22_X1 U2447 ( .A1(n9995), .A2(n371), .B1(n14739), .B2(n370), .ZN(n11117)
         );
  OAI22_X1 U2448 ( .A1(n9979), .A2(n371), .B1(n14699), .B2(n370), .ZN(n11118)
         );
  OAI22_X1 U2449 ( .A1(n9963), .A2(n371), .B1(n14659), .B2(n370), .ZN(n11119)
         );
  OAI22_X1 U2450 ( .A1(n9931), .A2(n374), .B1(n14899), .B2(n373), .ZN(n11121)
         );
  OAI22_X1 U2451 ( .A1(n9915), .A2(n374), .B1(n14859), .B2(n373), .ZN(n11122)
         );
  OAI22_X1 U2452 ( .A1(n9899), .A2(n374), .B1(n14819), .B2(n373), .ZN(n11123)
         );
  OAI22_X1 U2453 ( .A1(n9883), .A2(n374), .B1(n14779), .B2(n373), .ZN(n11124)
         );
  OAI22_X1 U2454 ( .A1(n9867), .A2(n374), .B1(n14739), .B2(n373), .ZN(n11125)
         );
  OAI22_X1 U2455 ( .A1(n9851), .A2(n374), .B1(n14699), .B2(n373), .ZN(n11126)
         );
  OAI22_X1 U2456 ( .A1(n9835), .A2(n374), .B1(n14659), .B2(n373), .ZN(n11127)
         );
  OAI22_X1 U2457 ( .A1(n9803), .A2(n376), .B1(n14900), .B2(n375), .ZN(n11129)
         );
  OAI22_X1 U2458 ( .A1(n9787), .A2(n376), .B1(n14860), .B2(n375), .ZN(n11130)
         );
  OAI22_X1 U2459 ( .A1(n9771), .A2(n376), .B1(n14820), .B2(n375), .ZN(n11131)
         );
  OAI22_X1 U2460 ( .A1(n9755), .A2(n376), .B1(n14780), .B2(n375), .ZN(n11132)
         );
  OAI22_X1 U2461 ( .A1(n9739), .A2(n376), .B1(n14740), .B2(n375), .ZN(n11133)
         );
  OAI22_X1 U2462 ( .A1(n9723), .A2(n376), .B1(n14700), .B2(n375), .ZN(n11134)
         );
  OAI22_X1 U2463 ( .A1(n9707), .A2(n376), .B1(n14660), .B2(n375), .ZN(n11135)
         );
  OAI22_X1 U2464 ( .A1(n9675), .A2(n378), .B1(n14900), .B2(n377), .ZN(n11137)
         );
  OAI22_X1 U2465 ( .A1(n9659), .A2(n378), .B1(n14860), .B2(n377), .ZN(n11138)
         );
  OAI22_X1 U2466 ( .A1(n9643), .A2(n378), .B1(n14820), .B2(n377), .ZN(n11139)
         );
  OAI22_X1 U2467 ( .A1(n9627), .A2(n378), .B1(n14780), .B2(n377), .ZN(n11140)
         );
  OAI22_X1 U2468 ( .A1(n9611), .A2(n378), .B1(n14740), .B2(n377), .ZN(n11141)
         );
  OAI22_X1 U2469 ( .A1(n9595), .A2(n378), .B1(n14700), .B2(n377), .ZN(n11142)
         );
  OAI22_X1 U2470 ( .A1(n9579), .A2(n378), .B1(n14660), .B2(n377), .ZN(n11143)
         );
  OAI22_X1 U2471 ( .A1(n9547), .A2(n380), .B1(n14900), .B2(n379), .ZN(n11145)
         );
  OAI22_X1 U2472 ( .A1(n9531), .A2(n380), .B1(n14860), .B2(n379), .ZN(n11146)
         );
  OAI22_X1 U2473 ( .A1(n9515), .A2(n380), .B1(n14820), .B2(n379), .ZN(n11147)
         );
  OAI22_X1 U2474 ( .A1(n9499), .A2(n380), .B1(n14780), .B2(n379), .ZN(n11148)
         );
  OAI22_X1 U2475 ( .A1(n9483), .A2(n380), .B1(n14740), .B2(n379), .ZN(n11149)
         );
  OAI22_X1 U2476 ( .A1(n9467), .A2(n380), .B1(n14700), .B2(n379), .ZN(n11150)
         );
  OAI22_X1 U2477 ( .A1(n9451), .A2(n380), .B1(n14660), .B2(n379), .ZN(n11151)
         );
  OAI22_X1 U2478 ( .A1(n9419), .A2(n382), .B1(n14900), .B2(n381), .ZN(n11153)
         );
  OAI22_X1 U2479 ( .A1(n9403), .A2(n382), .B1(n14860), .B2(n381), .ZN(n11154)
         );
  OAI22_X1 U2480 ( .A1(n9387), .A2(n382), .B1(n14820), .B2(n381), .ZN(n11155)
         );
  OAI22_X1 U2481 ( .A1(n9371), .A2(n382), .B1(n14780), .B2(n381), .ZN(n11156)
         );
  OAI22_X1 U2482 ( .A1(n9355), .A2(n382), .B1(n14740), .B2(n381), .ZN(n11157)
         );
  OAI22_X1 U2483 ( .A1(n9339), .A2(n382), .B1(n14700), .B2(n381), .ZN(n11158)
         );
  OAI22_X1 U2484 ( .A1(n9323), .A2(n382), .B1(n14660), .B2(n381), .ZN(n11159)
         );
  OAI22_X1 U2485 ( .A1(n6744), .A2(n685), .B1(n14937), .B2(n686), .ZN(n12344)
         );
  OAI22_X1 U2486 ( .A1(n6728), .A2(n685), .B1(n14911), .B2(n686), .ZN(n12345)
         );
  OAI22_X1 U2487 ( .A1(n6712), .A2(n685), .B1(n14871), .B2(n686), .ZN(n12346)
         );
  OAI22_X1 U2488 ( .A1(n6696), .A2(n685), .B1(n14831), .B2(n686), .ZN(n12347)
         );
  OAI22_X1 U2489 ( .A1(n6680), .A2(n685), .B1(n14791), .B2(n686), .ZN(n12348)
         );
  OAI22_X1 U2490 ( .A1(n6664), .A2(n685), .B1(n14751), .B2(n686), .ZN(n12349)
         );
  OAI22_X1 U2491 ( .A1(n6648), .A2(n685), .B1(n14711), .B2(n686), .ZN(n12350)
         );
  OAI22_X1 U2492 ( .A1(n6632), .A2(n685), .B1(n14671), .B2(n686), .ZN(n12351)
         );
  OAI22_X1 U2493 ( .A1(n6616), .A2(n687), .B1(n14937), .B2(n688), .ZN(n12352)
         );
  OAI22_X1 U2494 ( .A1(n6600), .A2(n687), .B1(n14911), .B2(n688), .ZN(n12353)
         );
  OAI22_X1 U2495 ( .A1(n6584), .A2(n687), .B1(n14871), .B2(n688), .ZN(n12354)
         );
  OAI22_X1 U2496 ( .A1(n6568), .A2(n687), .B1(n14831), .B2(n688), .ZN(n12355)
         );
  OAI22_X1 U2497 ( .A1(n6552), .A2(n687), .B1(n14791), .B2(n688), .ZN(n12356)
         );
  OAI22_X1 U2498 ( .A1(n6536), .A2(n687), .B1(n14751), .B2(n688), .ZN(n12357)
         );
  OAI22_X1 U2499 ( .A1(n6520), .A2(n687), .B1(n14711), .B2(n688), .ZN(n12358)
         );
  OAI22_X1 U2500 ( .A1(n6504), .A2(n687), .B1(n14671), .B2(n688), .ZN(n12359)
         );
  OAI22_X1 U2501 ( .A1(n6488), .A2(n689), .B1(n14937), .B2(n690), .ZN(n12360)
         );
  OAI22_X1 U2502 ( .A1(n6472), .A2(n689), .B1(n14911), .B2(n690), .ZN(n12361)
         );
  OAI22_X1 U2503 ( .A1(n6456), .A2(n689), .B1(n14871), .B2(n690), .ZN(n12362)
         );
  OAI22_X1 U2504 ( .A1(n6440), .A2(n689), .B1(n14831), .B2(n690), .ZN(n12363)
         );
  OAI22_X1 U2505 ( .A1(n6424), .A2(n689), .B1(n14791), .B2(n690), .ZN(n12364)
         );
  OAI22_X1 U2506 ( .A1(n6408), .A2(n689), .B1(n14751), .B2(n690), .ZN(n12365)
         );
  OAI22_X1 U2507 ( .A1(n6392), .A2(n689), .B1(n14711), .B2(n690), .ZN(n12366)
         );
  OAI22_X1 U2508 ( .A1(n6376), .A2(n689), .B1(n14671), .B2(n690), .ZN(n12367)
         );
  OAI22_X1 U2509 ( .A1(n6360), .A2(n691), .B1(n14937), .B2(n692), .ZN(n12368)
         );
  OAI22_X1 U2510 ( .A1(n6344), .A2(n691), .B1(n14911), .B2(n692), .ZN(n12369)
         );
  OAI22_X1 U2511 ( .A1(n6328), .A2(n691), .B1(n14871), .B2(n692), .ZN(n12370)
         );
  OAI22_X1 U2512 ( .A1(n6312), .A2(n691), .B1(n14831), .B2(n692), .ZN(n12371)
         );
  OAI22_X1 U2513 ( .A1(n6296), .A2(n691), .B1(n14791), .B2(n692), .ZN(n12372)
         );
  OAI22_X1 U2514 ( .A1(n6280), .A2(n691), .B1(n14751), .B2(n692), .ZN(n12373)
         );
  OAI22_X1 U2515 ( .A1(n6264), .A2(n691), .B1(n14711), .B2(n692), .ZN(n12374)
         );
  OAI22_X1 U2516 ( .A1(n6248), .A2(n691), .B1(n14671), .B2(n692), .ZN(n12375)
         );
  OAI22_X1 U2517 ( .A1(n6232), .A2(n693), .B1(n14937), .B2(n694), .ZN(n12376)
         );
  OAI22_X1 U2518 ( .A1(n6216), .A2(n693), .B1(n14912), .B2(n694), .ZN(n12377)
         );
  OAI22_X1 U2519 ( .A1(n6200), .A2(n693), .B1(n14872), .B2(n694), .ZN(n12378)
         );
  OAI22_X1 U2520 ( .A1(n6184), .A2(n693), .B1(n14832), .B2(n694), .ZN(n12379)
         );
  OAI22_X1 U2521 ( .A1(n6168), .A2(n693), .B1(n14792), .B2(n694), .ZN(n12380)
         );
  OAI22_X1 U2522 ( .A1(n6152), .A2(n693), .B1(n14752), .B2(n694), .ZN(n12381)
         );
  OAI22_X1 U2523 ( .A1(n6136), .A2(n693), .B1(n14712), .B2(n694), .ZN(n12382)
         );
  OAI22_X1 U2524 ( .A1(n6120), .A2(n693), .B1(n14672), .B2(n694), .ZN(n12383)
         );
  OAI22_X1 U2525 ( .A1(n6104), .A2(n695), .B1(n14937), .B2(n696), .ZN(n12384)
         );
  OAI22_X1 U2526 ( .A1(n6088), .A2(n695), .B1(n14912), .B2(n696), .ZN(n12385)
         );
  OAI22_X1 U2527 ( .A1(n6072), .A2(n695), .B1(n14872), .B2(n696), .ZN(n12386)
         );
  OAI22_X1 U2528 ( .A1(n6056), .A2(n695), .B1(n14832), .B2(n696), .ZN(n12387)
         );
  OAI22_X1 U2529 ( .A1(n6040), .A2(n695), .B1(n14792), .B2(n696), .ZN(n12388)
         );
  OAI22_X1 U2530 ( .A1(n6024), .A2(n695), .B1(n14752), .B2(n696), .ZN(n12389)
         );
  OAI22_X1 U2531 ( .A1(n6008), .A2(n695), .B1(n14712), .B2(n696), .ZN(n12390)
         );
  OAI22_X1 U2532 ( .A1(n5992), .A2(n695), .B1(n14672), .B2(n696), .ZN(n12391)
         );
  OAI22_X1 U2533 ( .A1(n6748), .A2(n751), .B1(n14935), .B2(n752), .ZN(n12600)
         );
  OAI22_X1 U2534 ( .A1(n6732), .A2(n751), .B1(n14914), .B2(n752), .ZN(n12601)
         );
  OAI22_X1 U2535 ( .A1(n6716), .A2(n751), .B1(n14874), .B2(n752), .ZN(n12602)
         );
  OAI22_X1 U2536 ( .A1(n6700), .A2(n751), .B1(n14834), .B2(n752), .ZN(n12603)
         );
  OAI22_X1 U2537 ( .A1(n6684), .A2(n751), .B1(n14794), .B2(n752), .ZN(n12604)
         );
  OAI22_X1 U2538 ( .A1(n6668), .A2(n751), .B1(n14754), .B2(n752), .ZN(n12605)
         );
  OAI22_X1 U2539 ( .A1(n6652), .A2(n751), .B1(n14714), .B2(n752), .ZN(n12606)
         );
  OAI22_X1 U2540 ( .A1(n6636), .A2(n751), .B1(n14674), .B2(n752), .ZN(n12607)
         );
  OAI22_X1 U2541 ( .A1(n6620), .A2(n753), .B1(n14935), .B2(n754), .ZN(n12608)
         );
  OAI22_X1 U2542 ( .A1(n6604), .A2(n753), .B1(n14914), .B2(n754), .ZN(n12609)
         );
  OAI22_X1 U2543 ( .A1(n6588), .A2(n753), .B1(n14874), .B2(n754), .ZN(n12610)
         );
  OAI22_X1 U2544 ( .A1(n6572), .A2(n753), .B1(n14834), .B2(n754), .ZN(n12611)
         );
  OAI22_X1 U2545 ( .A1(n6556), .A2(n753), .B1(n14794), .B2(n754), .ZN(n12612)
         );
  OAI22_X1 U2546 ( .A1(n6540), .A2(n753), .B1(n14754), .B2(n754), .ZN(n12613)
         );
  OAI22_X1 U2547 ( .A1(n6524), .A2(n753), .B1(n14714), .B2(n754), .ZN(n12614)
         );
  OAI22_X1 U2548 ( .A1(n6508), .A2(n753), .B1(n14674), .B2(n754), .ZN(n12615)
         );
  OAI22_X1 U2549 ( .A1(n6492), .A2(n755), .B1(n14935), .B2(n756), .ZN(n12616)
         );
  OAI22_X1 U2550 ( .A1(n6476), .A2(n755), .B1(n14914), .B2(n756), .ZN(n12617)
         );
  OAI22_X1 U2551 ( .A1(n6460), .A2(n755), .B1(n14874), .B2(n756), .ZN(n12618)
         );
  OAI22_X1 U2552 ( .A1(n6444), .A2(n755), .B1(n14834), .B2(n756), .ZN(n12619)
         );
  OAI22_X1 U2553 ( .A1(n6428), .A2(n755), .B1(n14794), .B2(n756), .ZN(n12620)
         );
  OAI22_X1 U2554 ( .A1(n6412), .A2(n755), .B1(n14754), .B2(n756), .ZN(n12621)
         );
  OAI22_X1 U2555 ( .A1(n6396), .A2(n755), .B1(n14714), .B2(n756), .ZN(n12622)
         );
  OAI22_X1 U2556 ( .A1(n6380), .A2(n755), .B1(n14674), .B2(n756), .ZN(n12623)
         );
  OAI22_X1 U2557 ( .A1(n6364), .A2(n757), .B1(n14935), .B2(n758), .ZN(n12624)
         );
  OAI22_X1 U2558 ( .A1(n6348), .A2(n757), .B1(n14914), .B2(n758), .ZN(n12625)
         );
  OAI22_X1 U2559 ( .A1(n6332), .A2(n757), .B1(n14874), .B2(n758), .ZN(n12626)
         );
  OAI22_X1 U2560 ( .A1(n6316), .A2(n757), .B1(n14834), .B2(n758), .ZN(n12627)
         );
  OAI22_X1 U2561 ( .A1(n6300), .A2(n757), .B1(n14794), .B2(n758), .ZN(n12628)
         );
  OAI22_X1 U2562 ( .A1(n6284), .A2(n757), .B1(n14754), .B2(n758), .ZN(n12629)
         );
  OAI22_X1 U2563 ( .A1(n6268), .A2(n757), .B1(n14714), .B2(n758), .ZN(n12630)
         );
  OAI22_X1 U2564 ( .A1(n6252), .A2(n757), .B1(n14674), .B2(n758), .ZN(n12631)
         );
  OAI22_X1 U2565 ( .A1(n6236), .A2(n759), .B1(n14935), .B2(n760), .ZN(n12632)
         );
  OAI22_X1 U2566 ( .A1(n6220), .A2(n759), .B1(n14914), .B2(n760), .ZN(n12633)
         );
  OAI22_X1 U2567 ( .A1(n6204), .A2(n759), .B1(n14874), .B2(n760), .ZN(n12634)
         );
  OAI22_X1 U2568 ( .A1(n6188), .A2(n759), .B1(n14834), .B2(n760), .ZN(n12635)
         );
  OAI22_X1 U2569 ( .A1(n6172), .A2(n759), .B1(n14794), .B2(n760), .ZN(n12636)
         );
  OAI22_X1 U2570 ( .A1(n6156), .A2(n759), .B1(n14754), .B2(n760), .ZN(n12637)
         );
  OAI22_X1 U2571 ( .A1(n6140), .A2(n759), .B1(n14714), .B2(n760), .ZN(n12638)
         );
  OAI22_X1 U2572 ( .A1(n6124), .A2(n759), .B1(n14674), .B2(n760), .ZN(n12639)
         );
  OAI22_X1 U2573 ( .A1(n6108), .A2(n761), .B1(n14935), .B2(n762), .ZN(n12640)
         );
  OAI22_X1 U2574 ( .A1(n6092), .A2(n761), .B1(n14914), .B2(n762), .ZN(n12641)
         );
  OAI22_X1 U2575 ( .A1(n6076), .A2(n761), .B1(n14874), .B2(n762), .ZN(n12642)
         );
  OAI22_X1 U2576 ( .A1(n6060), .A2(n761), .B1(n14834), .B2(n762), .ZN(n12643)
         );
  OAI22_X1 U2577 ( .A1(n6044), .A2(n761), .B1(n14794), .B2(n762), .ZN(n12644)
         );
  OAI22_X1 U2578 ( .A1(n6028), .A2(n761), .B1(n14754), .B2(n762), .ZN(n12645)
         );
  OAI22_X1 U2579 ( .A1(n6012), .A2(n761), .B1(n14714), .B2(n762), .ZN(n12646)
         );
  OAI22_X1 U2580 ( .A1(n5996), .A2(n761), .B1(n14674), .B2(n762), .ZN(n12647)
         );
  OAI22_X1 U2581 ( .A1(n6752), .A2(n817), .B1(n14932), .B2(n818), .ZN(n12856)
         );
  OAI22_X1 U2582 ( .A1(n6736), .A2(n817), .B1(n14916), .B2(n818), .ZN(n12857)
         );
  OAI22_X1 U2583 ( .A1(n6720), .A2(n817), .B1(n14876), .B2(n818), .ZN(n12858)
         );
  OAI22_X1 U2584 ( .A1(n6704), .A2(n817), .B1(n14836), .B2(n818), .ZN(n12859)
         );
  OAI22_X1 U2585 ( .A1(n6688), .A2(n817), .B1(n14796), .B2(n818), .ZN(n12860)
         );
  OAI22_X1 U2586 ( .A1(n6672), .A2(n817), .B1(n14756), .B2(n818), .ZN(n12861)
         );
  OAI22_X1 U2587 ( .A1(n6656), .A2(n817), .B1(n14716), .B2(n818), .ZN(n12862)
         );
  OAI22_X1 U2588 ( .A1(n6640), .A2(n817), .B1(n14676), .B2(n818), .ZN(n12863)
         );
  OAI22_X1 U2589 ( .A1(n6624), .A2(n819), .B1(n14932), .B2(n820), .ZN(n12864)
         );
  OAI22_X1 U2590 ( .A1(n6608), .A2(n819), .B1(n14916), .B2(n820), .ZN(n12865)
         );
  OAI22_X1 U2591 ( .A1(n6592), .A2(n819), .B1(n14876), .B2(n820), .ZN(n12866)
         );
  OAI22_X1 U2592 ( .A1(n6576), .A2(n819), .B1(n14836), .B2(n820), .ZN(n12867)
         );
  OAI22_X1 U2593 ( .A1(n6560), .A2(n819), .B1(n14796), .B2(n820), .ZN(n12868)
         );
  OAI22_X1 U2594 ( .A1(n6544), .A2(n819), .B1(n14756), .B2(n820), .ZN(n12869)
         );
  OAI22_X1 U2595 ( .A1(n6528), .A2(n819), .B1(n14716), .B2(n820), .ZN(n12870)
         );
  OAI22_X1 U2596 ( .A1(n6512), .A2(n819), .B1(n14676), .B2(n820), .ZN(n12871)
         );
  OAI22_X1 U2597 ( .A1(n6496), .A2(n821), .B1(n14932), .B2(n822), .ZN(n12872)
         );
  OAI22_X1 U2598 ( .A1(n6480), .A2(n821), .B1(n14916), .B2(n822), .ZN(n12873)
         );
  OAI22_X1 U2599 ( .A1(n6464), .A2(n821), .B1(n14876), .B2(n822), .ZN(n12874)
         );
  OAI22_X1 U2600 ( .A1(n6448), .A2(n821), .B1(n14836), .B2(n822), .ZN(n12875)
         );
  OAI22_X1 U2601 ( .A1(n6432), .A2(n821), .B1(n14796), .B2(n822), .ZN(n12876)
         );
  OAI22_X1 U2602 ( .A1(n6416), .A2(n821), .B1(n14756), .B2(n822), .ZN(n12877)
         );
  OAI22_X1 U2603 ( .A1(n6400), .A2(n821), .B1(n14716), .B2(n822), .ZN(n12878)
         );
  OAI22_X1 U2604 ( .A1(n6384), .A2(n821), .B1(n14676), .B2(n822), .ZN(n12879)
         );
  OAI22_X1 U2605 ( .A1(n6368), .A2(n823), .B1(n14932), .B2(n824), .ZN(n12880)
         );
  OAI22_X1 U2606 ( .A1(n6352), .A2(n823), .B1(n14916), .B2(n824), .ZN(n12881)
         );
  OAI22_X1 U2607 ( .A1(n6336), .A2(n823), .B1(n14876), .B2(n824), .ZN(n12882)
         );
  OAI22_X1 U2608 ( .A1(n6320), .A2(n823), .B1(n14836), .B2(n824), .ZN(n12883)
         );
  OAI22_X1 U2609 ( .A1(n6304), .A2(n823), .B1(n14796), .B2(n824), .ZN(n12884)
         );
  OAI22_X1 U2610 ( .A1(n6288), .A2(n823), .B1(n14756), .B2(n824), .ZN(n12885)
         );
  OAI22_X1 U2611 ( .A1(n6272), .A2(n823), .B1(n14716), .B2(n824), .ZN(n12886)
         );
  OAI22_X1 U2612 ( .A1(n6256), .A2(n823), .B1(n14676), .B2(n824), .ZN(n12887)
         );
  OAI22_X1 U2613 ( .A1(n6240), .A2(n825), .B1(n14932), .B2(n826), .ZN(n12888)
         );
  OAI22_X1 U2614 ( .A1(n6224), .A2(n825), .B1(n14916), .B2(n826), .ZN(n12889)
         );
  OAI22_X1 U2615 ( .A1(n6208), .A2(n825), .B1(n14876), .B2(n826), .ZN(n12890)
         );
  OAI22_X1 U2616 ( .A1(n6192), .A2(n825), .B1(n14836), .B2(n826), .ZN(n12891)
         );
  OAI22_X1 U2617 ( .A1(n6176), .A2(n825), .B1(n14796), .B2(n826), .ZN(n12892)
         );
  OAI22_X1 U2618 ( .A1(n6160), .A2(n825), .B1(n14756), .B2(n826), .ZN(n12893)
         );
  OAI22_X1 U2619 ( .A1(n6144), .A2(n825), .B1(n14716), .B2(n826), .ZN(n12894)
         );
  OAI22_X1 U2620 ( .A1(n6128), .A2(n825), .B1(n14676), .B2(n826), .ZN(n12895)
         );
  OAI22_X1 U2621 ( .A1(n6112), .A2(n827), .B1(n14932), .B2(n828), .ZN(n12896)
         );
  OAI22_X1 U2622 ( .A1(n6096), .A2(n827), .B1(n14917), .B2(n828), .ZN(n12897)
         );
  OAI22_X1 U2623 ( .A1(n6080), .A2(n827), .B1(n14877), .B2(n828), .ZN(n12898)
         );
  OAI22_X1 U2624 ( .A1(n6064), .A2(n827), .B1(n14837), .B2(n828), .ZN(n12899)
         );
  OAI22_X1 U2625 ( .A1(n6048), .A2(n827), .B1(n14797), .B2(n828), .ZN(n12900)
         );
  OAI22_X1 U2626 ( .A1(n6032), .A2(n827), .B1(n14757), .B2(n828), .ZN(n12901)
         );
  OAI22_X1 U2627 ( .A1(n6016), .A2(n827), .B1(n14717), .B2(n828), .ZN(n12902)
         );
  OAI22_X1 U2628 ( .A1(n6000), .A2(n827), .B1(n14677), .B2(n828), .ZN(n12903)
         );
  OAI22_X1 U2629 ( .A1(n6756), .A2(n882), .B1(n14930), .B2(n883), .ZN(n13112)
         );
  OAI22_X1 U2630 ( .A1(n6740), .A2(n882), .B1(n14919), .B2(n883), .ZN(n13113)
         );
  OAI22_X1 U2631 ( .A1(n6724), .A2(n882), .B1(n14879), .B2(n883), .ZN(n13114)
         );
  OAI22_X1 U2632 ( .A1(n6708), .A2(n882), .B1(n14839), .B2(n883), .ZN(n13115)
         );
  OAI22_X1 U2633 ( .A1(n6692), .A2(n882), .B1(n14799), .B2(n883), .ZN(n13116)
         );
  OAI22_X1 U2634 ( .A1(n6676), .A2(n882), .B1(n14759), .B2(n883), .ZN(n13117)
         );
  OAI22_X1 U2635 ( .A1(n6660), .A2(n882), .B1(n14719), .B2(n883), .ZN(n13118)
         );
  OAI22_X1 U2636 ( .A1(n6644), .A2(n882), .B1(n14679), .B2(n883), .ZN(n13119)
         );
  OAI22_X1 U2637 ( .A1(n6628), .A2(n884), .B1(n14930), .B2(n885), .ZN(n13120)
         );
  OAI22_X1 U2638 ( .A1(n6612), .A2(n884), .B1(n14919), .B2(n885), .ZN(n13121)
         );
  OAI22_X1 U2639 ( .A1(n6596), .A2(n884), .B1(n14879), .B2(n885), .ZN(n13122)
         );
  OAI22_X1 U2640 ( .A1(n6580), .A2(n884), .B1(n14839), .B2(n885), .ZN(n13123)
         );
  OAI22_X1 U2641 ( .A1(n6564), .A2(n884), .B1(n14799), .B2(n885), .ZN(n13124)
         );
  OAI22_X1 U2642 ( .A1(n6548), .A2(n884), .B1(n14759), .B2(n885), .ZN(n13125)
         );
  OAI22_X1 U2643 ( .A1(n6532), .A2(n884), .B1(n14719), .B2(n885), .ZN(n13126)
         );
  OAI22_X1 U2644 ( .A1(n6516), .A2(n884), .B1(n14679), .B2(n885), .ZN(n13127)
         );
  OAI22_X1 U2645 ( .A1(n6500), .A2(n886), .B1(n14930), .B2(n887), .ZN(n13128)
         );
  OAI22_X1 U2646 ( .A1(n6484), .A2(n886), .B1(n14919), .B2(n887), .ZN(n13129)
         );
  OAI22_X1 U2647 ( .A1(n6468), .A2(n886), .B1(n14879), .B2(n887), .ZN(n13130)
         );
  OAI22_X1 U2648 ( .A1(n6452), .A2(n886), .B1(n14839), .B2(n887), .ZN(n13131)
         );
  OAI22_X1 U2649 ( .A1(n6436), .A2(n886), .B1(n14799), .B2(n887), .ZN(n13132)
         );
  OAI22_X1 U2650 ( .A1(n6420), .A2(n886), .B1(n14759), .B2(n887), .ZN(n13133)
         );
  OAI22_X1 U2651 ( .A1(n6404), .A2(n886), .B1(n14719), .B2(n887), .ZN(n13134)
         );
  OAI22_X1 U2652 ( .A1(n6388), .A2(n886), .B1(n14679), .B2(n887), .ZN(n13135)
         );
  OAI22_X1 U2653 ( .A1(n6372), .A2(n888), .B1(n14930), .B2(n889), .ZN(n13136)
         );
  OAI22_X1 U2654 ( .A1(n6356), .A2(n888), .B1(n14919), .B2(n889), .ZN(n13137)
         );
  OAI22_X1 U2655 ( .A1(n6340), .A2(n888), .B1(n14879), .B2(n889), .ZN(n13138)
         );
  OAI22_X1 U2656 ( .A1(n6324), .A2(n888), .B1(n14839), .B2(n889), .ZN(n13139)
         );
  OAI22_X1 U2657 ( .A1(n6308), .A2(n888), .B1(n14799), .B2(n889), .ZN(n13140)
         );
  OAI22_X1 U2658 ( .A1(n6292), .A2(n888), .B1(n14759), .B2(n889), .ZN(n13141)
         );
  OAI22_X1 U2659 ( .A1(n6276), .A2(n888), .B1(n14719), .B2(n889), .ZN(n13142)
         );
  OAI22_X1 U2660 ( .A1(n6260), .A2(n888), .B1(n14679), .B2(n889), .ZN(n13143)
         );
  OAI22_X1 U2661 ( .A1(n6244), .A2(n890), .B1(n14930), .B2(n891), .ZN(n13144)
         );
  OAI22_X1 U2662 ( .A1(n6228), .A2(n890), .B1(n14919), .B2(n891), .ZN(n13145)
         );
  OAI22_X1 U2663 ( .A1(n6212), .A2(n890), .B1(n14879), .B2(n891), .ZN(n13146)
         );
  OAI22_X1 U2664 ( .A1(n6196), .A2(n890), .B1(n14839), .B2(n891), .ZN(n13147)
         );
  OAI22_X1 U2665 ( .A1(n6180), .A2(n890), .B1(n14799), .B2(n891), .ZN(n13148)
         );
  OAI22_X1 U2666 ( .A1(n6164), .A2(n890), .B1(n14759), .B2(n891), .ZN(n13149)
         );
  OAI22_X1 U2667 ( .A1(n6148), .A2(n890), .B1(n14719), .B2(n891), .ZN(n13150)
         );
  OAI22_X1 U2668 ( .A1(n6132), .A2(n890), .B1(n14679), .B2(n891), .ZN(n13151)
         );
  OAI22_X1 U2669 ( .A1(n6116), .A2(n892), .B1(n14934), .B2(n893), .ZN(n13152)
         );
  OAI22_X1 U2670 ( .A1(n6100), .A2(n892), .B1(n14919), .B2(n893), .ZN(n13153)
         );
  OAI22_X1 U2671 ( .A1(n6084), .A2(n892), .B1(n14879), .B2(n893), .ZN(n13154)
         );
  OAI22_X1 U2672 ( .A1(n6068), .A2(n892), .B1(n14839), .B2(n893), .ZN(n13155)
         );
  OAI22_X1 U2673 ( .A1(n6052), .A2(n892), .B1(n14799), .B2(n893), .ZN(n13156)
         );
  OAI22_X1 U2674 ( .A1(n6036), .A2(n892), .B1(n14759), .B2(n893), .ZN(n13157)
         );
  OAI22_X1 U2675 ( .A1(n6020), .A2(n892), .B1(n14719), .B2(n893), .ZN(n13158)
         );
  OAI22_X1 U2676 ( .A1(n6004), .A2(n892), .B1(n14679), .B2(n893), .ZN(n13159)
         );
  OAI22_X1 U2677 ( .A1(n6750), .A2(n1013), .B1(n14945), .B2(n1014), .ZN(n13624) );
  OAI22_X1 U2678 ( .A1(n6734), .A2(n1013), .B1(n14924), .B2(n1014), .ZN(n13625) );
  OAI22_X1 U2679 ( .A1(n6718), .A2(n1013), .B1(n14884), .B2(n1014), .ZN(n13626) );
  OAI22_X1 U2680 ( .A1(n6702), .A2(n1013), .B1(n14844), .B2(n1014), .ZN(n13627) );
  OAI22_X1 U2681 ( .A1(n6686), .A2(n1013), .B1(n14804), .B2(n1014), .ZN(n13628) );
  OAI22_X1 U2682 ( .A1(n6670), .A2(n1013), .B1(n14764), .B2(n1014), .ZN(n13629) );
  OAI22_X1 U2683 ( .A1(n6654), .A2(n1013), .B1(n14724), .B2(n1014), .ZN(n13630) );
  OAI22_X1 U2684 ( .A1(n6638), .A2(n1013), .B1(n14684), .B2(n1014), .ZN(n13631) );
  OAI22_X1 U2685 ( .A1(n6622), .A2(n1015), .B1(n14945), .B2(n1016), .ZN(n13632) );
  OAI22_X1 U2686 ( .A1(n6606), .A2(n1015), .B1(n14924), .B2(n1016), .ZN(n13633) );
  OAI22_X1 U2687 ( .A1(n6590), .A2(n1015), .B1(n14884), .B2(n1016), .ZN(n13634) );
  OAI22_X1 U2688 ( .A1(n6574), .A2(n1015), .B1(n14844), .B2(n1016), .ZN(n13635) );
  OAI22_X1 U2689 ( .A1(n6558), .A2(n1015), .B1(n14804), .B2(n1016), .ZN(n13636) );
  OAI22_X1 U2690 ( .A1(n6542), .A2(n1015), .B1(n14764), .B2(n1016), .ZN(n13637) );
  OAI22_X1 U2691 ( .A1(n6526), .A2(n1015), .B1(n14724), .B2(n1016), .ZN(n13638) );
  OAI22_X1 U2692 ( .A1(n6510), .A2(n1015), .B1(n14684), .B2(n1016), .ZN(n13639) );
  OAI22_X1 U2693 ( .A1(n6494), .A2(n1017), .B1(n14945), .B2(n1018), .ZN(n13640) );
  OAI22_X1 U2694 ( .A1(n6478), .A2(n1017), .B1(n14924), .B2(n1018), .ZN(n13641) );
  OAI22_X1 U2695 ( .A1(n6462), .A2(n1017), .B1(n14884), .B2(n1018), .ZN(n13642) );
  OAI22_X1 U2696 ( .A1(n6446), .A2(n1017), .B1(n14844), .B2(n1018), .ZN(n13643) );
  OAI22_X1 U2697 ( .A1(n6430), .A2(n1017), .B1(n14804), .B2(n1018), .ZN(n13644) );
  OAI22_X1 U2698 ( .A1(n6414), .A2(n1017), .B1(n14764), .B2(n1018), .ZN(n13645) );
  OAI22_X1 U2699 ( .A1(n6398), .A2(n1017), .B1(n14724), .B2(n1018), .ZN(n13646) );
  OAI22_X1 U2700 ( .A1(n6382), .A2(n1017), .B1(n14684), .B2(n1018), .ZN(n13647) );
  OAI22_X1 U2701 ( .A1(n6366), .A2(n1019), .B1(n14944), .B2(n1020), .ZN(n13648) );
  OAI22_X1 U2702 ( .A1(n6350), .A2(n1019), .B1(n14924), .B2(n1020), .ZN(n13649) );
  OAI22_X1 U2703 ( .A1(n6334), .A2(n1019), .B1(n14884), .B2(n1020), .ZN(n13650) );
  OAI22_X1 U2704 ( .A1(n6318), .A2(n1019), .B1(n14844), .B2(n1020), .ZN(n13651) );
  OAI22_X1 U2705 ( .A1(n6302), .A2(n1019), .B1(n14804), .B2(n1020), .ZN(n13652) );
  OAI22_X1 U2706 ( .A1(n6286), .A2(n1019), .B1(n14764), .B2(n1020), .ZN(n13653) );
  OAI22_X1 U2707 ( .A1(n6270), .A2(n1019), .B1(n14724), .B2(n1020), .ZN(n13654) );
  OAI22_X1 U2708 ( .A1(n6254), .A2(n1019), .B1(n14684), .B2(n1020), .ZN(n13655) );
  OAI22_X1 U2709 ( .A1(n6238), .A2(n1021), .B1(n14944), .B2(n1022), .ZN(n13656) );
  OAI22_X1 U2710 ( .A1(n6222), .A2(n1021), .B1(n14924), .B2(n1022), .ZN(n13657) );
  OAI22_X1 U2711 ( .A1(n6206), .A2(n1021), .B1(n14884), .B2(n1022), .ZN(n13658) );
  OAI22_X1 U2712 ( .A1(n6190), .A2(n1021), .B1(n14844), .B2(n1022), .ZN(n13659) );
  OAI22_X1 U2713 ( .A1(n6174), .A2(n1021), .B1(n14804), .B2(n1022), .ZN(n13660) );
  OAI22_X1 U2714 ( .A1(n6158), .A2(n1021), .B1(n14764), .B2(n1022), .ZN(n13661) );
  OAI22_X1 U2715 ( .A1(n6142), .A2(n1021), .B1(n14724), .B2(n1022), .ZN(n13662) );
  OAI22_X1 U2716 ( .A1(n6126), .A2(n1021), .B1(n14684), .B2(n1022), .ZN(n13663) );
  OAI22_X1 U2717 ( .A1(n6110), .A2(n1023), .B1(n14944), .B2(n1024), .ZN(n13664) );
  OAI22_X1 U2718 ( .A1(n6094), .A2(n1023), .B1(n14924), .B2(n1024), .ZN(n13665) );
  OAI22_X1 U2719 ( .A1(n6078), .A2(n1023), .B1(n14884), .B2(n1024), .ZN(n13666) );
  OAI22_X1 U2720 ( .A1(n6062), .A2(n1023), .B1(n14844), .B2(n1024), .ZN(n13667) );
  OAI22_X1 U2721 ( .A1(n6046), .A2(n1023), .B1(n14804), .B2(n1024), .ZN(n13668) );
  OAI22_X1 U2722 ( .A1(n6030), .A2(n1023), .B1(n14764), .B2(n1024), .ZN(n13669) );
  OAI22_X1 U2723 ( .A1(n6014), .A2(n1023), .B1(n14724), .B2(n1024), .ZN(n13670) );
  OAI22_X1 U2724 ( .A1(n5998), .A2(n1023), .B1(n14684), .B2(n1024), .ZN(n13671) );
  OAI22_X1 U2725 ( .A1(n6758), .A2(n1155), .B1(n14940), .B2(n1156), .ZN(n14136) );
  OAI22_X1 U2726 ( .A1(n6742), .A2(n1155), .B1(n14928), .B2(n1156), .ZN(n14137) );
  OAI22_X1 U2727 ( .A1(n6726), .A2(n1155), .B1(n14888), .B2(n1156), .ZN(n14138) );
  OAI22_X1 U2728 ( .A1(n6710), .A2(n1155), .B1(n14848), .B2(n1156), .ZN(n14139) );
  OAI22_X1 U2729 ( .A1(n6694), .A2(n1155), .B1(n14808), .B2(n1156), .ZN(n14140) );
  OAI22_X1 U2730 ( .A1(n6678), .A2(n1155), .B1(n14768), .B2(n1156), .ZN(n14141) );
  OAI22_X1 U2731 ( .A1(n6662), .A2(n1155), .B1(n14728), .B2(n1156), .ZN(n14142) );
  OAI22_X1 U2732 ( .A1(n6646), .A2(n1155), .B1(n14688), .B2(n1156), .ZN(n14143) );
  OAI22_X1 U2733 ( .A1(n6630), .A2(n1157), .B1(n14940), .B2(n1158), .ZN(n14144) );
  OAI22_X1 U2734 ( .A1(n6502), .A2(n1159), .B1(n14940), .B2(n1160), .ZN(n14152) );
  OAI22_X1 U2735 ( .A1(n6374), .A2(n1162), .B1(n14939), .B2(n1163), .ZN(n14160) );
  OAI22_X1 U2736 ( .A1(n6246), .A2(n1165), .B1(n14944), .B2(n1166), .ZN(n14168) );
  OAI22_X1 U2737 ( .A1(n6118), .A2(n1167), .B1(n14949), .B2(n1168), .ZN(n14176) );
  OAI22_X1 U2738 ( .A1(n10079), .A2(n436), .B1(n14966), .B2(n437), .ZN(n11368)
         );
  OAI22_X1 U2739 ( .A1(n10063), .A2(n436), .B1(n14902), .B2(n437), .ZN(n11369)
         );
  OAI22_X1 U2740 ( .A1(n10047), .A2(n436), .B1(n14862), .B2(n437), .ZN(n11370)
         );
  OAI22_X1 U2741 ( .A1(n10031), .A2(n436), .B1(n14822), .B2(n437), .ZN(n11371)
         );
  OAI22_X1 U2742 ( .A1(n10015), .A2(n436), .B1(n14782), .B2(n437), .ZN(n11372)
         );
  OAI22_X1 U2743 ( .A1(n9999), .A2(n436), .B1(n14742), .B2(n437), .ZN(n11373)
         );
  OAI22_X1 U2744 ( .A1(n9983), .A2(n436), .B1(n14702), .B2(n437), .ZN(n11374)
         );
  OAI22_X1 U2745 ( .A1(n9967), .A2(n436), .B1(n14662), .B2(n437), .ZN(n11375)
         );
  OAI22_X1 U2746 ( .A1(n9951), .A2(n439), .B1(n14966), .B2(n440), .ZN(n11376)
         );
  OAI22_X1 U2747 ( .A1(n9935), .A2(n439), .B1(n14902), .B2(n440), .ZN(n11377)
         );
  OAI22_X1 U2748 ( .A1(n9919), .A2(n439), .B1(n14862), .B2(n440), .ZN(n11378)
         );
  OAI22_X1 U2749 ( .A1(n9903), .A2(n439), .B1(n14822), .B2(n440), .ZN(n11379)
         );
  OAI22_X1 U2750 ( .A1(n9887), .A2(n439), .B1(n14782), .B2(n440), .ZN(n11380)
         );
  OAI22_X1 U2751 ( .A1(n9871), .A2(n439), .B1(n14742), .B2(n440), .ZN(n11381)
         );
  OAI22_X1 U2752 ( .A1(n9855), .A2(n439), .B1(n14702), .B2(n440), .ZN(n11382)
         );
  OAI22_X1 U2753 ( .A1(n9839), .A2(n439), .B1(n14662), .B2(n440), .ZN(n11383)
         );
  OAI22_X1 U2754 ( .A1(n9823), .A2(n441), .B1(n14966), .B2(n442), .ZN(n11384)
         );
  OAI22_X1 U2755 ( .A1(n9807), .A2(n441), .B1(n14902), .B2(n442), .ZN(n11385)
         );
  OAI22_X1 U2756 ( .A1(n9791), .A2(n441), .B1(n14862), .B2(n442), .ZN(n11386)
         );
  OAI22_X1 U2757 ( .A1(n9775), .A2(n441), .B1(n14822), .B2(n442), .ZN(n11387)
         );
  OAI22_X1 U2758 ( .A1(n9759), .A2(n441), .B1(n14782), .B2(n442), .ZN(n11388)
         );
  OAI22_X1 U2759 ( .A1(n9743), .A2(n441), .B1(n14742), .B2(n442), .ZN(n11389)
         );
  OAI22_X1 U2760 ( .A1(n9727), .A2(n441), .B1(n14702), .B2(n442), .ZN(n11390)
         );
  OAI22_X1 U2761 ( .A1(n9711), .A2(n441), .B1(n14662), .B2(n442), .ZN(n11391)
         );
  OAI22_X1 U2762 ( .A1(n9695), .A2(n443), .B1(n14966), .B2(n444), .ZN(n11392)
         );
  OAI22_X1 U2763 ( .A1(n9679), .A2(n443), .B1(n14902), .B2(n444), .ZN(n11393)
         );
  OAI22_X1 U2764 ( .A1(n9663), .A2(n443), .B1(n14862), .B2(n444), .ZN(n11394)
         );
  OAI22_X1 U2765 ( .A1(n9647), .A2(n443), .B1(n14822), .B2(n444), .ZN(n11395)
         );
  OAI22_X1 U2766 ( .A1(n9631), .A2(n443), .B1(n14782), .B2(n444), .ZN(n11396)
         );
  OAI22_X1 U2767 ( .A1(n9615), .A2(n443), .B1(n14742), .B2(n444), .ZN(n11397)
         );
  OAI22_X1 U2768 ( .A1(n9599), .A2(n443), .B1(n14702), .B2(n444), .ZN(n11398)
         );
  OAI22_X1 U2769 ( .A1(n9583), .A2(n443), .B1(n14662), .B2(n444), .ZN(n11399)
         );
  OAI22_X1 U2770 ( .A1(n9567), .A2(n445), .B1(n14966), .B2(n446), .ZN(n11400)
         );
  OAI22_X1 U2771 ( .A1(n9551), .A2(n445), .B1(n14902), .B2(n446), .ZN(n11401)
         );
  OAI22_X1 U2772 ( .A1(n9535), .A2(n445), .B1(n14862), .B2(n446), .ZN(n11402)
         );
  OAI22_X1 U2773 ( .A1(n9519), .A2(n445), .B1(n14822), .B2(n446), .ZN(n11403)
         );
  OAI22_X1 U2774 ( .A1(n9503), .A2(n445), .B1(n14782), .B2(n446), .ZN(n11404)
         );
  OAI22_X1 U2775 ( .A1(n9487), .A2(n445), .B1(n14742), .B2(n446), .ZN(n11405)
         );
  OAI22_X1 U2776 ( .A1(n9471), .A2(n445), .B1(n14702), .B2(n446), .ZN(n11406)
         );
  OAI22_X1 U2777 ( .A1(n9455), .A2(n445), .B1(n14662), .B2(n446), .ZN(n11407)
         );
  OAI22_X1 U2778 ( .A1(n9439), .A2(n447), .B1(n14966), .B2(n448), .ZN(n11408)
         );
  OAI22_X1 U2779 ( .A1(n9423), .A2(n447), .B1(n14902), .B2(n448), .ZN(n11409)
         );
  OAI22_X1 U2780 ( .A1(n9407), .A2(n447), .B1(n14862), .B2(n448), .ZN(n11410)
         );
  OAI22_X1 U2781 ( .A1(n9391), .A2(n447), .B1(n14822), .B2(n448), .ZN(n11411)
         );
  OAI22_X1 U2782 ( .A1(n9375), .A2(n447), .B1(n14782), .B2(n448), .ZN(n11412)
         );
  OAI22_X1 U2783 ( .A1(n9359), .A2(n447), .B1(n14742), .B2(n448), .ZN(n11413)
         );
  OAI22_X1 U2784 ( .A1(n9343), .A2(n447), .B1(n14702), .B2(n448), .ZN(n11414)
         );
  OAI22_X1 U2785 ( .A1(n9327), .A2(n447), .B1(n14662), .B2(n448), .ZN(n11415)
         );
  OAI22_X1 U2786 ( .A1(n10074), .A2(n894), .B1(n14949), .B2(n895), .ZN(n13160)
         );
  OAI22_X1 U2787 ( .A1(n10058), .A2(n894), .B1(n14919), .B2(n895), .ZN(n13161)
         );
  OAI22_X1 U2788 ( .A1(n10042), .A2(n894), .B1(n14879), .B2(n895), .ZN(n13162)
         );
  OAI22_X1 U2789 ( .A1(n10026), .A2(n894), .B1(n14839), .B2(n895), .ZN(n13163)
         );
  OAI22_X1 U2790 ( .A1(n10010), .A2(n894), .B1(n14799), .B2(n895), .ZN(n13164)
         );
  OAI22_X1 U2791 ( .A1(n9994), .A2(n894), .B1(n14759), .B2(n895), .ZN(n13165)
         );
  OAI22_X1 U2792 ( .A1(n9978), .A2(n894), .B1(n14719), .B2(n895), .ZN(n13166)
         );
  OAI22_X1 U2793 ( .A1(n9962), .A2(n894), .B1(n14679), .B2(n895), .ZN(n13167)
         );
  OAI22_X1 U2794 ( .A1(n9946), .A2(n897), .B1(n14949), .B2(n898), .ZN(n13168)
         );
  OAI22_X1 U2795 ( .A1(n9930), .A2(n897), .B1(n14919), .B2(n898), .ZN(n13169)
         );
  OAI22_X1 U2796 ( .A1(n9914), .A2(n897), .B1(n14879), .B2(n898), .ZN(n13170)
         );
  OAI22_X1 U2797 ( .A1(n9898), .A2(n897), .B1(n14839), .B2(n898), .ZN(n13171)
         );
  OAI22_X1 U2798 ( .A1(n9882), .A2(n897), .B1(n14799), .B2(n898), .ZN(n13172)
         );
  OAI22_X1 U2799 ( .A1(n9866), .A2(n897), .B1(n14759), .B2(n898), .ZN(n13173)
         );
  OAI22_X1 U2800 ( .A1(n9850), .A2(n897), .B1(n14719), .B2(n898), .ZN(n13174)
         );
  OAI22_X1 U2801 ( .A1(n9834), .A2(n897), .B1(n14679), .B2(n898), .ZN(n13175)
         );
  OAI22_X1 U2802 ( .A1(n9818), .A2(n899), .B1(n14949), .B2(n900), .ZN(n13176)
         );
  OAI22_X1 U2803 ( .A1(n9802), .A2(n899), .B1(n14919), .B2(n900), .ZN(n13177)
         );
  OAI22_X1 U2804 ( .A1(n9786), .A2(n899), .B1(n14879), .B2(n900), .ZN(n13178)
         );
  OAI22_X1 U2805 ( .A1(n9770), .A2(n899), .B1(n14839), .B2(n900), .ZN(n13179)
         );
  OAI22_X1 U2806 ( .A1(n9754), .A2(n899), .B1(n14799), .B2(n900), .ZN(n13180)
         );
  OAI22_X1 U2807 ( .A1(n9738), .A2(n899), .B1(n14759), .B2(n900), .ZN(n13181)
         );
  OAI22_X1 U2808 ( .A1(n9722), .A2(n899), .B1(n14719), .B2(n900), .ZN(n13182)
         );
  OAI22_X1 U2809 ( .A1(n9706), .A2(n899), .B1(n14679), .B2(n900), .ZN(n13183)
         );
  OAI22_X1 U2810 ( .A1(n9690), .A2(n901), .B1(n14949), .B2(n902), .ZN(n13184)
         );
  OAI22_X1 U2811 ( .A1(n9674), .A2(n901), .B1(n14919), .B2(n902), .ZN(n13185)
         );
  OAI22_X1 U2812 ( .A1(n9658), .A2(n901), .B1(n14879), .B2(n902), .ZN(n13186)
         );
  OAI22_X1 U2813 ( .A1(n9642), .A2(n901), .B1(n14839), .B2(n902), .ZN(n13187)
         );
  OAI22_X1 U2814 ( .A1(n9626), .A2(n901), .B1(n14799), .B2(n902), .ZN(n13188)
         );
  OAI22_X1 U2815 ( .A1(n9610), .A2(n901), .B1(n14759), .B2(n902), .ZN(n13189)
         );
  OAI22_X1 U2816 ( .A1(n9594), .A2(n901), .B1(n14719), .B2(n902), .ZN(n13190)
         );
  OAI22_X1 U2817 ( .A1(n9578), .A2(n901), .B1(n14679), .B2(n902), .ZN(n13191)
         );
  OAI22_X1 U2818 ( .A1(n9562), .A2(n903), .B1(n14949), .B2(n904), .ZN(n13192)
         );
  OAI22_X1 U2819 ( .A1(n9546), .A2(n903), .B1(n14919), .B2(n904), .ZN(n13193)
         );
  OAI22_X1 U2820 ( .A1(n9530), .A2(n903), .B1(n14879), .B2(n904), .ZN(n13194)
         );
  OAI22_X1 U2821 ( .A1(n9514), .A2(n903), .B1(n14839), .B2(n904), .ZN(n13195)
         );
  OAI22_X1 U2822 ( .A1(n9498), .A2(n903), .B1(n14799), .B2(n904), .ZN(n13196)
         );
  OAI22_X1 U2823 ( .A1(n9482), .A2(n903), .B1(n14759), .B2(n904), .ZN(n13197)
         );
  OAI22_X1 U2824 ( .A1(n9466), .A2(n903), .B1(n14719), .B2(n904), .ZN(n13198)
         );
  OAI22_X1 U2825 ( .A1(n9450), .A2(n903), .B1(n14679), .B2(n904), .ZN(n13199)
         );
  OAI22_X1 U2826 ( .A1(n9434), .A2(n905), .B1(n14949), .B2(n906), .ZN(n13200)
         );
  OAI22_X1 U2827 ( .A1(n9418), .A2(n905), .B1(n14919), .B2(n906), .ZN(n13201)
         );
  OAI22_X1 U2828 ( .A1(n9402), .A2(n905), .B1(n14879), .B2(n906), .ZN(n13202)
         );
  OAI22_X1 U2829 ( .A1(n9386), .A2(n905), .B1(n14839), .B2(n906), .ZN(n13203)
         );
  OAI22_X1 U2830 ( .A1(n9370), .A2(n905), .B1(n14799), .B2(n906), .ZN(n13204)
         );
  OAI22_X1 U2831 ( .A1(n9354), .A2(n905), .B1(n14759), .B2(n906), .ZN(n13205)
         );
  OAI22_X1 U2832 ( .A1(n9338), .A2(n905), .B1(n14719), .B2(n906), .ZN(n13206)
         );
  OAI22_X1 U2833 ( .A1(n9322), .A2(n905), .B1(n14679), .B2(n906), .ZN(n13207)
         );
  OAI22_X1 U2834 ( .A1(n10073), .A2(n66), .B1(n67), .B2(n14930), .ZN(n10088)
         );
  OAI22_X1 U2835 ( .A1(n9313), .A2(n253), .B1(n14954), .B2(n254), .ZN(n10648)
         );
  OAI22_X1 U2836 ( .A1(n9297), .A2(n253), .B1(n14895), .B2(n254), .ZN(n10649)
         );
  OAI22_X1 U2837 ( .A1(n9281), .A2(n253), .B1(n14855), .B2(n254), .ZN(n10650)
         );
  OAI22_X1 U2838 ( .A1(n9265), .A2(n253), .B1(n14815), .B2(n254), .ZN(n10651)
         );
  OAI22_X1 U2839 ( .A1(n9249), .A2(n253), .B1(n14775), .B2(n254), .ZN(n10652)
         );
  OAI22_X1 U2840 ( .A1(n9233), .A2(n253), .B1(n14735), .B2(n254), .ZN(n10653)
         );
  OAI22_X1 U2841 ( .A1(n9217), .A2(n253), .B1(n14695), .B2(n254), .ZN(n10654)
         );
  OAI22_X1 U2842 ( .A1(n9201), .A2(n253), .B1(n14655), .B2(n254), .ZN(n10655)
         );
  OAI22_X1 U2843 ( .A1(n9185), .A2(n255), .B1(n14954), .B2(n256), .ZN(n10656)
         );
  OAI22_X1 U2844 ( .A1(n9169), .A2(n255), .B1(n14895), .B2(n256), .ZN(n10657)
         );
  OAI22_X1 U2845 ( .A1(n9153), .A2(n255), .B1(n14855), .B2(n256), .ZN(n10658)
         );
  OAI22_X1 U2846 ( .A1(n9137), .A2(n255), .B1(n14815), .B2(n256), .ZN(n10659)
         );
  OAI22_X1 U2847 ( .A1(n9121), .A2(n255), .B1(n14775), .B2(n256), .ZN(n10660)
         );
  OAI22_X1 U2848 ( .A1(n9105), .A2(n255), .B1(n14735), .B2(n256), .ZN(n10661)
         );
  OAI22_X1 U2849 ( .A1(n9089), .A2(n255), .B1(n14695), .B2(n256), .ZN(n10662)
         );
  OAI22_X1 U2850 ( .A1(n9073), .A2(n255), .B1(n14655), .B2(n256), .ZN(n10663)
         );
  OAI22_X1 U2851 ( .A1(n9057), .A2(n257), .B1(n14953), .B2(n258), .ZN(n10664)
         );
  OAI22_X1 U2852 ( .A1(n9041), .A2(n257), .B1(n14895), .B2(n258), .ZN(n10665)
         );
  OAI22_X1 U2853 ( .A1(n9025), .A2(n257), .B1(n14855), .B2(n258), .ZN(n10666)
         );
  OAI22_X1 U2854 ( .A1(n9009), .A2(n257), .B1(n14815), .B2(n258), .ZN(n10667)
         );
  OAI22_X1 U2855 ( .A1(n8993), .A2(n257), .B1(n14775), .B2(n258), .ZN(n10668)
         );
  OAI22_X1 U2856 ( .A1(n8977), .A2(n257), .B1(n14735), .B2(n258), .ZN(n10669)
         );
  OAI22_X1 U2857 ( .A1(n8961), .A2(n257), .B1(n14695), .B2(n258), .ZN(n10670)
         );
  OAI22_X1 U2858 ( .A1(n8945), .A2(n257), .B1(n14655), .B2(n258), .ZN(n10671)
         );
  OAI22_X1 U2859 ( .A1(n8929), .A2(n259), .B1(n14953), .B2(n260), .ZN(n10672)
         );
  OAI22_X1 U2860 ( .A1(n8913), .A2(n259), .B1(n14895), .B2(n260), .ZN(n10673)
         );
  OAI22_X1 U2861 ( .A1(n8897), .A2(n259), .B1(n14855), .B2(n260), .ZN(n10674)
         );
  OAI22_X1 U2862 ( .A1(n8881), .A2(n259), .B1(n14815), .B2(n260), .ZN(n10675)
         );
  OAI22_X1 U2863 ( .A1(n8865), .A2(n259), .B1(n14775), .B2(n260), .ZN(n10676)
         );
  OAI22_X1 U2864 ( .A1(n8849), .A2(n259), .B1(n14735), .B2(n260), .ZN(n10677)
         );
  OAI22_X1 U2865 ( .A1(n8833), .A2(n259), .B1(n14695), .B2(n260), .ZN(n10678)
         );
  OAI22_X1 U2866 ( .A1(n8817), .A2(n259), .B1(n14655), .B2(n260), .ZN(n10679)
         );
  OAI22_X1 U2867 ( .A1(n8801), .A2(n261), .B1(n14953), .B2(n262), .ZN(n10680)
         );
  OAI22_X1 U2868 ( .A1(n8785), .A2(n261), .B1(n14895), .B2(n262), .ZN(n10681)
         );
  OAI22_X1 U2869 ( .A1(n8769), .A2(n261), .B1(n14855), .B2(n262), .ZN(n10682)
         );
  OAI22_X1 U2870 ( .A1(n8753), .A2(n261), .B1(n14815), .B2(n262), .ZN(n10683)
         );
  OAI22_X1 U2871 ( .A1(n8737), .A2(n261), .B1(n14775), .B2(n262), .ZN(n10684)
         );
  OAI22_X1 U2872 ( .A1(n8721), .A2(n261), .B1(n14735), .B2(n262), .ZN(n10685)
         );
  OAI22_X1 U2873 ( .A1(n8705), .A2(n261), .B1(n14695), .B2(n262), .ZN(n10686)
         );
  OAI22_X1 U2874 ( .A1(n8689), .A2(n261), .B1(n14655), .B2(n262), .ZN(n10687)
         );
  OAI22_X1 U2875 ( .A1(n8673), .A2(n263), .B1(n14953), .B2(n264), .ZN(n10688)
         );
  OAI22_X1 U2876 ( .A1(n8657), .A2(n263), .B1(n14895), .B2(n264), .ZN(n10689)
         );
  OAI22_X1 U2877 ( .A1(n8641), .A2(n263), .B1(n14855), .B2(n264), .ZN(n10690)
         );
  OAI22_X1 U2878 ( .A1(n8625), .A2(n263), .B1(n14815), .B2(n264), .ZN(n10691)
         );
  OAI22_X1 U2879 ( .A1(n8609), .A2(n263), .B1(n14775), .B2(n264), .ZN(n10692)
         );
  OAI22_X1 U2880 ( .A1(n8593), .A2(n263), .B1(n14735), .B2(n264), .ZN(n10693)
         );
  OAI22_X1 U2881 ( .A1(n8577), .A2(n263), .B1(n14695), .B2(n264), .ZN(n10694)
         );
  OAI22_X1 U2882 ( .A1(n8561), .A2(n263), .B1(n14655), .B2(n264), .ZN(n10695)
         );
  OAI22_X1 U2883 ( .A1(n8545), .A2(n265), .B1(n14953), .B2(n266), .ZN(n10696)
         );
  OAI22_X1 U2884 ( .A1(n8529), .A2(n265), .B1(n14895), .B2(n266), .ZN(n10697)
         );
  OAI22_X1 U2885 ( .A1(n8513), .A2(n265), .B1(n14855), .B2(n266), .ZN(n10698)
         );
  OAI22_X1 U2886 ( .A1(n8497), .A2(n265), .B1(n14815), .B2(n266), .ZN(n10699)
         );
  OAI22_X1 U2887 ( .A1(n8481), .A2(n265), .B1(n14775), .B2(n266), .ZN(n10700)
         );
  OAI22_X1 U2888 ( .A1(n8465), .A2(n265), .B1(n14735), .B2(n266), .ZN(n10701)
         );
  OAI22_X1 U2889 ( .A1(n8449), .A2(n265), .B1(n14695), .B2(n266), .ZN(n10702)
         );
  OAI22_X1 U2890 ( .A1(n8433), .A2(n265), .B1(n14655), .B2(n266), .ZN(n10703)
         );
  OAI22_X1 U2891 ( .A1(n8417), .A2(n267), .B1(n14953), .B2(n268), .ZN(n10704)
         );
  OAI22_X1 U2892 ( .A1(n8401), .A2(n267), .B1(n14895), .B2(n268), .ZN(n10705)
         );
  OAI22_X1 U2893 ( .A1(n8385), .A2(n267), .B1(n14855), .B2(n268), .ZN(n10706)
         );
  OAI22_X1 U2894 ( .A1(n8369), .A2(n267), .B1(n14815), .B2(n268), .ZN(n10707)
         );
  OAI22_X1 U2895 ( .A1(n8353), .A2(n267), .B1(n14775), .B2(n268), .ZN(n10708)
         );
  OAI22_X1 U2896 ( .A1(n8337), .A2(n267), .B1(n14735), .B2(n268), .ZN(n10709)
         );
  OAI22_X1 U2897 ( .A1(n8321), .A2(n267), .B1(n14695), .B2(n268), .ZN(n10710)
         );
  OAI22_X1 U2898 ( .A1(n8305), .A2(n267), .B1(n14655), .B2(n268), .ZN(n10711)
         );
  OAI22_X1 U2899 ( .A1(n8289), .A2(n269), .B1(n14953), .B2(n270), .ZN(n10712)
         );
  OAI22_X1 U2900 ( .A1(n8273), .A2(n269), .B1(n14896), .B2(n270), .ZN(n10713)
         );
  OAI22_X1 U2901 ( .A1(n8257), .A2(n269), .B1(n14856), .B2(n270), .ZN(n10714)
         );
  OAI22_X1 U2902 ( .A1(n8241), .A2(n269), .B1(n14816), .B2(n270), .ZN(n10715)
         );
  OAI22_X1 U2903 ( .A1(n8225), .A2(n269), .B1(n14776), .B2(n270), .ZN(n10716)
         );
  OAI22_X1 U2904 ( .A1(n8209), .A2(n269), .B1(n14736), .B2(n270), .ZN(n10717)
         );
  OAI22_X1 U2905 ( .A1(n8193), .A2(n269), .B1(n14696), .B2(n270), .ZN(n10718)
         );
  OAI22_X1 U2906 ( .A1(n8177), .A2(n269), .B1(n14656), .B2(n270), .ZN(n10719)
         );
  OAI22_X1 U2907 ( .A1(n8161), .A2(n271), .B1(n14953), .B2(n272), .ZN(n10720)
         );
  OAI22_X1 U2908 ( .A1(n8145), .A2(n271), .B1(n14896), .B2(n272), .ZN(n10721)
         );
  OAI22_X1 U2909 ( .A1(n8129), .A2(n271), .B1(n14856), .B2(n272), .ZN(n10722)
         );
  OAI22_X1 U2910 ( .A1(n8113), .A2(n271), .B1(n14816), .B2(n272), .ZN(n10723)
         );
  OAI22_X1 U2911 ( .A1(n8097), .A2(n271), .B1(n14776), .B2(n272), .ZN(n10724)
         );
  OAI22_X1 U2912 ( .A1(n8081), .A2(n271), .B1(n14736), .B2(n272), .ZN(n10725)
         );
  OAI22_X1 U2913 ( .A1(n8065), .A2(n271), .B1(n14696), .B2(n272), .ZN(n10726)
         );
  OAI22_X1 U2914 ( .A1(n8049), .A2(n271), .B1(n14656), .B2(n272), .ZN(n10727)
         );
  OAI22_X1 U2915 ( .A1(n8033), .A2(n273), .B1(n14953), .B2(n274), .ZN(n10728)
         );
  OAI22_X1 U2916 ( .A1(n8017), .A2(n273), .B1(n14896), .B2(n274), .ZN(n10729)
         );
  OAI22_X1 U2917 ( .A1(n8001), .A2(n273), .B1(n14856), .B2(n274), .ZN(n10730)
         );
  OAI22_X1 U2918 ( .A1(n7985), .A2(n273), .B1(n14816), .B2(n274), .ZN(n10731)
         );
  OAI22_X1 U2919 ( .A1(n7969), .A2(n273), .B1(n14776), .B2(n274), .ZN(n10732)
         );
  OAI22_X1 U2920 ( .A1(n7953), .A2(n273), .B1(n14736), .B2(n274), .ZN(n10733)
         );
  OAI22_X1 U2921 ( .A1(n7937), .A2(n273), .B1(n14696), .B2(n274), .ZN(n10734)
         );
  OAI22_X1 U2922 ( .A1(n7921), .A2(n273), .B1(n14656), .B2(n274), .ZN(n10735)
         );
  OAI22_X1 U2923 ( .A1(n7905), .A2(n275), .B1(n14953), .B2(n276), .ZN(n10736)
         );
  OAI22_X1 U2924 ( .A1(n7889), .A2(n275), .B1(n14896), .B2(n276), .ZN(n10737)
         );
  OAI22_X1 U2925 ( .A1(n7873), .A2(n275), .B1(n14856), .B2(n276), .ZN(n10738)
         );
  OAI22_X1 U2926 ( .A1(n7857), .A2(n275), .B1(n14816), .B2(n276), .ZN(n10739)
         );
  OAI22_X1 U2927 ( .A1(n7841), .A2(n275), .B1(n14776), .B2(n276), .ZN(n10740)
         );
  OAI22_X1 U2928 ( .A1(n7825), .A2(n275), .B1(n14736), .B2(n276), .ZN(n10741)
         );
  OAI22_X1 U2929 ( .A1(n7809), .A2(n275), .B1(n14696), .B2(n276), .ZN(n10742)
         );
  OAI22_X1 U2930 ( .A1(n7793), .A2(n275), .B1(n14656), .B2(n276), .ZN(n10743)
         );
  OAI22_X1 U2931 ( .A1(n7777), .A2(n277), .B1(n14953), .B2(n278), .ZN(n10744)
         );
  OAI22_X1 U2932 ( .A1(n7761), .A2(n277), .B1(n14896), .B2(n278), .ZN(n10745)
         );
  OAI22_X1 U2933 ( .A1(n7745), .A2(n277), .B1(n14856), .B2(n278), .ZN(n10746)
         );
  OAI22_X1 U2934 ( .A1(n7729), .A2(n277), .B1(n14816), .B2(n278), .ZN(n10747)
         );
  OAI22_X1 U2935 ( .A1(n7713), .A2(n277), .B1(n14776), .B2(n278), .ZN(n10748)
         );
  OAI22_X1 U2936 ( .A1(n7697), .A2(n277), .B1(n14736), .B2(n278), .ZN(n10749)
         );
  OAI22_X1 U2937 ( .A1(n7681), .A2(n277), .B1(n14696), .B2(n278), .ZN(n10750)
         );
  OAI22_X1 U2938 ( .A1(n7665), .A2(n277), .B1(n14656), .B2(n278), .ZN(n10751)
         );
  OAI22_X1 U2939 ( .A1(n7649), .A2(n279), .B1(n14953), .B2(n280), .ZN(n10752)
         );
  OAI22_X1 U2940 ( .A1(n7633), .A2(n279), .B1(n14896), .B2(n280), .ZN(n10753)
         );
  OAI22_X1 U2941 ( .A1(n7617), .A2(n279), .B1(n14856), .B2(n280), .ZN(n10754)
         );
  OAI22_X1 U2942 ( .A1(n7601), .A2(n279), .B1(n14816), .B2(n280), .ZN(n10755)
         );
  OAI22_X1 U2943 ( .A1(n7585), .A2(n279), .B1(n14776), .B2(n280), .ZN(n10756)
         );
  OAI22_X1 U2944 ( .A1(n7569), .A2(n279), .B1(n14736), .B2(n280), .ZN(n10757)
         );
  OAI22_X1 U2945 ( .A1(n7553), .A2(n279), .B1(n14696), .B2(n280), .ZN(n10758)
         );
  OAI22_X1 U2946 ( .A1(n7537), .A2(n279), .B1(n14656), .B2(n280), .ZN(n10759)
         );
  OAI22_X1 U2947 ( .A1(n7521), .A2(n281), .B1(n14953), .B2(n282), .ZN(n10760)
         );
  OAI22_X1 U2948 ( .A1(n7505), .A2(n281), .B1(n14896), .B2(n282), .ZN(n10761)
         );
  OAI22_X1 U2949 ( .A1(n7489), .A2(n281), .B1(n14856), .B2(n282), .ZN(n10762)
         );
  OAI22_X1 U2950 ( .A1(n7473), .A2(n281), .B1(n14816), .B2(n282), .ZN(n10763)
         );
  OAI22_X1 U2951 ( .A1(n7457), .A2(n281), .B1(n14776), .B2(n282), .ZN(n10764)
         );
  OAI22_X1 U2952 ( .A1(n7441), .A2(n281), .B1(n14736), .B2(n282), .ZN(n10765)
         );
  OAI22_X1 U2953 ( .A1(n7425), .A2(n281), .B1(n14696), .B2(n282), .ZN(n10766)
         );
  OAI22_X1 U2954 ( .A1(n7409), .A2(n281), .B1(n14656), .B2(n282), .ZN(n10767)
         );
  OAI22_X1 U2955 ( .A1(n7393), .A2(n283), .B1(n14952), .B2(n284), .ZN(n10768)
         );
  OAI22_X1 U2956 ( .A1(n7377), .A2(n283), .B1(n14896), .B2(n284), .ZN(n10769)
         );
  OAI22_X1 U2957 ( .A1(n7361), .A2(n283), .B1(n14856), .B2(n284), .ZN(n10770)
         );
  OAI22_X1 U2958 ( .A1(n7345), .A2(n283), .B1(n14816), .B2(n284), .ZN(n10771)
         );
  OAI22_X1 U2959 ( .A1(n7329), .A2(n283), .B1(n14776), .B2(n284), .ZN(n10772)
         );
  OAI22_X1 U2960 ( .A1(n7313), .A2(n283), .B1(n14736), .B2(n284), .ZN(n10773)
         );
  OAI22_X1 U2961 ( .A1(n7297), .A2(n283), .B1(n14696), .B2(n284), .ZN(n10774)
         );
  OAI22_X1 U2962 ( .A1(n7281), .A2(n283), .B1(n14656), .B2(n284), .ZN(n10775)
         );
  OAI22_X1 U2963 ( .A1(n7265), .A2(n285), .B1(n14952), .B2(n286), .ZN(n10776)
         );
  OAI22_X1 U2964 ( .A1(n7249), .A2(n285), .B1(n14896), .B2(n286), .ZN(n10777)
         );
  OAI22_X1 U2965 ( .A1(n7233), .A2(n285), .B1(n14856), .B2(n286), .ZN(n10778)
         );
  OAI22_X1 U2966 ( .A1(n7217), .A2(n285), .B1(n14816), .B2(n286), .ZN(n10779)
         );
  OAI22_X1 U2967 ( .A1(n7201), .A2(n285), .B1(n14776), .B2(n286), .ZN(n10780)
         );
  OAI22_X1 U2968 ( .A1(n7185), .A2(n285), .B1(n14736), .B2(n286), .ZN(n10781)
         );
  OAI22_X1 U2969 ( .A1(n7169), .A2(n285), .B1(n14696), .B2(n286), .ZN(n10782)
         );
  OAI22_X1 U2970 ( .A1(n7153), .A2(n285), .B1(n14656), .B2(n286), .ZN(n10783)
         );
  OAI22_X1 U2971 ( .A1(n7137), .A2(n287), .B1(n14952), .B2(n288), .ZN(n10784)
         );
  OAI22_X1 U2972 ( .A1(n7121), .A2(n287), .B1(n14896), .B2(n288), .ZN(n10785)
         );
  OAI22_X1 U2973 ( .A1(n7105), .A2(n287), .B1(n14856), .B2(n288), .ZN(n10786)
         );
  OAI22_X1 U2974 ( .A1(n7089), .A2(n287), .B1(n14816), .B2(n288), .ZN(n10787)
         );
  OAI22_X1 U2975 ( .A1(n7073), .A2(n287), .B1(n14776), .B2(n288), .ZN(n10788)
         );
  OAI22_X1 U2976 ( .A1(n7057), .A2(n287), .B1(n14736), .B2(n288), .ZN(n10789)
         );
  OAI22_X1 U2977 ( .A1(n7041), .A2(n287), .B1(n14696), .B2(n288), .ZN(n10790)
         );
  OAI22_X1 U2978 ( .A1(n7025), .A2(n287), .B1(n14656), .B2(n288), .ZN(n10791)
         );
  OAI22_X1 U2979 ( .A1(n7009), .A2(n289), .B1(n14952), .B2(n290), .ZN(n10792)
         );
  OAI22_X1 U2980 ( .A1(n6993), .A2(n289), .B1(n14896), .B2(n290), .ZN(n10793)
         );
  OAI22_X1 U2981 ( .A1(n6977), .A2(n289), .B1(n14856), .B2(n290), .ZN(n10794)
         );
  OAI22_X1 U2982 ( .A1(n6961), .A2(n289), .B1(n14816), .B2(n290), .ZN(n10795)
         );
  OAI22_X1 U2983 ( .A1(n6945), .A2(n289), .B1(n14776), .B2(n290), .ZN(n10796)
         );
  OAI22_X1 U2984 ( .A1(n6929), .A2(n289), .B1(n14736), .B2(n290), .ZN(n10797)
         );
  OAI22_X1 U2985 ( .A1(n6913), .A2(n289), .B1(n14696), .B2(n290), .ZN(n10798)
         );
  OAI22_X1 U2986 ( .A1(n6897), .A2(n289), .B1(n14656), .B2(n290), .ZN(n10799)
         );
  OAI22_X1 U2987 ( .A1(n6881), .A2(n291), .B1(n14952), .B2(n292), .ZN(n10800)
         );
  OAI22_X1 U2988 ( .A1(n6865), .A2(n291), .B1(n14896), .B2(n292), .ZN(n10801)
         );
  OAI22_X1 U2989 ( .A1(n6849), .A2(n291), .B1(n14856), .B2(n292), .ZN(n10802)
         );
  OAI22_X1 U2990 ( .A1(n6833), .A2(n291), .B1(n14816), .B2(n292), .ZN(n10803)
         );
  OAI22_X1 U2991 ( .A1(n6817), .A2(n291), .B1(n14776), .B2(n292), .ZN(n10804)
         );
  OAI22_X1 U2992 ( .A1(n6801), .A2(n291), .B1(n14736), .B2(n292), .ZN(n10805)
         );
  OAI22_X1 U2993 ( .A1(n6785), .A2(n291), .B1(n14696), .B2(n292), .ZN(n10806)
         );
  OAI22_X1 U2994 ( .A1(n6769), .A2(n291), .B1(n14656), .B2(n292), .ZN(n10807)
         );
  OAI22_X1 U2995 ( .A1(n6753), .A2(n293), .B1(n14952), .B2(n294), .ZN(n10808)
         );
  OAI22_X1 U2996 ( .A1(n6737), .A2(n293), .B1(n14896), .B2(n294), .ZN(n10809)
         );
  OAI22_X1 U2997 ( .A1(n6721), .A2(n293), .B1(n14856), .B2(n294), .ZN(n10810)
         );
  OAI22_X1 U2998 ( .A1(n6705), .A2(n293), .B1(n14816), .B2(n294), .ZN(n10811)
         );
  OAI22_X1 U2999 ( .A1(n6689), .A2(n293), .B1(n14776), .B2(n294), .ZN(n10812)
         );
  OAI22_X1 U3000 ( .A1(n6673), .A2(n293), .B1(n14736), .B2(n294), .ZN(n10813)
         );
  OAI22_X1 U3001 ( .A1(n6657), .A2(n293), .B1(n14696), .B2(n294), .ZN(n10814)
         );
  OAI22_X1 U3002 ( .A1(n6641), .A2(n293), .B1(n14656), .B2(n294), .ZN(n10815)
         );
  OAI22_X1 U3003 ( .A1(n6625), .A2(n295), .B1(n14952), .B2(n296), .ZN(n10816)
         );
  OAI22_X1 U3004 ( .A1(n6609), .A2(n295), .B1(n14897), .B2(n296), .ZN(n10817)
         );
  OAI22_X1 U3005 ( .A1(n6593), .A2(n295), .B1(n14857), .B2(n296), .ZN(n10818)
         );
  OAI22_X1 U3006 ( .A1(n6577), .A2(n295), .B1(n14817), .B2(n296), .ZN(n10819)
         );
  OAI22_X1 U3007 ( .A1(n6561), .A2(n295), .B1(n14777), .B2(n296), .ZN(n10820)
         );
  OAI22_X1 U3008 ( .A1(n6545), .A2(n295), .B1(n14737), .B2(n296), .ZN(n10821)
         );
  OAI22_X1 U3009 ( .A1(n6529), .A2(n295), .B1(n14697), .B2(n296), .ZN(n10822)
         );
  OAI22_X1 U3010 ( .A1(n6513), .A2(n295), .B1(n14657), .B2(n296), .ZN(n10823)
         );
  OAI22_X1 U3011 ( .A1(n6497), .A2(n297), .B1(n14952), .B2(n298), .ZN(n10824)
         );
  OAI22_X1 U3012 ( .A1(n6481), .A2(n297), .B1(n14897), .B2(n298), .ZN(n10825)
         );
  OAI22_X1 U3013 ( .A1(n6465), .A2(n297), .B1(n14857), .B2(n298), .ZN(n10826)
         );
  OAI22_X1 U3014 ( .A1(n6449), .A2(n297), .B1(n14817), .B2(n298), .ZN(n10827)
         );
  OAI22_X1 U3015 ( .A1(n6433), .A2(n297), .B1(n14777), .B2(n298), .ZN(n10828)
         );
  OAI22_X1 U3016 ( .A1(n6417), .A2(n297), .B1(n14737), .B2(n298), .ZN(n10829)
         );
  OAI22_X1 U3017 ( .A1(n6401), .A2(n297), .B1(n14697), .B2(n298), .ZN(n10830)
         );
  OAI22_X1 U3018 ( .A1(n6385), .A2(n297), .B1(n14657), .B2(n298), .ZN(n10831)
         );
  OAI22_X1 U3019 ( .A1(n6369), .A2(n299), .B1(n14952), .B2(n300), .ZN(n10832)
         );
  OAI22_X1 U3020 ( .A1(n6353), .A2(n299), .B1(n14897), .B2(n300), .ZN(n10833)
         );
  OAI22_X1 U3021 ( .A1(n6337), .A2(n299), .B1(n14857), .B2(n300), .ZN(n10834)
         );
  OAI22_X1 U3022 ( .A1(n6321), .A2(n299), .B1(n14817), .B2(n300), .ZN(n10835)
         );
  OAI22_X1 U3023 ( .A1(n6305), .A2(n299), .B1(n14777), .B2(n300), .ZN(n10836)
         );
  OAI22_X1 U3024 ( .A1(n6289), .A2(n299), .B1(n14737), .B2(n300), .ZN(n10837)
         );
  OAI22_X1 U3025 ( .A1(n6273), .A2(n299), .B1(n14697), .B2(n300), .ZN(n10838)
         );
  OAI22_X1 U3026 ( .A1(n6257), .A2(n299), .B1(n14657), .B2(n300), .ZN(n10839)
         );
  OAI22_X1 U3027 ( .A1(n6241), .A2(n301), .B1(n14952), .B2(n302), .ZN(n10840)
         );
  OAI22_X1 U3028 ( .A1(n6225), .A2(n301), .B1(n14897), .B2(n302), .ZN(n10841)
         );
  OAI22_X1 U3029 ( .A1(n6209), .A2(n301), .B1(n14857), .B2(n302), .ZN(n10842)
         );
  OAI22_X1 U3030 ( .A1(n6193), .A2(n301), .B1(n14817), .B2(n302), .ZN(n10843)
         );
  OAI22_X1 U3031 ( .A1(n6177), .A2(n301), .B1(n14777), .B2(n302), .ZN(n10844)
         );
  OAI22_X1 U3032 ( .A1(n6161), .A2(n301), .B1(n14737), .B2(n302), .ZN(n10845)
         );
  OAI22_X1 U3033 ( .A1(n6145), .A2(n301), .B1(n14697), .B2(n302), .ZN(n10846)
         );
  OAI22_X1 U3034 ( .A1(n6129), .A2(n301), .B1(n14657), .B2(n302), .ZN(n10847)
         );
  OAI22_X1 U3035 ( .A1(n6113), .A2(n303), .B1(n14952), .B2(n304), .ZN(n10848)
         );
  OAI22_X1 U3036 ( .A1(n6097), .A2(n303), .B1(n14897), .B2(n304), .ZN(n10849)
         );
  OAI22_X1 U3037 ( .A1(n6081), .A2(n303), .B1(n14857), .B2(n304), .ZN(n10850)
         );
  OAI22_X1 U3038 ( .A1(n6065), .A2(n303), .B1(n14817), .B2(n304), .ZN(n10851)
         );
  OAI22_X1 U3039 ( .A1(n6049), .A2(n303), .B1(n14777), .B2(n304), .ZN(n10852)
         );
  OAI22_X1 U3040 ( .A1(n6033), .A2(n303), .B1(n14737), .B2(n304), .ZN(n10853)
         );
  OAI22_X1 U3041 ( .A1(n6017), .A2(n303), .B1(n14697), .B2(n304), .ZN(n10854)
         );
  OAI22_X1 U3042 ( .A1(n6001), .A2(n303), .B1(n14657), .B2(n304), .ZN(n10855)
         );
  OAI22_X1 U3043 ( .A1(n9315), .A2(n515), .B1(n14963), .B2(n516), .ZN(n11672)
         );
  OAI22_X1 U3044 ( .A1(n9299), .A2(n515), .B1(n14905), .B2(n516), .ZN(n11673)
         );
  OAI22_X1 U3045 ( .A1(n9283), .A2(n515), .B1(n14865), .B2(n516), .ZN(n11674)
         );
  OAI22_X1 U3046 ( .A1(n9267), .A2(n515), .B1(n14825), .B2(n516), .ZN(n11675)
         );
  OAI22_X1 U3047 ( .A1(n9251), .A2(n515), .B1(n14785), .B2(n516), .ZN(n11676)
         );
  OAI22_X1 U3048 ( .A1(n9235), .A2(n515), .B1(n14745), .B2(n516), .ZN(n11677)
         );
  OAI22_X1 U3049 ( .A1(n9219), .A2(n515), .B1(n14705), .B2(n516), .ZN(n11678)
         );
  OAI22_X1 U3050 ( .A1(n9203), .A2(n515), .B1(n14665), .B2(n516), .ZN(n11679)
         );
  OAI22_X1 U3051 ( .A1(n9187), .A2(n517), .B1(n14963), .B2(n518), .ZN(n11680)
         );
  OAI22_X1 U3052 ( .A1(n9171), .A2(n517), .B1(n14905), .B2(n518), .ZN(n11681)
         );
  OAI22_X1 U3053 ( .A1(n9155), .A2(n517), .B1(n14865), .B2(n518), .ZN(n11682)
         );
  OAI22_X1 U3054 ( .A1(n9139), .A2(n517), .B1(n14825), .B2(n518), .ZN(n11683)
         );
  OAI22_X1 U3055 ( .A1(n9123), .A2(n517), .B1(n14785), .B2(n518), .ZN(n11684)
         );
  OAI22_X1 U3056 ( .A1(n9107), .A2(n517), .B1(n14745), .B2(n518), .ZN(n11685)
         );
  OAI22_X1 U3057 ( .A1(n9091), .A2(n517), .B1(n14705), .B2(n518), .ZN(n11686)
         );
  OAI22_X1 U3058 ( .A1(n9075), .A2(n517), .B1(n14665), .B2(n518), .ZN(n11687)
         );
  OAI22_X1 U3059 ( .A1(n9059), .A2(n519), .B1(n14963), .B2(n520), .ZN(n11688)
         );
  OAI22_X1 U3060 ( .A1(n9043), .A2(n519), .B1(n14905), .B2(n520), .ZN(n11689)
         );
  OAI22_X1 U3061 ( .A1(n9027), .A2(n519), .B1(n14865), .B2(n520), .ZN(n11690)
         );
  OAI22_X1 U3062 ( .A1(n9011), .A2(n519), .B1(n14825), .B2(n520), .ZN(n11691)
         );
  OAI22_X1 U3063 ( .A1(n8995), .A2(n519), .B1(n14785), .B2(n520), .ZN(n11692)
         );
  OAI22_X1 U3064 ( .A1(n8979), .A2(n519), .B1(n14745), .B2(n520), .ZN(n11693)
         );
  OAI22_X1 U3065 ( .A1(n8963), .A2(n519), .B1(n14705), .B2(n520), .ZN(n11694)
         );
  OAI22_X1 U3066 ( .A1(n8947), .A2(n519), .B1(n14665), .B2(n520), .ZN(n11695)
         );
  OAI22_X1 U3067 ( .A1(n8931), .A2(n521), .B1(n14963), .B2(n522), .ZN(n11696)
         );
  OAI22_X1 U3068 ( .A1(n8915), .A2(n521), .B1(n14905), .B2(n522), .ZN(n11697)
         );
  OAI22_X1 U3069 ( .A1(n8899), .A2(n521), .B1(n14865), .B2(n522), .ZN(n11698)
         );
  OAI22_X1 U3070 ( .A1(n8883), .A2(n521), .B1(n14825), .B2(n522), .ZN(n11699)
         );
  OAI22_X1 U3071 ( .A1(n8867), .A2(n521), .B1(n14785), .B2(n522), .ZN(n11700)
         );
  OAI22_X1 U3072 ( .A1(n8851), .A2(n521), .B1(n14745), .B2(n522), .ZN(n11701)
         );
  OAI22_X1 U3073 ( .A1(n8835), .A2(n521), .B1(n14705), .B2(n522), .ZN(n11702)
         );
  OAI22_X1 U3074 ( .A1(n8819), .A2(n521), .B1(n14665), .B2(n522), .ZN(n11703)
         );
  OAI22_X1 U3075 ( .A1(n8803), .A2(n523), .B1(n14963), .B2(n524), .ZN(n11704)
         );
  OAI22_X1 U3076 ( .A1(n8787), .A2(n523), .B1(n14905), .B2(n524), .ZN(n11705)
         );
  OAI22_X1 U3077 ( .A1(n8771), .A2(n523), .B1(n14865), .B2(n524), .ZN(n11706)
         );
  OAI22_X1 U3078 ( .A1(n8755), .A2(n523), .B1(n14825), .B2(n524), .ZN(n11707)
         );
  OAI22_X1 U3079 ( .A1(n8739), .A2(n523), .B1(n14785), .B2(n524), .ZN(n11708)
         );
  OAI22_X1 U3080 ( .A1(n8723), .A2(n523), .B1(n14745), .B2(n524), .ZN(n11709)
         );
  OAI22_X1 U3081 ( .A1(n8707), .A2(n523), .B1(n14705), .B2(n524), .ZN(n11710)
         );
  OAI22_X1 U3082 ( .A1(n8691), .A2(n523), .B1(n14665), .B2(n524), .ZN(n11711)
         );
  OAI22_X1 U3083 ( .A1(n8675), .A2(n525), .B1(n14963), .B2(n526), .ZN(n11712)
         );
  OAI22_X1 U3084 ( .A1(n8659), .A2(n525), .B1(n14905), .B2(n526), .ZN(n11713)
         );
  OAI22_X1 U3085 ( .A1(n8643), .A2(n525), .B1(n14865), .B2(n526), .ZN(n11714)
         );
  OAI22_X1 U3086 ( .A1(n8627), .A2(n525), .B1(n14825), .B2(n526), .ZN(n11715)
         );
  OAI22_X1 U3087 ( .A1(n8611), .A2(n525), .B1(n14785), .B2(n526), .ZN(n11716)
         );
  OAI22_X1 U3088 ( .A1(n8595), .A2(n525), .B1(n14745), .B2(n526), .ZN(n11717)
         );
  OAI22_X1 U3089 ( .A1(n8579), .A2(n525), .B1(n14705), .B2(n526), .ZN(n11718)
         );
  OAI22_X1 U3090 ( .A1(n8563), .A2(n525), .B1(n14665), .B2(n526), .ZN(n11719)
         );
  OAI22_X1 U3091 ( .A1(n8547), .A2(n527), .B1(n14963), .B2(n528), .ZN(n11720)
         );
  OAI22_X1 U3092 ( .A1(n8531), .A2(n527), .B1(n14905), .B2(n528), .ZN(n11721)
         );
  OAI22_X1 U3093 ( .A1(n8515), .A2(n527), .B1(n14865), .B2(n528), .ZN(n11722)
         );
  OAI22_X1 U3094 ( .A1(n8499), .A2(n527), .B1(n14825), .B2(n528), .ZN(n11723)
         );
  OAI22_X1 U3095 ( .A1(n8483), .A2(n527), .B1(n14785), .B2(n528), .ZN(n11724)
         );
  OAI22_X1 U3096 ( .A1(n8467), .A2(n527), .B1(n14745), .B2(n528), .ZN(n11725)
         );
  OAI22_X1 U3097 ( .A1(n8451), .A2(n527), .B1(n14705), .B2(n528), .ZN(n11726)
         );
  OAI22_X1 U3098 ( .A1(n8435), .A2(n527), .B1(n14665), .B2(n528), .ZN(n11727)
         );
  OAI22_X1 U3099 ( .A1(n8419), .A2(n529), .B1(n14963), .B2(n530), .ZN(n11728)
         );
  OAI22_X1 U3100 ( .A1(n8403), .A2(n529), .B1(n14905), .B2(n530), .ZN(n11729)
         );
  OAI22_X1 U3101 ( .A1(n8387), .A2(n529), .B1(n14865), .B2(n530), .ZN(n11730)
         );
  OAI22_X1 U3102 ( .A1(n8371), .A2(n529), .B1(n14825), .B2(n530), .ZN(n11731)
         );
  OAI22_X1 U3103 ( .A1(n8355), .A2(n529), .B1(n14785), .B2(n530), .ZN(n11732)
         );
  OAI22_X1 U3104 ( .A1(n8339), .A2(n529), .B1(n14745), .B2(n530), .ZN(n11733)
         );
  OAI22_X1 U3105 ( .A1(n8323), .A2(n529), .B1(n14705), .B2(n530), .ZN(n11734)
         );
  OAI22_X1 U3106 ( .A1(n8307), .A2(n529), .B1(n14665), .B2(n530), .ZN(n11735)
         );
  OAI22_X1 U3107 ( .A1(n8291), .A2(n531), .B1(n14963), .B2(n532), .ZN(n11736)
         );
  OAI22_X1 U3108 ( .A1(n8275), .A2(n531), .B1(n14905), .B2(n532), .ZN(n11737)
         );
  OAI22_X1 U3109 ( .A1(n8259), .A2(n531), .B1(n14865), .B2(n532), .ZN(n11738)
         );
  OAI22_X1 U3110 ( .A1(n8243), .A2(n531), .B1(n14825), .B2(n532), .ZN(n11739)
         );
  OAI22_X1 U3111 ( .A1(n8227), .A2(n531), .B1(n14785), .B2(n532), .ZN(n11740)
         );
  OAI22_X1 U3112 ( .A1(n8211), .A2(n531), .B1(n14745), .B2(n532), .ZN(n11741)
         );
  OAI22_X1 U3113 ( .A1(n8195), .A2(n531), .B1(n14705), .B2(n532), .ZN(n11742)
         );
  OAI22_X1 U3114 ( .A1(n8179), .A2(n531), .B1(n14665), .B2(n532), .ZN(n11743)
         );
  OAI22_X1 U3115 ( .A1(n8163), .A2(n533), .B1(n14963), .B2(n534), .ZN(n11744)
         );
  OAI22_X1 U3116 ( .A1(n8147), .A2(n533), .B1(n14905), .B2(n534), .ZN(n11745)
         );
  OAI22_X1 U3117 ( .A1(n8131), .A2(n533), .B1(n14865), .B2(n534), .ZN(n11746)
         );
  OAI22_X1 U3118 ( .A1(n8115), .A2(n533), .B1(n14825), .B2(n534), .ZN(n11747)
         );
  OAI22_X1 U3119 ( .A1(n8099), .A2(n533), .B1(n14785), .B2(n534), .ZN(n11748)
         );
  OAI22_X1 U3120 ( .A1(n8083), .A2(n533), .B1(n14745), .B2(n534), .ZN(n11749)
         );
  OAI22_X1 U3121 ( .A1(n8067), .A2(n533), .B1(n14705), .B2(n534), .ZN(n11750)
         );
  OAI22_X1 U3122 ( .A1(n8051), .A2(n533), .B1(n14665), .B2(n534), .ZN(n11751)
         );
  OAI22_X1 U3123 ( .A1(n8035), .A2(n535), .B1(n14963), .B2(n536), .ZN(n11752)
         );
  OAI22_X1 U3124 ( .A1(n8019), .A2(n535), .B1(n14906), .B2(n536), .ZN(n11753)
         );
  OAI22_X1 U3125 ( .A1(n8003), .A2(n535), .B1(n14866), .B2(n536), .ZN(n11754)
         );
  OAI22_X1 U3126 ( .A1(n7987), .A2(n535), .B1(n14826), .B2(n536), .ZN(n11755)
         );
  OAI22_X1 U3127 ( .A1(n7971), .A2(n535), .B1(n14786), .B2(n536), .ZN(n11756)
         );
  OAI22_X1 U3128 ( .A1(n7955), .A2(n535), .B1(n14746), .B2(n536), .ZN(n11757)
         );
  OAI22_X1 U3129 ( .A1(n7939), .A2(n535), .B1(n14706), .B2(n536), .ZN(n11758)
         );
  OAI22_X1 U3130 ( .A1(n7923), .A2(n535), .B1(n14666), .B2(n536), .ZN(n11759)
         );
  OAI22_X1 U3131 ( .A1(n7907), .A2(n537), .B1(n14963), .B2(n538), .ZN(n11760)
         );
  OAI22_X1 U3132 ( .A1(n7891), .A2(n537), .B1(n14906), .B2(n538), .ZN(n11761)
         );
  OAI22_X1 U3133 ( .A1(n7875), .A2(n537), .B1(n14866), .B2(n538), .ZN(n11762)
         );
  OAI22_X1 U3134 ( .A1(n7859), .A2(n537), .B1(n14826), .B2(n538), .ZN(n11763)
         );
  OAI22_X1 U3135 ( .A1(n7843), .A2(n537), .B1(n14786), .B2(n538), .ZN(n11764)
         );
  OAI22_X1 U3136 ( .A1(n7827), .A2(n537), .B1(n14746), .B2(n538), .ZN(n11765)
         );
  OAI22_X1 U3137 ( .A1(n7811), .A2(n537), .B1(n14706), .B2(n538), .ZN(n11766)
         );
  OAI22_X1 U3138 ( .A1(n7795), .A2(n537), .B1(n14666), .B2(n538), .ZN(n11767)
         );
  OAI22_X1 U3139 ( .A1(n7779), .A2(n539), .B1(n14962), .B2(n540), .ZN(n11768)
         );
  OAI22_X1 U3140 ( .A1(n7763), .A2(n539), .B1(n14906), .B2(n540), .ZN(n11769)
         );
  OAI22_X1 U3141 ( .A1(n7747), .A2(n539), .B1(n14866), .B2(n540), .ZN(n11770)
         );
  OAI22_X1 U3142 ( .A1(n7731), .A2(n539), .B1(n14826), .B2(n540), .ZN(n11771)
         );
  OAI22_X1 U3143 ( .A1(n7715), .A2(n539), .B1(n14786), .B2(n540), .ZN(n11772)
         );
  OAI22_X1 U3144 ( .A1(n7699), .A2(n539), .B1(n14746), .B2(n540), .ZN(n11773)
         );
  OAI22_X1 U3145 ( .A1(n7683), .A2(n539), .B1(n14706), .B2(n540), .ZN(n11774)
         );
  OAI22_X1 U3146 ( .A1(n7667), .A2(n539), .B1(n14666), .B2(n540), .ZN(n11775)
         );
  OAI22_X1 U3147 ( .A1(n7651), .A2(n541), .B1(n14962), .B2(n542), .ZN(n11776)
         );
  OAI22_X1 U3148 ( .A1(n7635), .A2(n541), .B1(n14906), .B2(n542), .ZN(n11777)
         );
  OAI22_X1 U3149 ( .A1(n7619), .A2(n541), .B1(n14866), .B2(n542), .ZN(n11778)
         );
  OAI22_X1 U3150 ( .A1(n7603), .A2(n541), .B1(n14826), .B2(n542), .ZN(n11779)
         );
  OAI22_X1 U3151 ( .A1(n7587), .A2(n541), .B1(n14786), .B2(n542), .ZN(n11780)
         );
  OAI22_X1 U3152 ( .A1(n7571), .A2(n541), .B1(n14746), .B2(n542), .ZN(n11781)
         );
  OAI22_X1 U3153 ( .A1(n7555), .A2(n541), .B1(n14706), .B2(n542), .ZN(n11782)
         );
  OAI22_X1 U3154 ( .A1(n7539), .A2(n541), .B1(n14666), .B2(n542), .ZN(n11783)
         );
  OAI22_X1 U3155 ( .A1(n7523), .A2(n543), .B1(n14962), .B2(n544), .ZN(n11784)
         );
  OAI22_X1 U3156 ( .A1(n7507), .A2(n543), .B1(n14906), .B2(n544), .ZN(n11785)
         );
  OAI22_X1 U3157 ( .A1(n7491), .A2(n543), .B1(n14866), .B2(n544), .ZN(n11786)
         );
  OAI22_X1 U3158 ( .A1(n7475), .A2(n543), .B1(n14826), .B2(n544), .ZN(n11787)
         );
  OAI22_X1 U3159 ( .A1(n7459), .A2(n543), .B1(n14786), .B2(n544), .ZN(n11788)
         );
  OAI22_X1 U3160 ( .A1(n7443), .A2(n543), .B1(n14746), .B2(n544), .ZN(n11789)
         );
  OAI22_X1 U3161 ( .A1(n7427), .A2(n543), .B1(n14706), .B2(n544), .ZN(n11790)
         );
  OAI22_X1 U3162 ( .A1(n7411), .A2(n543), .B1(n14666), .B2(n544), .ZN(n11791)
         );
  OAI22_X1 U3163 ( .A1(n7395), .A2(n545), .B1(n14962), .B2(n546), .ZN(n11792)
         );
  OAI22_X1 U3164 ( .A1(n7379), .A2(n545), .B1(n14906), .B2(n546), .ZN(n11793)
         );
  OAI22_X1 U3165 ( .A1(n7363), .A2(n545), .B1(n14866), .B2(n546), .ZN(n11794)
         );
  OAI22_X1 U3166 ( .A1(n7347), .A2(n545), .B1(n14826), .B2(n546), .ZN(n11795)
         );
  OAI22_X1 U3167 ( .A1(n7331), .A2(n545), .B1(n14786), .B2(n546), .ZN(n11796)
         );
  OAI22_X1 U3168 ( .A1(n7315), .A2(n545), .B1(n14746), .B2(n546), .ZN(n11797)
         );
  OAI22_X1 U3169 ( .A1(n7299), .A2(n545), .B1(n14706), .B2(n546), .ZN(n11798)
         );
  OAI22_X1 U3170 ( .A1(n7283), .A2(n545), .B1(n14666), .B2(n546), .ZN(n11799)
         );
  OAI22_X1 U3171 ( .A1(n7267), .A2(n547), .B1(n14962), .B2(n548), .ZN(n11800)
         );
  OAI22_X1 U3172 ( .A1(n7251), .A2(n547), .B1(n14906), .B2(n548), .ZN(n11801)
         );
  OAI22_X1 U3173 ( .A1(n7235), .A2(n547), .B1(n14866), .B2(n548), .ZN(n11802)
         );
  OAI22_X1 U3174 ( .A1(n7219), .A2(n547), .B1(n14826), .B2(n548), .ZN(n11803)
         );
  OAI22_X1 U3175 ( .A1(n7203), .A2(n547), .B1(n14786), .B2(n548), .ZN(n11804)
         );
  OAI22_X1 U3176 ( .A1(n7187), .A2(n547), .B1(n14746), .B2(n548), .ZN(n11805)
         );
  OAI22_X1 U3177 ( .A1(n7171), .A2(n547), .B1(n14706), .B2(n548), .ZN(n11806)
         );
  OAI22_X1 U3178 ( .A1(n7155), .A2(n547), .B1(n14666), .B2(n548), .ZN(n11807)
         );
  OAI22_X1 U3179 ( .A1(n7139), .A2(n549), .B1(n14962), .B2(n550), .ZN(n11808)
         );
  OAI22_X1 U3180 ( .A1(n7123), .A2(n549), .B1(n14906), .B2(n550), .ZN(n11809)
         );
  OAI22_X1 U3181 ( .A1(n7107), .A2(n549), .B1(n14866), .B2(n550), .ZN(n11810)
         );
  OAI22_X1 U3182 ( .A1(n7091), .A2(n549), .B1(n14826), .B2(n550), .ZN(n11811)
         );
  OAI22_X1 U3183 ( .A1(n7075), .A2(n549), .B1(n14786), .B2(n550), .ZN(n11812)
         );
  OAI22_X1 U3184 ( .A1(n7059), .A2(n549), .B1(n14746), .B2(n550), .ZN(n11813)
         );
  OAI22_X1 U3185 ( .A1(n7043), .A2(n549), .B1(n14706), .B2(n550), .ZN(n11814)
         );
  OAI22_X1 U3186 ( .A1(n7027), .A2(n549), .B1(n14666), .B2(n550), .ZN(n11815)
         );
  OAI22_X1 U3187 ( .A1(n7011), .A2(n551), .B1(n14962), .B2(n552), .ZN(n11816)
         );
  OAI22_X1 U3188 ( .A1(n6995), .A2(n551), .B1(n14906), .B2(n552), .ZN(n11817)
         );
  OAI22_X1 U3189 ( .A1(n6979), .A2(n551), .B1(n14866), .B2(n552), .ZN(n11818)
         );
  OAI22_X1 U3190 ( .A1(n6963), .A2(n551), .B1(n14826), .B2(n552), .ZN(n11819)
         );
  OAI22_X1 U3191 ( .A1(n6947), .A2(n551), .B1(n14786), .B2(n552), .ZN(n11820)
         );
  OAI22_X1 U3192 ( .A1(n6931), .A2(n551), .B1(n14746), .B2(n552), .ZN(n11821)
         );
  OAI22_X1 U3193 ( .A1(n6915), .A2(n551), .B1(n14706), .B2(n552), .ZN(n11822)
         );
  OAI22_X1 U3194 ( .A1(n6899), .A2(n551), .B1(n14666), .B2(n552), .ZN(n11823)
         );
  OAI22_X1 U3195 ( .A1(n6883), .A2(n553), .B1(n14962), .B2(n554), .ZN(n11824)
         );
  OAI22_X1 U3196 ( .A1(n6867), .A2(n553), .B1(n14906), .B2(n554), .ZN(n11825)
         );
  OAI22_X1 U3197 ( .A1(n6851), .A2(n553), .B1(n14866), .B2(n554), .ZN(n11826)
         );
  OAI22_X1 U3198 ( .A1(n6835), .A2(n553), .B1(n14826), .B2(n554), .ZN(n11827)
         );
  OAI22_X1 U3199 ( .A1(n6819), .A2(n553), .B1(n14786), .B2(n554), .ZN(n11828)
         );
  OAI22_X1 U3200 ( .A1(n6803), .A2(n553), .B1(n14746), .B2(n554), .ZN(n11829)
         );
  OAI22_X1 U3201 ( .A1(n6787), .A2(n553), .B1(n14706), .B2(n554), .ZN(n11830)
         );
  OAI22_X1 U3202 ( .A1(n6771), .A2(n553), .B1(n14666), .B2(n554), .ZN(n11831)
         );
  OAI22_X1 U3203 ( .A1(n6755), .A2(n555), .B1(n14962), .B2(n556), .ZN(n11832)
         );
  OAI22_X1 U3204 ( .A1(n6739), .A2(n555), .B1(n14906), .B2(n556), .ZN(n11833)
         );
  OAI22_X1 U3205 ( .A1(n6723), .A2(n555), .B1(n14866), .B2(n556), .ZN(n11834)
         );
  OAI22_X1 U3206 ( .A1(n6707), .A2(n555), .B1(n14826), .B2(n556), .ZN(n11835)
         );
  OAI22_X1 U3207 ( .A1(n6691), .A2(n555), .B1(n14786), .B2(n556), .ZN(n11836)
         );
  OAI22_X1 U3208 ( .A1(n6675), .A2(n555), .B1(n14746), .B2(n556), .ZN(n11837)
         );
  OAI22_X1 U3209 ( .A1(n6659), .A2(n555), .B1(n14706), .B2(n556), .ZN(n11838)
         );
  OAI22_X1 U3210 ( .A1(n6643), .A2(n555), .B1(n14666), .B2(n556), .ZN(n11839)
         );
  OAI22_X1 U3211 ( .A1(n6627), .A2(n557), .B1(n14962), .B2(n558), .ZN(n11840)
         );
  OAI22_X1 U3212 ( .A1(n6611), .A2(n557), .B1(n14906), .B2(n558), .ZN(n11841)
         );
  OAI22_X1 U3213 ( .A1(n6595), .A2(n557), .B1(n14866), .B2(n558), .ZN(n11842)
         );
  OAI22_X1 U3214 ( .A1(n6579), .A2(n557), .B1(n14826), .B2(n558), .ZN(n11843)
         );
  OAI22_X1 U3215 ( .A1(n6563), .A2(n557), .B1(n14786), .B2(n558), .ZN(n11844)
         );
  OAI22_X1 U3216 ( .A1(n6547), .A2(n557), .B1(n14746), .B2(n558), .ZN(n11845)
         );
  OAI22_X1 U3217 ( .A1(n6531), .A2(n557), .B1(n14706), .B2(n558), .ZN(n11846)
         );
  OAI22_X1 U3218 ( .A1(n6515), .A2(n557), .B1(n14666), .B2(n558), .ZN(n11847)
         );
  OAI22_X1 U3219 ( .A1(n6499), .A2(n559), .B1(n14962), .B2(n560), .ZN(n11848)
         );
  OAI22_X1 U3220 ( .A1(n6483), .A2(n559), .B1(n14906), .B2(n560), .ZN(n11849)
         );
  OAI22_X1 U3221 ( .A1(n6467), .A2(n559), .B1(n14866), .B2(n560), .ZN(n11850)
         );
  OAI22_X1 U3222 ( .A1(n6451), .A2(n559), .B1(n14826), .B2(n560), .ZN(n11851)
         );
  OAI22_X1 U3223 ( .A1(n6435), .A2(n559), .B1(n14786), .B2(n560), .ZN(n11852)
         );
  OAI22_X1 U3224 ( .A1(n6419), .A2(n559), .B1(n14746), .B2(n560), .ZN(n11853)
         );
  OAI22_X1 U3225 ( .A1(n6403), .A2(n559), .B1(n14706), .B2(n560), .ZN(n11854)
         );
  OAI22_X1 U3226 ( .A1(n6387), .A2(n559), .B1(n14666), .B2(n560), .ZN(n11855)
         );
  OAI22_X1 U3227 ( .A1(n6371), .A2(n561), .B1(n14962), .B2(n562), .ZN(n11856)
         );
  OAI22_X1 U3228 ( .A1(n6355), .A2(n561), .B1(n14907), .B2(n562), .ZN(n11857)
         );
  OAI22_X1 U3229 ( .A1(n6339), .A2(n561), .B1(n14867), .B2(n562), .ZN(n11858)
         );
  OAI22_X1 U3230 ( .A1(n6323), .A2(n561), .B1(n14827), .B2(n562), .ZN(n11859)
         );
  OAI22_X1 U3231 ( .A1(n6307), .A2(n561), .B1(n14787), .B2(n562), .ZN(n11860)
         );
  OAI22_X1 U3232 ( .A1(n6291), .A2(n561), .B1(n14747), .B2(n562), .ZN(n11861)
         );
  OAI22_X1 U3233 ( .A1(n6275), .A2(n561), .B1(n14707), .B2(n562), .ZN(n11862)
         );
  OAI22_X1 U3234 ( .A1(n6259), .A2(n561), .B1(n14667), .B2(n562), .ZN(n11863)
         );
  OAI22_X1 U3235 ( .A1(n6243), .A2(n563), .B1(n14962), .B2(n564), .ZN(n11864)
         );
  OAI22_X1 U3236 ( .A1(n6227), .A2(n563), .B1(n14907), .B2(n564), .ZN(n11865)
         );
  OAI22_X1 U3237 ( .A1(n6211), .A2(n563), .B1(n14867), .B2(n564), .ZN(n11866)
         );
  OAI22_X1 U3238 ( .A1(n6195), .A2(n563), .B1(n14827), .B2(n564), .ZN(n11867)
         );
  OAI22_X1 U3239 ( .A1(n6179), .A2(n563), .B1(n14787), .B2(n564), .ZN(n11868)
         );
  OAI22_X1 U3240 ( .A1(n6163), .A2(n563), .B1(n14747), .B2(n564), .ZN(n11869)
         );
  OAI22_X1 U3241 ( .A1(n6147), .A2(n563), .B1(n14707), .B2(n564), .ZN(n11870)
         );
  OAI22_X1 U3242 ( .A1(n6131), .A2(n563), .B1(n14667), .B2(n564), .ZN(n11871)
         );
  OAI22_X1 U3243 ( .A1(n6115), .A2(n565), .B1(n14961), .B2(n566), .ZN(n11872)
         );
  OAI22_X1 U3244 ( .A1(n6099), .A2(n565), .B1(n14907), .B2(n566), .ZN(n11873)
         );
  OAI22_X1 U3245 ( .A1(n6083), .A2(n565), .B1(n14867), .B2(n566), .ZN(n11874)
         );
  OAI22_X1 U3246 ( .A1(n6067), .A2(n565), .B1(n14827), .B2(n566), .ZN(n11875)
         );
  OAI22_X1 U3247 ( .A1(n6051), .A2(n565), .B1(n14787), .B2(n566), .ZN(n11876)
         );
  OAI22_X1 U3248 ( .A1(n6035), .A2(n565), .B1(n14747), .B2(n566), .ZN(n11877)
         );
  OAI22_X1 U3249 ( .A1(n6019), .A2(n565), .B1(n14707), .B2(n566), .ZN(n11878)
         );
  OAI22_X1 U3250 ( .A1(n6003), .A2(n565), .B1(n14667), .B2(n566), .ZN(n11879)
         );
  OAI22_X1 U3251 ( .A1(n9319), .A2(n580), .B1(n14961), .B2(n581), .ZN(n11928)
         );
  OAI22_X1 U3252 ( .A1(n9303), .A2(n580), .B1(n14907), .B2(n581), .ZN(n11929)
         );
  OAI22_X1 U3253 ( .A1(n9287), .A2(n580), .B1(n14867), .B2(n581), .ZN(n11930)
         );
  OAI22_X1 U3254 ( .A1(n9271), .A2(n580), .B1(n14827), .B2(n581), .ZN(n11931)
         );
  OAI22_X1 U3255 ( .A1(n9255), .A2(n580), .B1(n14787), .B2(n581), .ZN(n11932)
         );
  OAI22_X1 U3256 ( .A1(n9239), .A2(n580), .B1(n14747), .B2(n581), .ZN(n11933)
         );
  OAI22_X1 U3257 ( .A1(n9223), .A2(n580), .B1(n14707), .B2(n581), .ZN(n11934)
         );
  OAI22_X1 U3258 ( .A1(n9207), .A2(n580), .B1(n14667), .B2(n581), .ZN(n11935)
         );
  OAI22_X1 U3259 ( .A1(n9191), .A2(n582), .B1(n14961), .B2(n583), .ZN(n11936)
         );
  OAI22_X1 U3260 ( .A1(n9175), .A2(n582), .B1(n14907), .B2(n583), .ZN(n11937)
         );
  OAI22_X1 U3261 ( .A1(n9159), .A2(n582), .B1(n14867), .B2(n583), .ZN(n11938)
         );
  OAI22_X1 U3262 ( .A1(n9143), .A2(n582), .B1(n14827), .B2(n583), .ZN(n11939)
         );
  OAI22_X1 U3263 ( .A1(n9127), .A2(n582), .B1(n14787), .B2(n583), .ZN(n11940)
         );
  OAI22_X1 U3264 ( .A1(n9111), .A2(n582), .B1(n14747), .B2(n583), .ZN(n11941)
         );
  OAI22_X1 U3265 ( .A1(n9095), .A2(n582), .B1(n14707), .B2(n583), .ZN(n11942)
         );
  OAI22_X1 U3266 ( .A1(n9079), .A2(n582), .B1(n14667), .B2(n583), .ZN(n11943)
         );
  OAI22_X1 U3267 ( .A1(n9063), .A2(n584), .B1(n14961), .B2(n585), .ZN(n11944)
         );
  OAI22_X1 U3268 ( .A1(n9047), .A2(n584), .B1(n14907), .B2(n585), .ZN(n11945)
         );
  OAI22_X1 U3269 ( .A1(n9031), .A2(n584), .B1(n14867), .B2(n585), .ZN(n11946)
         );
  OAI22_X1 U3270 ( .A1(n9015), .A2(n584), .B1(n14827), .B2(n585), .ZN(n11947)
         );
  OAI22_X1 U3271 ( .A1(n8999), .A2(n584), .B1(n14787), .B2(n585), .ZN(n11948)
         );
  OAI22_X1 U3272 ( .A1(n8983), .A2(n584), .B1(n14747), .B2(n585), .ZN(n11949)
         );
  OAI22_X1 U3273 ( .A1(n8967), .A2(n584), .B1(n14707), .B2(n585), .ZN(n11950)
         );
  OAI22_X1 U3274 ( .A1(n8951), .A2(n584), .B1(n14667), .B2(n585), .ZN(n11951)
         );
  OAI22_X1 U3275 ( .A1(n8935), .A2(n586), .B1(n14961), .B2(n587), .ZN(n11952)
         );
  OAI22_X1 U3276 ( .A1(n8919), .A2(n586), .B1(n14907), .B2(n587), .ZN(n11953)
         );
  OAI22_X1 U3277 ( .A1(n8903), .A2(n586), .B1(n14867), .B2(n587), .ZN(n11954)
         );
  OAI22_X1 U3278 ( .A1(n8887), .A2(n586), .B1(n14827), .B2(n587), .ZN(n11955)
         );
  OAI22_X1 U3279 ( .A1(n8871), .A2(n586), .B1(n14787), .B2(n587), .ZN(n11956)
         );
  OAI22_X1 U3280 ( .A1(n8855), .A2(n586), .B1(n14747), .B2(n587), .ZN(n11957)
         );
  OAI22_X1 U3281 ( .A1(n8839), .A2(n586), .B1(n14707), .B2(n587), .ZN(n11958)
         );
  OAI22_X1 U3282 ( .A1(n8823), .A2(n586), .B1(n14667), .B2(n587), .ZN(n11959)
         );
  OAI22_X1 U3283 ( .A1(n8807), .A2(n588), .B1(n14961), .B2(n589), .ZN(n11960)
         );
  OAI22_X1 U3284 ( .A1(n8791), .A2(n588), .B1(n14908), .B2(n589), .ZN(n11961)
         );
  OAI22_X1 U3285 ( .A1(n8775), .A2(n588), .B1(n14868), .B2(n589), .ZN(n11962)
         );
  OAI22_X1 U3286 ( .A1(n8759), .A2(n588), .B1(n14828), .B2(n589), .ZN(n11963)
         );
  OAI22_X1 U3287 ( .A1(n8743), .A2(n588), .B1(n14788), .B2(n589), .ZN(n11964)
         );
  OAI22_X1 U3288 ( .A1(n8727), .A2(n588), .B1(n14748), .B2(n589), .ZN(n11965)
         );
  OAI22_X1 U3289 ( .A1(n8711), .A2(n588), .B1(n14708), .B2(n589), .ZN(n11966)
         );
  OAI22_X1 U3290 ( .A1(n8695), .A2(n588), .B1(n14668), .B2(n589), .ZN(n11967)
         );
  OAI22_X1 U3291 ( .A1(n8679), .A2(n590), .B1(n14961), .B2(n591), .ZN(n11968)
         );
  OAI22_X1 U3292 ( .A1(n8663), .A2(n590), .B1(n14908), .B2(n591), .ZN(n11969)
         );
  OAI22_X1 U3293 ( .A1(n8647), .A2(n590), .B1(n14868), .B2(n591), .ZN(n11970)
         );
  OAI22_X1 U3294 ( .A1(n8631), .A2(n590), .B1(n14828), .B2(n591), .ZN(n11971)
         );
  OAI22_X1 U3295 ( .A1(n8615), .A2(n590), .B1(n14788), .B2(n591), .ZN(n11972)
         );
  OAI22_X1 U3296 ( .A1(n8599), .A2(n590), .B1(n14748), .B2(n591), .ZN(n11973)
         );
  OAI22_X1 U3297 ( .A1(n8583), .A2(n590), .B1(n14708), .B2(n591), .ZN(n11974)
         );
  OAI22_X1 U3298 ( .A1(n8567), .A2(n590), .B1(n14668), .B2(n591), .ZN(n11975)
         );
  OAI22_X1 U3299 ( .A1(n8551), .A2(n592), .B1(n14960), .B2(n593), .ZN(n11976)
         );
  OAI22_X1 U3300 ( .A1(n8535), .A2(n592), .B1(n14908), .B2(n593), .ZN(n11977)
         );
  OAI22_X1 U3301 ( .A1(n8519), .A2(n592), .B1(n14868), .B2(n593), .ZN(n11978)
         );
  OAI22_X1 U3302 ( .A1(n8503), .A2(n592), .B1(n14828), .B2(n593), .ZN(n11979)
         );
  OAI22_X1 U3303 ( .A1(n8487), .A2(n592), .B1(n14788), .B2(n593), .ZN(n11980)
         );
  OAI22_X1 U3304 ( .A1(n8471), .A2(n592), .B1(n14748), .B2(n593), .ZN(n11981)
         );
  OAI22_X1 U3305 ( .A1(n8455), .A2(n592), .B1(n14708), .B2(n593), .ZN(n11982)
         );
  OAI22_X1 U3306 ( .A1(n8439), .A2(n592), .B1(n14668), .B2(n593), .ZN(n11983)
         );
  OAI22_X1 U3307 ( .A1(n8423), .A2(n594), .B1(n14960), .B2(n595), .ZN(n11984)
         );
  OAI22_X1 U3308 ( .A1(n8407), .A2(n594), .B1(n14908), .B2(n595), .ZN(n11985)
         );
  OAI22_X1 U3309 ( .A1(n8391), .A2(n594), .B1(n14868), .B2(n595), .ZN(n11986)
         );
  OAI22_X1 U3310 ( .A1(n8375), .A2(n594), .B1(n14828), .B2(n595), .ZN(n11987)
         );
  OAI22_X1 U3311 ( .A1(n8359), .A2(n594), .B1(n14788), .B2(n595), .ZN(n11988)
         );
  OAI22_X1 U3312 ( .A1(n8343), .A2(n594), .B1(n14748), .B2(n595), .ZN(n11989)
         );
  OAI22_X1 U3313 ( .A1(n8327), .A2(n594), .B1(n14708), .B2(n595), .ZN(n11990)
         );
  OAI22_X1 U3314 ( .A1(n8311), .A2(n594), .B1(n14668), .B2(n595), .ZN(n11991)
         );
  OAI22_X1 U3315 ( .A1(n8295), .A2(n596), .B1(n14960), .B2(n597), .ZN(n11992)
         );
  OAI22_X1 U3316 ( .A1(n8279), .A2(n596), .B1(n14908), .B2(n597), .ZN(n11993)
         );
  OAI22_X1 U3317 ( .A1(n8263), .A2(n596), .B1(n14868), .B2(n597), .ZN(n11994)
         );
  OAI22_X1 U3318 ( .A1(n8247), .A2(n596), .B1(n14828), .B2(n597), .ZN(n11995)
         );
  OAI22_X1 U3319 ( .A1(n8231), .A2(n596), .B1(n14788), .B2(n597), .ZN(n11996)
         );
  OAI22_X1 U3320 ( .A1(n8215), .A2(n596), .B1(n14748), .B2(n597), .ZN(n11997)
         );
  OAI22_X1 U3321 ( .A1(n8199), .A2(n596), .B1(n14708), .B2(n597), .ZN(n11998)
         );
  OAI22_X1 U3322 ( .A1(n8183), .A2(n596), .B1(n14668), .B2(n597), .ZN(n11999)
         );
  OAI22_X1 U3323 ( .A1(n8167), .A2(n598), .B1(n14960), .B2(n599), .ZN(n12000)
         );
  OAI22_X1 U3324 ( .A1(n8151), .A2(n598), .B1(n14908), .B2(n599), .ZN(n12001)
         );
  OAI22_X1 U3325 ( .A1(n8135), .A2(n598), .B1(n14868), .B2(n599), .ZN(n12002)
         );
  OAI22_X1 U3326 ( .A1(n8119), .A2(n598), .B1(n14828), .B2(n599), .ZN(n12003)
         );
  OAI22_X1 U3327 ( .A1(n8103), .A2(n598), .B1(n14788), .B2(n599), .ZN(n12004)
         );
  OAI22_X1 U3328 ( .A1(n8087), .A2(n598), .B1(n14748), .B2(n599), .ZN(n12005)
         );
  OAI22_X1 U3329 ( .A1(n8071), .A2(n598), .B1(n14708), .B2(n599), .ZN(n12006)
         );
  OAI22_X1 U3330 ( .A1(n8055), .A2(n598), .B1(n14668), .B2(n599), .ZN(n12007)
         );
  OAI22_X1 U3331 ( .A1(n8039), .A2(n600), .B1(n14960), .B2(n601), .ZN(n12008)
         );
  OAI22_X1 U3332 ( .A1(n8023), .A2(n600), .B1(n14908), .B2(n601), .ZN(n12009)
         );
  OAI22_X1 U3333 ( .A1(n8007), .A2(n600), .B1(n14868), .B2(n601), .ZN(n12010)
         );
  OAI22_X1 U3334 ( .A1(n7991), .A2(n600), .B1(n14828), .B2(n601), .ZN(n12011)
         );
  OAI22_X1 U3335 ( .A1(n7975), .A2(n600), .B1(n14788), .B2(n601), .ZN(n12012)
         );
  OAI22_X1 U3336 ( .A1(n7959), .A2(n600), .B1(n14748), .B2(n601), .ZN(n12013)
         );
  OAI22_X1 U3337 ( .A1(n7943), .A2(n600), .B1(n14708), .B2(n601), .ZN(n12014)
         );
  OAI22_X1 U3338 ( .A1(n7927), .A2(n600), .B1(n14668), .B2(n601), .ZN(n12015)
         );
  OAI22_X1 U3339 ( .A1(n7911), .A2(n602), .B1(n14960), .B2(n603), .ZN(n12016)
         );
  OAI22_X1 U3340 ( .A1(n7895), .A2(n602), .B1(n14908), .B2(n603), .ZN(n12017)
         );
  OAI22_X1 U3341 ( .A1(n7879), .A2(n602), .B1(n14868), .B2(n603), .ZN(n12018)
         );
  OAI22_X1 U3342 ( .A1(n7863), .A2(n602), .B1(n14828), .B2(n603), .ZN(n12019)
         );
  OAI22_X1 U3343 ( .A1(n7847), .A2(n602), .B1(n14788), .B2(n603), .ZN(n12020)
         );
  OAI22_X1 U3344 ( .A1(n7831), .A2(n602), .B1(n14748), .B2(n603), .ZN(n12021)
         );
  OAI22_X1 U3345 ( .A1(n7815), .A2(n602), .B1(n14708), .B2(n603), .ZN(n12022)
         );
  OAI22_X1 U3346 ( .A1(n7799), .A2(n602), .B1(n14668), .B2(n603), .ZN(n12023)
         );
  OAI22_X1 U3347 ( .A1(n7783), .A2(n604), .B1(n14960), .B2(n605), .ZN(n12024)
         );
  OAI22_X1 U3348 ( .A1(n7767), .A2(n604), .B1(n14908), .B2(n605), .ZN(n12025)
         );
  OAI22_X1 U3349 ( .A1(n7751), .A2(n604), .B1(n14868), .B2(n605), .ZN(n12026)
         );
  OAI22_X1 U3350 ( .A1(n7735), .A2(n604), .B1(n14828), .B2(n605), .ZN(n12027)
         );
  OAI22_X1 U3351 ( .A1(n7719), .A2(n604), .B1(n14788), .B2(n605), .ZN(n12028)
         );
  OAI22_X1 U3352 ( .A1(n7703), .A2(n604), .B1(n14748), .B2(n605), .ZN(n12029)
         );
  OAI22_X1 U3353 ( .A1(n7687), .A2(n604), .B1(n14708), .B2(n605), .ZN(n12030)
         );
  OAI22_X1 U3354 ( .A1(n7671), .A2(n604), .B1(n14668), .B2(n605), .ZN(n12031)
         );
  OAI22_X1 U3355 ( .A1(n7655), .A2(n606), .B1(n14960), .B2(n607), .ZN(n12032)
         );
  OAI22_X1 U3356 ( .A1(n7639), .A2(n606), .B1(n14908), .B2(n607), .ZN(n12033)
         );
  OAI22_X1 U3357 ( .A1(n7623), .A2(n606), .B1(n14868), .B2(n607), .ZN(n12034)
         );
  OAI22_X1 U3358 ( .A1(n7607), .A2(n606), .B1(n14828), .B2(n607), .ZN(n12035)
         );
  OAI22_X1 U3359 ( .A1(n7591), .A2(n606), .B1(n14788), .B2(n607), .ZN(n12036)
         );
  OAI22_X1 U3360 ( .A1(n7575), .A2(n606), .B1(n14748), .B2(n607), .ZN(n12037)
         );
  OAI22_X1 U3361 ( .A1(n7559), .A2(n606), .B1(n14708), .B2(n607), .ZN(n12038)
         );
  OAI22_X1 U3362 ( .A1(n7543), .A2(n606), .B1(n14668), .B2(n607), .ZN(n12039)
         );
  OAI22_X1 U3363 ( .A1(n7527), .A2(n608), .B1(n14960), .B2(n609), .ZN(n12040)
         );
  OAI22_X1 U3364 ( .A1(n7511), .A2(n608), .B1(n14908), .B2(n609), .ZN(n12041)
         );
  OAI22_X1 U3365 ( .A1(n7495), .A2(n608), .B1(n14868), .B2(n609), .ZN(n12042)
         );
  OAI22_X1 U3366 ( .A1(n7479), .A2(n608), .B1(n14828), .B2(n609), .ZN(n12043)
         );
  OAI22_X1 U3367 ( .A1(n7463), .A2(n608), .B1(n14788), .B2(n609), .ZN(n12044)
         );
  OAI22_X1 U3368 ( .A1(n7447), .A2(n608), .B1(n14748), .B2(n609), .ZN(n12045)
         );
  OAI22_X1 U3369 ( .A1(n7431), .A2(n608), .B1(n14708), .B2(n609), .ZN(n12046)
         );
  OAI22_X1 U3370 ( .A1(n7415), .A2(n608), .B1(n14668), .B2(n609), .ZN(n12047)
         );
  OAI22_X1 U3371 ( .A1(n7399), .A2(n610), .B1(n14960), .B2(n611), .ZN(n12048)
         );
  OAI22_X1 U3372 ( .A1(n7383), .A2(n610), .B1(n14908), .B2(n611), .ZN(n12049)
         );
  OAI22_X1 U3373 ( .A1(n7367), .A2(n610), .B1(n14868), .B2(n611), .ZN(n12050)
         );
  OAI22_X1 U3374 ( .A1(n7351), .A2(n610), .B1(n14828), .B2(n611), .ZN(n12051)
         );
  OAI22_X1 U3375 ( .A1(n7335), .A2(n610), .B1(n14788), .B2(n611), .ZN(n12052)
         );
  OAI22_X1 U3376 ( .A1(n7319), .A2(n610), .B1(n14748), .B2(n611), .ZN(n12053)
         );
  OAI22_X1 U3377 ( .A1(n7303), .A2(n610), .B1(n14708), .B2(n611), .ZN(n12054)
         );
  OAI22_X1 U3378 ( .A1(n7287), .A2(n610), .B1(n14668), .B2(n611), .ZN(n12055)
         );
  OAI22_X1 U3379 ( .A1(n7271), .A2(n612), .B1(n14960), .B2(n613), .ZN(n12056)
         );
  OAI22_X1 U3380 ( .A1(n7255), .A2(n612), .B1(n14908), .B2(n613), .ZN(n12057)
         );
  OAI22_X1 U3381 ( .A1(n7239), .A2(n612), .B1(n14868), .B2(n613), .ZN(n12058)
         );
  OAI22_X1 U3382 ( .A1(n7223), .A2(n612), .B1(n14828), .B2(n613), .ZN(n12059)
         );
  OAI22_X1 U3383 ( .A1(n7207), .A2(n612), .B1(n14788), .B2(n613), .ZN(n12060)
         );
  OAI22_X1 U3384 ( .A1(n7191), .A2(n612), .B1(n14748), .B2(n613), .ZN(n12061)
         );
  OAI22_X1 U3385 ( .A1(n7175), .A2(n612), .B1(n14708), .B2(n613), .ZN(n12062)
         );
  OAI22_X1 U3386 ( .A1(n7159), .A2(n612), .B1(n14668), .B2(n613), .ZN(n12063)
         );
  OAI22_X1 U3387 ( .A1(n7143), .A2(n614), .B1(n14960), .B2(n615), .ZN(n12064)
         );
  OAI22_X1 U3388 ( .A1(n7127), .A2(n614), .B1(n14909), .B2(n615), .ZN(n12065)
         );
  OAI22_X1 U3389 ( .A1(n7111), .A2(n614), .B1(n14869), .B2(n615), .ZN(n12066)
         );
  OAI22_X1 U3390 ( .A1(n7095), .A2(n614), .B1(n14829), .B2(n615), .ZN(n12067)
         );
  OAI22_X1 U3391 ( .A1(n7079), .A2(n614), .B1(n14789), .B2(n615), .ZN(n12068)
         );
  OAI22_X1 U3392 ( .A1(n7063), .A2(n614), .B1(n14749), .B2(n615), .ZN(n12069)
         );
  OAI22_X1 U3393 ( .A1(n7047), .A2(n614), .B1(n14709), .B2(n615), .ZN(n12070)
         );
  OAI22_X1 U3394 ( .A1(n7031), .A2(n614), .B1(n14669), .B2(n615), .ZN(n12071)
         );
  OAI22_X1 U3395 ( .A1(n7015), .A2(n616), .B1(n14960), .B2(n617), .ZN(n12072)
         );
  OAI22_X1 U3396 ( .A1(n6999), .A2(n616), .B1(n14909), .B2(n617), .ZN(n12073)
         );
  OAI22_X1 U3397 ( .A1(n6983), .A2(n616), .B1(n14869), .B2(n617), .ZN(n12074)
         );
  OAI22_X1 U3398 ( .A1(n6967), .A2(n616), .B1(n14829), .B2(n617), .ZN(n12075)
         );
  OAI22_X1 U3399 ( .A1(n6951), .A2(n616), .B1(n14789), .B2(n617), .ZN(n12076)
         );
  OAI22_X1 U3400 ( .A1(n6935), .A2(n616), .B1(n14749), .B2(n617), .ZN(n12077)
         );
  OAI22_X1 U3401 ( .A1(n6919), .A2(n616), .B1(n14709), .B2(n617), .ZN(n12078)
         );
  OAI22_X1 U3402 ( .A1(n6903), .A2(n616), .B1(n14669), .B2(n617), .ZN(n12079)
         );
  OAI22_X1 U3403 ( .A1(n6887), .A2(n618), .B1(n14959), .B2(n619), .ZN(n12080)
         );
  OAI22_X1 U3404 ( .A1(n6871), .A2(n618), .B1(n14909), .B2(n619), .ZN(n12081)
         );
  OAI22_X1 U3405 ( .A1(n6855), .A2(n618), .B1(n14869), .B2(n619), .ZN(n12082)
         );
  OAI22_X1 U3406 ( .A1(n6839), .A2(n618), .B1(n14829), .B2(n619), .ZN(n12083)
         );
  OAI22_X1 U3407 ( .A1(n6823), .A2(n618), .B1(n14789), .B2(n619), .ZN(n12084)
         );
  OAI22_X1 U3408 ( .A1(n6807), .A2(n618), .B1(n14749), .B2(n619), .ZN(n12085)
         );
  OAI22_X1 U3409 ( .A1(n6791), .A2(n618), .B1(n14709), .B2(n619), .ZN(n12086)
         );
  OAI22_X1 U3410 ( .A1(n6775), .A2(n618), .B1(n14669), .B2(n619), .ZN(n12087)
         );
  OAI22_X1 U3411 ( .A1(n6759), .A2(n620), .B1(n14959), .B2(n621), .ZN(n12088)
         );
  OAI22_X1 U3412 ( .A1(n6743), .A2(n620), .B1(n14909), .B2(n621), .ZN(n12089)
         );
  OAI22_X1 U3413 ( .A1(n6727), .A2(n620), .B1(n14869), .B2(n621), .ZN(n12090)
         );
  OAI22_X1 U3414 ( .A1(n6711), .A2(n620), .B1(n14829), .B2(n621), .ZN(n12091)
         );
  OAI22_X1 U3415 ( .A1(n6695), .A2(n620), .B1(n14789), .B2(n621), .ZN(n12092)
         );
  OAI22_X1 U3416 ( .A1(n6679), .A2(n620), .B1(n14749), .B2(n621), .ZN(n12093)
         );
  OAI22_X1 U3417 ( .A1(n6663), .A2(n620), .B1(n14709), .B2(n621), .ZN(n12094)
         );
  OAI22_X1 U3418 ( .A1(n6647), .A2(n620), .B1(n14669), .B2(n621), .ZN(n12095)
         );
  OAI22_X1 U3419 ( .A1(n6631), .A2(n622), .B1(n14959), .B2(n623), .ZN(n12096)
         );
  OAI22_X1 U3420 ( .A1(n6615), .A2(n622), .B1(n14909), .B2(n623), .ZN(n12097)
         );
  OAI22_X1 U3421 ( .A1(n6599), .A2(n622), .B1(n14869), .B2(n623), .ZN(n12098)
         );
  OAI22_X1 U3422 ( .A1(n6583), .A2(n622), .B1(n14829), .B2(n623), .ZN(n12099)
         );
  OAI22_X1 U3423 ( .A1(n6567), .A2(n622), .B1(n14789), .B2(n623), .ZN(n12100)
         );
  OAI22_X1 U3424 ( .A1(n6551), .A2(n622), .B1(n14749), .B2(n623), .ZN(n12101)
         );
  OAI22_X1 U3425 ( .A1(n6535), .A2(n622), .B1(n14709), .B2(n623), .ZN(n12102)
         );
  OAI22_X1 U3426 ( .A1(n6519), .A2(n622), .B1(n14669), .B2(n623), .ZN(n12103)
         );
  OAI22_X1 U3427 ( .A1(n6503), .A2(n624), .B1(n14959), .B2(n625), .ZN(n12104)
         );
  OAI22_X1 U3428 ( .A1(n6487), .A2(n624), .B1(n14909), .B2(n625), .ZN(n12105)
         );
  OAI22_X1 U3429 ( .A1(n6471), .A2(n624), .B1(n14869), .B2(n625), .ZN(n12106)
         );
  OAI22_X1 U3430 ( .A1(n6455), .A2(n624), .B1(n14829), .B2(n625), .ZN(n12107)
         );
  OAI22_X1 U3431 ( .A1(n6439), .A2(n624), .B1(n14789), .B2(n625), .ZN(n12108)
         );
  OAI22_X1 U3432 ( .A1(n6423), .A2(n624), .B1(n14749), .B2(n625), .ZN(n12109)
         );
  OAI22_X1 U3433 ( .A1(n6407), .A2(n624), .B1(n14709), .B2(n625), .ZN(n12110)
         );
  OAI22_X1 U3434 ( .A1(n6391), .A2(n624), .B1(n14669), .B2(n625), .ZN(n12111)
         );
  OAI22_X1 U3435 ( .A1(n6375), .A2(n626), .B1(n14959), .B2(n627), .ZN(n12112)
         );
  OAI22_X1 U3436 ( .A1(n6359), .A2(n626), .B1(n14909), .B2(n627), .ZN(n12113)
         );
  OAI22_X1 U3437 ( .A1(n6343), .A2(n626), .B1(n14869), .B2(n627), .ZN(n12114)
         );
  OAI22_X1 U3438 ( .A1(n6327), .A2(n626), .B1(n14829), .B2(n627), .ZN(n12115)
         );
  OAI22_X1 U3439 ( .A1(n6311), .A2(n626), .B1(n14789), .B2(n627), .ZN(n12116)
         );
  OAI22_X1 U3440 ( .A1(n6295), .A2(n626), .B1(n14749), .B2(n627), .ZN(n12117)
         );
  OAI22_X1 U3441 ( .A1(n6279), .A2(n626), .B1(n14709), .B2(n627), .ZN(n12118)
         );
  OAI22_X1 U3442 ( .A1(n6263), .A2(n626), .B1(n14669), .B2(n627), .ZN(n12119)
         );
  OAI22_X1 U3443 ( .A1(n6247), .A2(n628), .B1(n14959), .B2(n629), .ZN(n12120)
         );
  OAI22_X1 U3444 ( .A1(n6231), .A2(n628), .B1(n14909), .B2(n629), .ZN(n12121)
         );
  OAI22_X1 U3445 ( .A1(n6215), .A2(n628), .B1(n14869), .B2(n629), .ZN(n12122)
         );
  OAI22_X1 U3446 ( .A1(n6199), .A2(n628), .B1(n14829), .B2(n629), .ZN(n12123)
         );
  OAI22_X1 U3447 ( .A1(n6183), .A2(n628), .B1(n14789), .B2(n629), .ZN(n12124)
         );
  OAI22_X1 U3448 ( .A1(n6167), .A2(n628), .B1(n14749), .B2(n629), .ZN(n12125)
         );
  OAI22_X1 U3449 ( .A1(n6151), .A2(n628), .B1(n14709), .B2(n629), .ZN(n12126)
         );
  OAI22_X1 U3450 ( .A1(n6135), .A2(n628), .B1(n14669), .B2(n629), .ZN(n12127)
         );
  OAI22_X1 U3451 ( .A1(n6119), .A2(n630), .B1(n14959), .B2(n631), .ZN(n12128)
         );
  OAI22_X1 U3452 ( .A1(n6103), .A2(n630), .B1(n14909), .B2(n631), .ZN(n12129)
         );
  OAI22_X1 U3453 ( .A1(n6087), .A2(n630), .B1(n14869), .B2(n631), .ZN(n12130)
         );
  OAI22_X1 U3454 ( .A1(n6071), .A2(n630), .B1(n14829), .B2(n631), .ZN(n12131)
         );
  OAI22_X1 U3455 ( .A1(n6055), .A2(n630), .B1(n14789), .B2(n631), .ZN(n12132)
         );
  OAI22_X1 U3456 ( .A1(n6039), .A2(n630), .B1(n14749), .B2(n631), .ZN(n12133)
         );
  OAI22_X1 U3457 ( .A1(n6023), .A2(n630), .B1(n14709), .B2(n631), .ZN(n12134)
         );
  OAI22_X1 U3458 ( .A1(n6007), .A2(n630), .B1(n14669), .B2(n631), .ZN(n12135)
         );
  OAI22_X1 U3459 ( .A1(n9314), .A2(n1039), .B1(n14944), .B2(n1040), .ZN(n13720) );
  OAI22_X1 U3460 ( .A1(n9298), .A2(n1039), .B1(n14924), .B2(n1040), .ZN(n13721) );
  OAI22_X1 U3461 ( .A1(n9282), .A2(n1039), .B1(n14884), .B2(n1040), .ZN(n13722) );
  OAI22_X1 U3462 ( .A1(n9266), .A2(n1039), .B1(n14844), .B2(n1040), .ZN(n13723) );
  OAI22_X1 U3463 ( .A1(n9250), .A2(n1039), .B1(n14804), .B2(n1040), .ZN(n13724) );
  OAI22_X1 U3464 ( .A1(n9234), .A2(n1039), .B1(n14764), .B2(n1040), .ZN(n13725) );
  OAI22_X1 U3465 ( .A1(n9218), .A2(n1039), .B1(n14724), .B2(n1040), .ZN(n13726) );
  OAI22_X1 U3466 ( .A1(n9202), .A2(n1039), .B1(n14684), .B2(n1040), .ZN(n13727) );
  OAI22_X1 U3467 ( .A1(n9186), .A2(n1041), .B1(n14944), .B2(n1042), .ZN(n13728) );
  OAI22_X1 U3468 ( .A1(n9170), .A2(n1041), .B1(n14925), .B2(n1042), .ZN(n13729) );
  OAI22_X1 U3469 ( .A1(n9154), .A2(n1041), .B1(n14885), .B2(n1042), .ZN(n13730) );
  OAI22_X1 U3470 ( .A1(n9138), .A2(n1041), .B1(n14845), .B2(n1042), .ZN(n13731) );
  OAI22_X1 U3471 ( .A1(n9122), .A2(n1041), .B1(n14805), .B2(n1042), .ZN(n13732) );
  OAI22_X1 U3472 ( .A1(n9106), .A2(n1041), .B1(n14765), .B2(n1042), .ZN(n13733) );
  OAI22_X1 U3473 ( .A1(n9090), .A2(n1041), .B1(n14725), .B2(n1042), .ZN(n13734) );
  OAI22_X1 U3474 ( .A1(n9074), .A2(n1041), .B1(n14685), .B2(n1042), .ZN(n13735) );
  OAI22_X1 U3475 ( .A1(n9058), .A2(n1043), .B1(n14944), .B2(n1044), .ZN(n13736) );
  OAI22_X1 U3476 ( .A1(n9042), .A2(n1043), .B1(n14925), .B2(n1044), .ZN(n13737) );
  OAI22_X1 U3477 ( .A1(n9026), .A2(n1043), .B1(n14885), .B2(n1044), .ZN(n13738) );
  OAI22_X1 U3478 ( .A1(n9010), .A2(n1043), .B1(n14845), .B2(n1044), .ZN(n13739) );
  OAI22_X1 U3479 ( .A1(n8994), .A2(n1043), .B1(n14805), .B2(n1044), .ZN(n13740) );
  OAI22_X1 U3480 ( .A1(n8978), .A2(n1043), .B1(n14765), .B2(n1044), .ZN(n13741) );
  OAI22_X1 U3481 ( .A1(n8962), .A2(n1043), .B1(n14725), .B2(n1044), .ZN(n13742) );
  OAI22_X1 U3482 ( .A1(n8946), .A2(n1043), .B1(n14685), .B2(n1044), .ZN(n13743) );
  OAI22_X1 U3483 ( .A1(n8930), .A2(n1045), .B1(n14943), .B2(n1046), .ZN(n13744) );
  OAI22_X1 U3484 ( .A1(n8914), .A2(n1045), .B1(n14925), .B2(n1046), .ZN(n13745) );
  OAI22_X1 U3485 ( .A1(n8898), .A2(n1045), .B1(n14885), .B2(n1046), .ZN(n13746) );
  OAI22_X1 U3486 ( .A1(n8882), .A2(n1045), .B1(n14845), .B2(n1046), .ZN(n13747) );
  OAI22_X1 U3487 ( .A1(n8866), .A2(n1045), .B1(n14805), .B2(n1046), .ZN(n13748) );
  OAI22_X1 U3488 ( .A1(n8850), .A2(n1045), .B1(n14765), .B2(n1046), .ZN(n13749) );
  OAI22_X1 U3489 ( .A1(n8834), .A2(n1045), .B1(n14725), .B2(n1046), .ZN(n13750) );
  OAI22_X1 U3490 ( .A1(n8818), .A2(n1045), .B1(n14685), .B2(n1046), .ZN(n13751) );
  OAI22_X1 U3491 ( .A1(n8802), .A2(n1047), .B1(n14943), .B2(n1048), .ZN(n13752) );
  OAI22_X1 U3492 ( .A1(n8786), .A2(n1047), .B1(n14925), .B2(n1048), .ZN(n13753) );
  OAI22_X1 U3493 ( .A1(n8770), .A2(n1047), .B1(n14885), .B2(n1048), .ZN(n13754) );
  OAI22_X1 U3494 ( .A1(n8754), .A2(n1047), .B1(n14845), .B2(n1048), .ZN(n13755) );
  OAI22_X1 U3495 ( .A1(n8738), .A2(n1047), .B1(n14805), .B2(n1048), .ZN(n13756) );
  OAI22_X1 U3496 ( .A1(n8722), .A2(n1047), .B1(n14765), .B2(n1048), .ZN(n13757) );
  OAI22_X1 U3497 ( .A1(n8706), .A2(n1047), .B1(n14725), .B2(n1048), .ZN(n13758) );
  OAI22_X1 U3498 ( .A1(n8690), .A2(n1047), .B1(n14685), .B2(n1048), .ZN(n13759) );
  OAI22_X1 U3499 ( .A1(n8674), .A2(n1049), .B1(n14943), .B2(n1050), .ZN(n13760) );
  OAI22_X1 U3500 ( .A1(n8658), .A2(n1049), .B1(n14925), .B2(n1050), .ZN(n13761) );
  OAI22_X1 U3501 ( .A1(n8642), .A2(n1049), .B1(n14885), .B2(n1050), .ZN(n13762) );
  OAI22_X1 U3502 ( .A1(n8626), .A2(n1049), .B1(n14845), .B2(n1050), .ZN(n13763) );
  OAI22_X1 U3503 ( .A1(n8610), .A2(n1049), .B1(n14805), .B2(n1050), .ZN(n13764) );
  OAI22_X1 U3504 ( .A1(n8594), .A2(n1049), .B1(n14765), .B2(n1050), .ZN(n13765) );
  OAI22_X1 U3505 ( .A1(n8578), .A2(n1049), .B1(n14725), .B2(n1050), .ZN(n13766) );
  OAI22_X1 U3506 ( .A1(n8562), .A2(n1049), .B1(n14685), .B2(n1050), .ZN(n13767) );
  OAI22_X1 U3507 ( .A1(n8546), .A2(n1051), .B1(n14943), .B2(n1052), .ZN(n13768) );
  OAI22_X1 U3508 ( .A1(n8530), .A2(n1051), .B1(n14925), .B2(n1052), .ZN(n13769) );
  OAI22_X1 U3509 ( .A1(n8514), .A2(n1051), .B1(n14885), .B2(n1052), .ZN(n13770) );
  OAI22_X1 U3510 ( .A1(n8498), .A2(n1051), .B1(n14845), .B2(n1052), .ZN(n13771) );
  OAI22_X1 U3511 ( .A1(n8482), .A2(n1051), .B1(n14805), .B2(n1052), .ZN(n13772) );
  OAI22_X1 U3512 ( .A1(n8466), .A2(n1051), .B1(n14765), .B2(n1052), .ZN(n13773) );
  OAI22_X1 U3513 ( .A1(n8450), .A2(n1051), .B1(n14725), .B2(n1052), .ZN(n13774) );
  OAI22_X1 U3514 ( .A1(n8434), .A2(n1051), .B1(n14685), .B2(n1052), .ZN(n13775) );
  OAI22_X1 U3515 ( .A1(n8418), .A2(n1053), .B1(n14943), .B2(n1054), .ZN(n13776) );
  OAI22_X1 U3516 ( .A1(n8402), .A2(n1053), .B1(n14925), .B2(n1054), .ZN(n13777) );
  OAI22_X1 U3517 ( .A1(n8386), .A2(n1053), .B1(n14885), .B2(n1054), .ZN(n13778) );
  OAI22_X1 U3518 ( .A1(n8370), .A2(n1053), .B1(n14845), .B2(n1054), .ZN(n13779) );
  OAI22_X1 U3519 ( .A1(n8354), .A2(n1053), .B1(n14805), .B2(n1054), .ZN(n13780) );
  OAI22_X1 U3520 ( .A1(n8338), .A2(n1053), .B1(n14765), .B2(n1054), .ZN(n13781) );
  OAI22_X1 U3521 ( .A1(n8322), .A2(n1053), .B1(n14725), .B2(n1054), .ZN(n13782) );
  OAI22_X1 U3522 ( .A1(n8306), .A2(n1053), .B1(n14685), .B2(n1054), .ZN(n13783) );
  OAI22_X1 U3523 ( .A1(n8290), .A2(n1055), .B1(n14943), .B2(n1056), .ZN(n13784) );
  OAI22_X1 U3524 ( .A1(n8274), .A2(n1055), .B1(n14925), .B2(n1056), .ZN(n13785) );
  OAI22_X1 U3525 ( .A1(n8258), .A2(n1055), .B1(n14885), .B2(n1056), .ZN(n13786) );
  OAI22_X1 U3526 ( .A1(n8242), .A2(n1055), .B1(n14845), .B2(n1056), .ZN(n13787) );
  OAI22_X1 U3527 ( .A1(n8226), .A2(n1055), .B1(n14805), .B2(n1056), .ZN(n13788) );
  OAI22_X1 U3528 ( .A1(n8210), .A2(n1055), .B1(n14765), .B2(n1056), .ZN(n13789) );
  OAI22_X1 U3529 ( .A1(n8194), .A2(n1055), .B1(n14725), .B2(n1056), .ZN(n13790) );
  OAI22_X1 U3530 ( .A1(n8178), .A2(n1055), .B1(n14685), .B2(n1056), .ZN(n13791) );
  OAI22_X1 U3531 ( .A1(n8162), .A2(n1057), .B1(n14943), .B2(n1058), .ZN(n13792) );
  OAI22_X1 U3532 ( .A1(n8146), .A2(n1057), .B1(n14925), .B2(n1058), .ZN(n13793) );
  OAI22_X1 U3533 ( .A1(n8130), .A2(n1057), .B1(n14885), .B2(n1058), .ZN(n13794) );
  OAI22_X1 U3534 ( .A1(n8114), .A2(n1057), .B1(n14845), .B2(n1058), .ZN(n13795) );
  OAI22_X1 U3535 ( .A1(n8098), .A2(n1057), .B1(n14805), .B2(n1058), .ZN(n13796) );
  OAI22_X1 U3536 ( .A1(n8082), .A2(n1057), .B1(n14765), .B2(n1058), .ZN(n13797) );
  OAI22_X1 U3537 ( .A1(n8066), .A2(n1057), .B1(n14725), .B2(n1058), .ZN(n13798) );
  OAI22_X1 U3538 ( .A1(n8050), .A2(n1057), .B1(n14685), .B2(n1058), .ZN(n13799) );
  OAI22_X1 U3539 ( .A1(n8034), .A2(n1059), .B1(n14943), .B2(n1060), .ZN(n13800) );
  OAI22_X1 U3540 ( .A1(n8018), .A2(n1059), .B1(n14925), .B2(n1060), .ZN(n13801) );
  OAI22_X1 U3541 ( .A1(n8002), .A2(n1059), .B1(n14885), .B2(n1060), .ZN(n13802) );
  OAI22_X1 U3542 ( .A1(n7986), .A2(n1059), .B1(n14845), .B2(n1060), .ZN(n13803) );
  OAI22_X1 U3543 ( .A1(n7970), .A2(n1059), .B1(n14805), .B2(n1060), .ZN(n13804) );
  OAI22_X1 U3544 ( .A1(n7954), .A2(n1059), .B1(n14765), .B2(n1060), .ZN(n13805) );
  OAI22_X1 U3545 ( .A1(n7938), .A2(n1059), .B1(n14725), .B2(n1060), .ZN(n13806) );
  OAI22_X1 U3546 ( .A1(n7922), .A2(n1059), .B1(n14685), .B2(n1060), .ZN(n13807) );
  OAI22_X1 U3547 ( .A1(n7906), .A2(n1061), .B1(n14943), .B2(n1062), .ZN(n13808) );
  OAI22_X1 U3548 ( .A1(n7890), .A2(n1061), .B1(n14925), .B2(n1062), .ZN(n13809) );
  OAI22_X1 U3549 ( .A1(n7874), .A2(n1061), .B1(n14885), .B2(n1062), .ZN(n13810) );
  OAI22_X1 U3550 ( .A1(n7858), .A2(n1061), .B1(n14845), .B2(n1062), .ZN(n13811) );
  OAI22_X1 U3551 ( .A1(n7842), .A2(n1061), .B1(n14805), .B2(n1062), .ZN(n13812) );
  OAI22_X1 U3552 ( .A1(n7826), .A2(n1061), .B1(n14765), .B2(n1062), .ZN(n13813) );
  OAI22_X1 U3553 ( .A1(n7810), .A2(n1061), .B1(n14725), .B2(n1062), .ZN(n13814) );
  OAI22_X1 U3554 ( .A1(n7794), .A2(n1061), .B1(n14685), .B2(n1062), .ZN(n13815) );
  OAI22_X1 U3555 ( .A1(n7778), .A2(n1063), .B1(n14943), .B2(n1064), .ZN(n13816) );
  OAI22_X1 U3556 ( .A1(n7762), .A2(n1063), .B1(n14925), .B2(n1064), .ZN(n13817) );
  OAI22_X1 U3557 ( .A1(n7746), .A2(n1063), .B1(n14885), .B2(n1064), .ZN(n13818) );
  OAI22_X1 U3558 ( .A1(n7730), .A2(n1063), .B1(n14845), .B2(n1064), .ZN(n13819) );
  OAI22_X1 U3559 ( .A1(n7714), .A2(n1063), .B1(n14805), .B2(n1064), .ZN(n13820) );
  OAI22_X1 U3560 ( .A1(n7698), .A2(n1063), .B1(n14765), .B2(n1064), .ZN(n13821) );
  OAI22_X1 U3561 ( .A1(n7682), .A2(n1063), .B1(n14725), .B2(n1064), .ZN(n13822) );
  OAI22_X1 U3562 ( .A1(n7666), .A2(n1063), .B1(n14685), .B2(n1064), .ZN(n13823) );
  OAI22_X1 U3563 ( .A1(n7650), .A2(n1065), .B1(n14943), .B2(n1066), .ZN(n13824) );
  OAI22_X1 U3564 ( .A1(n7634), .A2(n1065), .B1(n14925), .B2(n1066), .ZN(n13825) );
  OAI22_X1 U3565 ( .A1(n7618), .A2(n1065), .B1(n14885), .B2(n1066), .ZN(n13826) );
  OAI22_X1 U3566 ( .A1(n7602), .A2(n1065), .B1(n14845), .B2(n1066), .ZN(n13827) );
  OAI22_X1 U3567 ( .A1(n7586), .A2(n1065), .B1(n14805), .B2(n1066), .ZN(n13828) );
  OAI22_X1 U3568 ( .A1(n7570), .A2(n1065), .B1(n14765), .B2(n1066), .ZN(n13829) );
  OAI22_X1 U3569 ( .A1(n7554), .A2(n1065), .B1(n14725), .B2(n1066), .ZN(n13830) );
  OAI22_X1 U3570 ( .A1(n7538), .A2(n1065), .B1(n14685), .B2(n1066), .ZN(n13831) );
  OAI22_X1 U3571 ( .A1(n7522), .A2(n1067), .B1(n14943), .B2(n1068), .ZN(n13832) );
  OAI22_X1 U3572 ( .A1(n7506), .A2(n1067), .B1(n14926), .B2(n1068), .ZN(n13833) );
  OAI22_X1 U3573 ( .A1(n7490), .A2(n1067), .B1(n14886), .B2(n1068), .ZN(n13834) );
  OAI22_X1 U3574 ( .A1(n7474), .A2(n1067), .B1(n14846), .B2(n1068), .ZN(n13835) );
  OAI22_X1 U3575 ( .A1(n7458), .A2(n1067), .B1(n14806), .B2(n1068), .ZN(n13836) );
  OAI22_X1 U3576 ( .A1(n7442), .A2(n1067), .B1(n14766), .B2(n1068), .ZN(n13837) );
  OAI22_X1 U3577 ( .A1(n7426), .A2(n1067), .B1(n14726), .B2(n1068), .ZN(n13838) );
  OAI22_X1 U3578 ( .A1(n7410), .A2(n1067), .B1(n14686), .B2(n1068), .ZN(n13839) );
  OAI22_X1 U3579 ( .A1(n7394), .A2(n1069), .B1(n14943), .B2(n1070), .ZN(n13840) );
  OAI22_X1 U3580 ( .A1(n7378), .A2(n1069), .B1(n14926), .B2(n1070), .ZN(n13841) );
  OAI22_X1 U3581 ( .A1(n7362), .A2(n1069), .B1(n14886), .B2(n1070), .ZN(n13842) );
  OAI22_X1 U3582 ( .A1(n7346), .A2(n1069), .B1(n14846), .B2(n1070), .ZN(n13843) );
  OAI22_X1 U3583 ( .A1(n7330), .A2(n1069), .B1(n14806), .B2(n1070), .ZN(n13844) );
  OAI22_X1 U3584 ( .A1(n7314), .A2(n1069), .B1(n14766), .B2(n1070), .ZN(n13845) );
  OAI22_X1 U3585 ( .A1(n7298), .A2(n1069), .B1(n14726), .B2(n1070), .ZN(n13846) );
  OAI22_X1 U3586 ( .A1(n7282), .A2(n1069), .B1(n14686), .B2(n1070), .ZN(n13847) );
  OAI22_X1 U3587 ( .A1(n7266), .A2(n1071), .B1(n14942), .B2(n1072), .ZN(n13848) );
  OAI22_X1 U3588 ( .A1(n7250), .A2(n1071), .B1(n14926), .B2(n1072), .ZN(n13849) );
  OAI22_X1 U3589 ( .A1(n7234), .A2(n1071), .B1(n14886), .B2(n1072), .ZN(n13850) );
  OAI22_X1 U3590 ( .A1(n7218), .A2(n1071), .B1(n14846), .B2(n1072), .ZN(n13851) );
  OAI22_X1 U3591 ( .A1(n7202), .A2(n1071), .B1(n14806), .B2(n1072), .ZN(n13852) );
  OAI22_X1 U3592 ( .A1(n7186), .A2(n1071), .B1(n14766), .B2(n1072), .ZN(n13853) );
  OAI22_X1 U3593 ( .A1(n7170), .A2(n1071), .B1(n14726), .B2(n1072), .ZN(n13854) );
  OAI22_X1 U3594 ( .A1(n7154), .A2(n1071), .B1(n14686), .B2(n1072), .ZN(n13855) );
  OAI22_X1 U3595 ( .A1(n7138), .A2(n1073), .B1(n14942), .B2(n1074), .ZN(n13856) );
  OAI22_X1 U3596 ( .A1(n7122), .A2(n1073), .B1(n14926), .B2(n1074), .ZN(n13857) );
  OAI22_X1 U3597 ( .A1(n7106), .A2(n1073), .B1(n14886), .B2(n1074), .ZN(n13858) );
  OAI22_X1 U3598 ( .A1(n7090), .A2(n1073), .B1(n14846), .B2(n1074), .ZN(n13859) );
  OAI22_X1 U3599 ( .A1(n7074), .A2(n1073), .B1(n14806), .B2(n1074), .ZN(n13860) );
  OAI22_X1 U3600 ( .A1(n7058), .A2(n1073), .B1(n14766), .B2(n1074), .ZN(n13861) );
  OAI22_X1 U3601 ( .A1(n7042), .A2(n1073), .B1(n14726), .B2(n1074), .ZN(n13862) );
  OAI22_X1 U3602 ( .A1(n7026), .A2(n1073), .B1(n14686), .B2(n1074), .ZN(n13863) );
  OAI22_X1 U3603 ( .A1(n7010), .A2(n1075), .B1(n14942), .B2(n1076), .ZN(n13864) );
  OAI22_X1 U3604 ( .A1(n6994), .A2(n1075), .B1(n14926), .B2(n1076), .ZN(n13865) );
  OAI22_X1 U3605 ( .A1(n6978), .A2(n1075), .B1(n14886), .B2(n1076), .ZN(n13866) );
  OAI22_X1 U3606 ( .A1(n6962), .A2(n1075), .B1(n14846), .B2(n1076), .ZN(n13867) );
  OAI22_X1 U3607 ( .A1(n6946), .A2(n1075), .B1(n14806), .B2(n1076), .ZN(n13868) );
  OAI22_X1 U3608 ( .A1(n6930), .A2(n1075), .B1(n14766), .B2(n1076), .ZN(n13869) );
  OAI22_X1 U3609 ( .A1(n6914), .A2(n1075), .B1(n14726), .B2(n1076), .ZN(n13870) );
  OAI22_X1 U3610 ( .A1(n6898), .A2(n1075), .B1(n14686), .B2(n1076), .ZN(n13871) );
  OAI22_X1 U3611 ( .A1(n6882), .A2(n1077), .B1(n14942), .B2(n1078), .ZN(n13872) );
  OAI22_X1 U3612 ( .A1(n6866), .A2(n1077), .B1(n14926), .B2(n1078), .ZN(n13873) );
  OAI22_X1 U3613 ( .A1(n6850), .A2(n1077), .B1(n14886), .B2(n1078), .ZN(n13874) );
  OAI22_X1 U3614 ( .A1(n6834), .A2(n1077), .B1(n14846), .B2(n1078), .ZN(n13875) );
  OAI22_X1 U3615 ( .A1(n6818), .A2(n1077), .B1(n14806), .B2(n1078), .ZN(n13876) );
  OAI22_X1 U3616 ( .A1(n6802), .A2(n1077), .B1(n14766), .B2(n1078), .ZN(n13877) );
  OAI22_X1 U3617 ( .A1(n6786), .A2(n1077), .B1(n14726), .B2(n1078), .ZN(n13878) );
  OAI22_X1 U3618 ( .A1(n6770), .A2(n1077), .B1(n14686), .B2(n1078), .ZN(n13879) );
  OAI22_X1 U3619 ( .A1(n6754), .A2(n1079), .B1(n14942), .B2(n1080), .ZN(n13880) );
  OAI22_X1 U3620 ( .A1(n6738), .A2(n1079), .B1(n14926), .B2(n1080), .ZN(n13881) );
  OAI22_X1 U3621 ( .A1(n6722), .A2(n1079), .B1(n14886), .B2(n1080), .ZN(n13882) );
  OAI22_X1 U3622 ( .A1(n6706), .A2(n1079), .B1(n14846), .B2(n1080), .ZN(n13883) );
  OAI22_X1 U3623 ( .A1(n6690), .A2(n1079), .B1(n14806), .B2(n1080), .ZN(n13884) );
  OAI22_X1 U3624 ( .A1(n6674), .A2(n1079), .B1(n14766), .B2(n1080), .ZN(n13885) );
  OAI22_X1 U3625 ( .A1(n6658), .A2(n1079), .B1(n14726), .B2(n1080), .ZN(n13886) );
  OAI22_X1 U3626 ( .A1(n6642), .A2(n1079), .B1(n14686), .B2(n1080), .ZN(n13887) );
  OAI22_X1 U3627 ( .A1(n6626), .A2(n1081), .B1(n14942), .B2(n1082), .ZN(n13888) );
  OAI22_X1 U3628 ( .A1(n6610), .A2(n1081), .B1(n14926), .B2(n1082), .ZN(n13889) );
  OAI22_X1 U3629 ( .A1(n6594), .A2(n1081), .B1(n14886), .B2(n1082), .ZN(n13890) );
  OAI22_X1 U3630 ( .A1(n6578), .A2(n1081), .B1(n14846), .B2(n1082), .ZN(n13891) );
  OAI22_X1 U3631 ( .A1(n6562), .A2(n1081), .B1(n14806), .B2(n1082), .ZN(n13892) );
  OAI22_X1 U3632 ( .A1(n6546), .A2(n1081), .B1(n14766), .B2(n1082), .ZN(n13893) );
  OAI22_X1 U3633 ( .A1(n6530), .A2(n1081), .B1(n14726), .B2(n1082), .ZN(n13894) );
  OAI22_X1 U3634 ( .A1(n6514), .A2(n1081), .B1(n14686), .B2(n1082), .ZN(n13895) );
  OAI22_X1 U3635 ( .A1(n6498), .A2(n1083), .B1(n14942), .B2(n1084), .ZN(n13896) );
  OAI22_X1 U3636 ( .A1(n6482), .A2(n1083), .B1(n14926), .B2(n1084), .ZN(n13897) );
  OAI22_X1 U3637 ( .A1(n6466), .A2(n1083), .B1(n14886), .B2(n1084), .ZN(n13898) );
  OAI22_X1 U3638 ( .A1(n6450), .A2(n1083), .B1(n14846), .B2(n1084), .ZN(n13899) );
  OAI22_X1 U3639 ( .A1(n6434), .A2(n1083), .B1(n14806), .B2(n1084), .ZN(n13900) );
  OAI22_X1 U3640 ( .A1(n6418), .A2(n1083), .B1(n14766), .B2(n1084), .ZN(n13901) );
  OAI22_X1 U3641 ( .A1(n6402), .A2(n1083), .B1(n14726), .B2(n1084), .ZN(n13902) );
  OAI22_X1 U3642 ( .A1(n6386), .A2(n1083), .B1(n14686), .B2(n1084), .ZN(n13903) );
  OAI22_X1 U3643 ( .A1(n6370), .A2(n1085), .B1(n14942), .B2(n1086), .ZN(n13904) );
  OAI22_X1 U3644 ( .A1(n6354), .A2(n1085), .B1(n14926), .B2(n1086), .ZN(n13905) );
  OAI22_X1 U3645 ( .A1(n6338), .A2(n1085), .B1(n14886), .B2(n1086), .ZN(n13906) );
  OAI22_X1 U3646 ( .A1(n6322), .A2(n1085), .B1(n14846), .B2(n1086), .ZN(n13907) );
  OAI22_X1 U3647 ( .A1(n6306), .A2(n1085), .B1(n14806), .B2(n1086), .ZN(n13908) );
  OAI22_X1 U3648 ( .A1(n6290), .A2(n1085), .B1(n14766), .B2(n1086), .ZN(n13909) );
  OAI22_X1 U3649 ( .A1(n6274), .A2(n1085), .B1(n14726), .B2(n1086), .ZN(n13910) );
  OAI22_X1 U3650 ( .A1(n6258), .A2(n1085), .B1(n14686), .B2(n1086), .ZN(n13911) );
  OAI22_X1 U3651 ( .A1(n6242), .A2(n1087), .B1(n14942), .B2(n1088), .ZN(n13912) );
  OAI22_X1 U3652 ( .A1(n6226), .A2(n1087), .B1(n14926), .B2(n1088), .ZN(n13913) );
  OAI22_X1 U3653 ( .A1(n6210), .A2(n1087), .B1(n14886), .B2(n1088), .ZN(n13914) );
  OAI22_X1 U3654 ( .A1(n6194), .A2(n1087), .B1(n14846), .B2(n1088), .ZN(n13915) );
  OAI22_X1 U3655 ( .A1(n6178), .A2(n1087), .B1(n14806), .B2(n1088), .ZN(n13916) );
  OAI22_X1 U3656 ( .A1(n6162), .A2(n1087), .B1(n14766), .B2(n1088), .ZN(n13917) );
  OAI22_X1 U3657 ( .A1(n6146), .A2(n1087), .B1(n14726), .B2(n1088), .ZN(n13918) );
  OAI22_X1 U3658 ( .A1(n6130), .A2(n1087), .B1(n14686), .B2(n1088), .ZN(n13919) );
  OAI22_X1 U3659 ( .A1(n6114), .A2(n1089), .B1(n14942), .B2(n1090), .ZN(n13920) );
  OAI22_X1 U3660 ( .A1(n6098), .A2(n1089), .B1(n14926), .B2(n1090), .ZN(n13921) );
  OAI22_X1 U3661 ( .A1(n6082), .A2(n1089), .B1(n14886), .B2(n1090), .ZN(n13922) );
  OAI22_X1 U3662 ( .A1(n6066), .A2(n1089), .B1(n14846), .B2(n1090), .ZN(n13923) );
  OAI22_X1 U3663 ( .A1(n6050), .A2(n1089), .B1(n14806), .B2(n1090), .ZN(n13924) );
  OAI22_X1 U3664 ( .A1(n6034), .A2(n1089), .B1(n14766), .B2(n1090), .ZN(n13925) );
  OAI22_X1 U3665 ( .A1(n6018), .A2(n1089), .B1(n14726), .B2(n1090), .ZN(n13926) );
  OAI22_X1 U3666 ( .A1(n6002), .A2(n1089), .B1(n14686), .B2(n1090), .ZN(n13927) );
  OAI22_X1 U3667 ( .A1(n7643), .A2(n409), .B1(n14967), .B2(n410), .ZN(n11264)
         );
  OAI22_X1 U3668 ( .A1(n7627), .A2(n409), .B1(n14901), .B2(n410), .ZN(n11265)
         );
  OAI22_X1 U3669 ( .A1(n7611), .A2(n409), .B1(n14861), .B2(n410), .ZN(n11266)
         );
  OAI22_X1 U3670 ( .A1(n7595), .A2(n409), .B1(n14821), .B2(n410), .ZN(n11267)
         );
  OAI22_X1 U3671 ( .A1(n7579), .A2(n409), .B1(n14781), .B2(n410), .ZN(n11268)
         );
  OAI22_X1 U3672 ( .A1(n7563), .A2(n409), .B1(n14741), .B2(n410), .ZN(n11269)
         );
  OAI22_X1 U3673 ( .A1(n7547), .A2(n409), .B1(n14701), .B2(n410), .ZN(n11270)
         );
  OAI22_X1 U3674 ( .A1(n7531), .A2(n409), .B1(n14661), .B2(n410), .ZN(n11271)
         );
  OAI22_X1 U3675 ( .A1(n7515), .A2(n411), .B1(n14967), .B2(n412), .ZN(n11272)
         );
  OAI22_X1 U3676 ( .A1(n7499), .A2(n411), .B1(n14901), .B2(n412), .ZN(n11273)
         );
  OAI22_X1 U3677 ( .A1(n7483), .A2(n411), .B1(n14861), .B2(n412), .ZN(n11274)
         );
  OAI22_X1 U3678 ( .A1(n7467), .A2(n411), .B1(n14821), .B2(n412), .ZN(n11275)
         );
  OAI22_X1 U3679 ( .A1(n7451), .A2(n411), .B1(n14781), .B2(n412), .ZN(n11276)
         );
  OAI22_X1 U3680 ( .A1(n7435), .A2(n411), .B1(n14741), .B2(n412), .ZN(n11277)
         );
  OAI22_X1 U3681 ( .A1(n7419), .A2(n411), .B1(n14701), .B2(n412), .ZN(n11278)
         );
  OAI22_X1 U3682 ( .A1(n7403), .A2(n411), .B1(n14661), .B2(n412), .ZN(n11279)
         );
  OAI22_X1 U3683 ( .A1(n7387), .A2(n413), .B1(n14967), .B2(n414), .ZN(n11280)
         );
  OAI22_X1 U3684 ( .A1(n7371), .A2(n413), .B1(n14901), .B2(n414), .ZN(n11281)
         );
  OAI22_X1 U3685 ( .A1(n7355), .A2(n413), .B1(n14861), .B2(n414), .ZN(n11282)
         );
  OAI22_X1 U3686 ( .A1(n7339), .A2(n413), .B1(n14821), .B2(n414), .ZN(n11283)
         );
  OAI22_X1 U3687 ( .A1(n7323), .A2(n413), .B1(n14781), .B2(n414), .ZN(n11284)
         );
  OAI22_X1 U3688 ( .A1(n7307), .A2(n413), .B1(n14741), .B2(n414), .ZN(n11285)
         );
  OAI22_X1 U3689 ( .A1(n7291), .A2(n413), .B1(n14701), .B2(n414), .ZN(n11286)
         );
  OAI22_X1 U3690 ( .A1(n7275), .A2(n413), .B1(n14661), .B2(n414), .ZN(n11287)
         );
  OAI22_X1 U3691 ( .A1(n7259), .A2(n415), .B1(n14967), .B2(n416), .ZN(n11288)
         );
  OAI22_X1 U3692 ( .A1(n7243), .A2(n415), .B1(n14901), .B2(n416), .ZN(n11289)
         );
  OAI22_X1 U3693 ( .A1(n7227), .A2(n415), .B1(n14861), .B2(n416), .ZN(n11290)
         );
  OAI22_X1 U3694 ( .A1(n7211), .A2(n415), .B1(n14821), .B2(n416), .ZN(n11291)
         );
  OAI22_X1 U3695 ( .A1(n7195), .A2(n415), .B1(n14781), .B2(n416), .ZN(n11292)
         );
  OAI22_X1 U3696 ( .A1(n7179), .A2(n415), .B1(n14741), .B2(n416), .ZN(n11293)
         );
  OAI22_X1 U3697 ( .A1(n7163), .A2(n415), .B1(n14701), .B2(n416), .ZN(n11294)
         );
  OAI22_X1 U3698 ( .A1(n7147), .A2(n415), .B1(n14661), .B2(n416), .ZN(n11295)
         );
  OAI22_X1 U3699 ( .A1(n7131), .A2(n417), .B1(n14967), .B2(n418), .ZN(n11296)
         );
  OAI22_X1 U3700 ( .A1(n7115), .A2(n417), .B1(n14901), .B2(n418), .ZN(n11297)
         );
  OAI22_X1 U3701 ( .A1(n7099), .A2(n417), .B1(n14861), .B2(n418), .ZN(n11298)
         );
  OAI22_X1 U3702 ( .A1(n7083), .A2(n417), .B1(n14821), .B2(n418), .ZN(n11299)
         );
  OAI22_X1 U3703 ( .A1(n7067), .A2(n417), .B1(n14781), .B2(n418), .ZN(n11300)
         );
  OAI22_X1 U3704 ( .A1(n7051), .A2(n417), .B1(n14741), .B2(n418), .ZN(n11301)
         );
  OAI22_X1 U3705 ( .A1(n7035), .A2(n417), .B1(n14701), .B2(n418), .ZN(n11302)
         );
  OAI22_X1 U3706 ( .A1(n7019), .A2(n417), .B1(n14661), .B2(n418), .ZN(n11303)
         );
  OAI22_X1 U3707 ( .A1(n7003), .A2(n419), .B1(n14967), .B2(n420), .ZN(n11304)
         );
  OAI22_X1 U3708 ( .A1(n6987), .A2(n419), .B1(n14901), .B2(n420), .ZN(n11305)
         );
  OAI22_X1 U3709 ( .A1(n6971), .A2(n419), .B1(n14861), .B2(n420), .ZN(n11306)
         );
  OAI22_X1 U3710 ( .A1(n6955), .A2(n419), .B1(n14821), .B2(n420), .ZN(n11307)
         );
  OAI22_X1 U3711 ( .A1(n6939), .A2(n419), .B1(n14781), .B2(n420), .ZN(n11308)
         );
  OAI22_X1 U3712 ( .A1(n6923), .A2(n419), .B1(n14741), .B2(n420), .ZN(n11309)
         );
  OAI22_X1 U3713 ( .A1(n6907), .A2(n419), .B1(n14701), .B2(n420), .ZN(n11310)
         );
  OAI22_X1 U3714 ( .A1(n6891), .A2(n419), .B1(n14661), .B2(n420), .ZN(n11311)
         );
  OAI22_X1 U3715 ( .A1(n6875), .A2(n421), .B1(n14967), .B2(n422), .ZN(n11312)
         );
  OAI22_X1 U3716 ( .A1(n6859), .A2(n421), .B1(n14901), .B2(n422), .ZN(n11313)
         );
  OAI22_X1 U3717 ( .A1(n6843), .A2(n421), .B1(n14861), .B2(n422), .ZN(n11314)
         );
  OAI22_X1 U3718 ( .A1(n6827), .A2(n421), .B1(n14821), .B2(n422), .ZN(n11315)
         );
  OAI22_X1 U3719 ( .A1(n6811), .A2(n421), .B1(n14781), .B2(n422), .ZN(n11316)
         );
  OAI22_X1 U3720 ( .A1(n6795), .A2(n421), .B1(n14741), .B2(n422), .ZN(n11317)
         );
  OAI22_X1 U3721 ( .A1(n6779), .A2(n421), .B1(n14701), .B2(n422), .ZN(n11318)
         );
  OAI22_X1 U3722 ( .A1(n6763), .A2(n421), .B1(n14661), .B2(n422), .ZN(n11319)
         );
  OAI22_X1 U3723 ( .A1(n6747), .A2(n423), .B1(n14967), .B2(n424), .ZN(n11320)
         );
  OAI22_X1 U3724 ( .A1(n6731), .A2(n423), .B1(n14901), .B2(n424), .ZN(n11321)
         );
  OAI22_X1 U3725 ( .A1(n6715), .A2(n423), .B1(n14861), .B2(n424), .ZN(n11322)
         );
  OAI22_X1 U3726 ( .A1(n6699), .A2(n423), .B1(n14821), .B2(n424), .ZN(n11323)
         );
  OAI22_X1 U3727 ( .A1(n6683), .A2(n423), .B1(n14781), .B2(n424), .ZN(n11324)
         );
  OAI22_X1 U3728 ( .A1(n6667), .A2(n423), .B1(n14741), .B2(n424), .ZN(n11325)
         );
  OAI22_X1 U3729 ( .A1(n6651), .A2(n423), .B1(n14701), .B2(n424), .ZN(n11326)
         );
  OAI22_X1 U3730 ( .A1(n6635), .A2(n423), .B1(n14661), .B2(n424), .ZN(n11327)
         );
  OAI22_X1 U3731 ( .A1(n6619), .A2(n425), .B1(n14967), .B2(n426), .ZN(n11328)
         );
  OAI22_X1 U3732 ( .A1(n6603), .A2(n425), .B1(n14901), .B2(n426), .ZN(n11329)
         );
  OAI22_X1 U3733 ( .A1(n6587), .A2(n425), .B1(n14861), .B2(n426), .ZN(n11330)
         );
  OAI22_X1 U3734 ( .A1(n6571), .A2(n425), .B1(n14821), .B2(n426), .ZN(n11331)
         );
  OAI22_X1 U3735 ( .A1(n6555), .A2(n425), .B1(n14781), .B2(n426), .ZN(n11332)
         );
  OAI22_X1 U3736 ( .A1(n6539), .A2(n425), .B1(n14741), .B2(n426), .ZN(n11333)
         );
  OAI22_X1 U3737 ( .A1(n6523), .A2(n425), .B1(n14701), .B2(n426), .ZN(n11334)
         );
  OAI22_X1 U3738 ( .A1(n6507), .A2(n425), .B1(n14661), .B2(n426), .ZN(n11335)
         );
  OAI22_X1 U3739 ( .A1(n6491), .A2(n427), .B1(n14967), .B2(n428), .ZN(n11336)
         );
  OAI22_X1 U3740 ( .A1(n6475), .A2(n427), .B1(n14902), .B2(n428), .ZN(n11337)
         );
  OAI22_X1 U3741 ( .A1(n6459), .A2(n427), .B1(n14862), .B2(n428), .ZN(n11338)
         );
  OAI22_X1 U3742 ( .A1(n6443), .A2(n427), .B1(n14822), .B2(n428), .ZN(n11339)
         );
  OAI22_X1 U3743 ( .A1(n6427), .A2(n427), .B1(n14782), .B2(n428), .ZN(n11340)
         );
  OAI22_X1 U3744 ( .A1(n6411), .A2(n427), .B1(n14742), .B2(n428), .ZN(n11341)
         );
  OAI22_X1 U3745 ( .A1(n6395), .A2(n427), .B1(n14702), .B2(n428), .ZN(n11342)
         );
  OAI22_X1 U3746 ( .A1(n6379), .A2(n427), .B1(n14662), .B2(n428), .ZN(n11343)
         );
  OAI22_X1 U3747 ( .A1(n6363), .A2(n429), .B1(n14967), .B2(n430), .ZN(n11344)
         );
  OAI22_X1 U3748 ( .A1(n6347), .A2(n429), .B1(n14902), .B2(n430), .ZN(n11345)
         );
  OAI22_X1 U3749 ( .A1(n6331), .A2(n429), .B1(n14862), .B2(n430), .ZN(n11346)
         );
  OAI22_X1 U3750 ( .A1(n6315), .A2(n429), .B1(n14822), .B2(n430), .ZN(n11347)
         );
  OAI22_X1 U3751 ( .A1(n6299), .A2(n429), .B1(n14782), .B2(n430), .ZN(n11348)
         );
  OAI22_X1 U3752 ( .A1(n6283), .A2(n429), .B1(n14742), .B2(n430), .ZN(n11349)
         );
  OAI22_X1 U3753 ( .A1(n6267), .A2(n429), .B1(n14702), .B2(n430), .ZN(n11350)
         );
  OAI22_X1 U3754 ( .A1(n6251), .A2(n429), .B1(n14662), .B2(n430), .ZN(n11351)
         );
  OAI22_X1 U3755 ( .A1(n6235), .A2(n431), .B1(n14967), .B2(n432), .ZN(n11352)
         );
  OAI22_X1 U3756 ( .A1(n6219), .A2(n431), .B1(n14902), .B2(n432), .ZN(n11353)
         );
  OAI22_X1 U3757 ( .A1(n6203), .A2(n431), .B1(n14862), .B2(n432), .ZN(n11354)
         );
  OAI22_X1 U3758 ( .A1(n6187), .A2(n431), .B1(n14822), .B2(n432), .ZN(n11355)
         );
  OAI22_X1 U3759 ( .A1(n6171), .A2(n431), .B1(n14782), .B2(n432), .ZN(n11356)
         );
  OAI22_X1 U3760 ( .A1(n6155), .A2(n431), .B1(n14742), .B2(n432), .ZN(n11357)
         );
  OAI22_X1 U3761 ( .A1(n6139), .A2(n431), .B1(n14702), .B2(n432), .ZN(n11358)
         );
  OAI22_X1 U3762 ( .A1(n6123), .A2(n431), .B1(n14662), .B2(n432), .ZN(n11359)
         );
  OAI22_X1 U3763 ( .A1(n6107), .A2(n433), .B1(n14966), .B2(n434), .ZN(n11360)
         );
  OAI22_X1 U3764 ( .A1(n6091), .A2(n433), .B1(n14902), .B2(n434), .ZN(n11361)
         );
  OAI22_X1 U3765 ( .A1(n6075), .A2(n433), .B1(n14862), .B2(n434), .ZN(n11362)
         );
  OAI22_X1 U3766 ( .A1(n6059), .A2(n433), .B1(n14822), .B2(n434), .ZN(n11363)
         );
  OAI22_X1 U3767 ( .A1(n6043), .A2(n433), .B1(n14782), .B2(n434), .ZN(n11364)
         );
  OAI22_X1 U3768 ( .A1(n6027), .A2(n433), .B1(n14742), .B2(n434), .ZN(n11365)
         );
  OAI22_X1 U3769 ( .A1(n6011), .A2(n433), .B1(n14702), .B2(n434), .ZN(n11366)
         );
  OAI22_X1 U3770 ( .A1(n5995), .A2(n433), .B1(n14662), .B2(n434), .ZN(n11367)
         );
  OAI22_X1 U3771 ( .A1(n7647), .A2(n475), .B1(n14965), .B2(n476), .ZN(n11520)
         );
  OAI22_X1 U3772 ( .A1(n7631), .A2(n475), .B1(n14903), .B2(n476), .ZN(n11521)
         );
  OAI22_X1 U3773 ( .A1(n7615), .A2(n475), .B1(n14863), .B2(n476), .ZN(n11522)
         );
  OAI22_X1 U3774 ( .A1(n7599), .A2(n475), .B1(n14823), .B2(n476), .ZN(n11523)
         );
  OAI22_X1 U3775 ( .A1(n7583), .A2(n475), .B1(n14783), .B2(n476), .ZN(n11524)
         );
  OAI22_X1 U3776 ( .A1(n7567), .A2(n475), .B1(n14743), .B2(n476), .ZN(n11525)
         );
  OAI22_X1 U3777 ( .A1(n7551), .A2(n475), .B1(n14703), .B2(n476), .ZN(n11526)
         );
  OAI22_X1 U3778 ( .A1(n7535), .A2(n475), .B1(n14663), .B2(n476), .ZN(n11527)
         );
  OAI22_X1 U3779 ( .A1(n7519), .A2(n477), .B1(n14965), .B2(n478), .ZN(n11528)
         );
  OAI22_X1 U3780 ( .A1(n7503), .A2(n477), .B1(n14903), .B2(n478), .ZN(n11529)
         );
  OAI22_X1 U3781 ( .A1(n7487), .A2(n477), .B1(n14863), .B2(n478), .ZN(n11530)
         );
  OAI22_X1 U3782 ( .A1(n7471), .A2(n477), .B1(n14823), .B2(n478), .ZN(n11531)
         );
  OAI22_X1 U3783 ( .A1(n7455), .A2(n477), .B1(n14783), .B2(n478), .ZN(n11532)
         );
  OAI22_X1 U3784 ( .A1(n7439), .A2(n477), .B1(n14743), .B2(n478), .ZN(n11533)
         );
  OAI22_X1 U3785 ( .A1(n7423), .A2(n477), .B1(n14703), .B2(n478), .ZN(n11534)
         );
  OAI22_X1 U3786 ( .A1(n7407), .A2(n477), .B1(n14663), .B2(n478), .ZN(n11535)
         );
  OAI22_X1 U3787 ( .A1(n7391), .A2(n479), .B1(n14965), .B2(n480), .ZN(n11536)
         );
  OAI22_X1 U3788 ( .A1(n7375), .A2(n479), .B1(n14903), .B2(n480), .ZN(n11537)
         );
  OAI22_X1 U3789 ( .A1(n7359), .A2(n479), .B1(n14863), .B2(n480), .ZN(n11538)
         );
  OAI22_X1 U3790 ( .A1(n7343), .A2(n479), .B1(n14823), .B2(n480), .ZN(n11539)
         );
  OAI22_X1 U3791 ( .A1(n7327), .A2(n479), .B1(n14783), .B2(n480), .ZN(n11540)
         );
  OAI22_X1 U3792 ( .A1(n7311), .A2(n479), .B1(n14743), .B2(n480), .ZN(n11541)
         );
  OAI22_X1 U3793 ( .A1(n7295), .A2(n479), .B1(n14703), .B2(n480), .ZN(n11542)
         );
  OAI22_X1 U3794 ( .A1(n7279), .A2(n479), .B1(n14663), .B2(n480), .ZN(n11543)
         );
  OAI22_X1 U3795 ( .A1(n7263), .A2(n481), .B1(n14965), .B2(n482), .ZN(n11544)
         );
  OAI22_X1 U3796 ( .A1(n7247), .A2(n481), .B1(n14904), .B2(n482), .ZN(n11545)
         );
  OAI22_X1 U3797 ( .A1(n7231), .A2(n481), .B1(n14864), .B2(n482), .ZN(n11546)
         );
  OAI22_X1 U3798 ( .A1(n7215), .A2(n481), .B1(n14824), .B2(n482), .ZN(n11547)
         );
  OAI22_X1 U3799 ( .A1(n7199), .A2(n481), .B1(n14784), .B2(n482), .ZN(n11548)
         );
  OAI22_X1 U3800 ( .A1(n7183), .A2(n481), .B1(n14744), .B2(n482), .ZN(n11549)
         );
  OAI22_X1 U3801 ( .A1(n7167), .A2(n481), .B1(n14704), .B2(n482), .ZN(n11550)
         );
  OAI22_X1 U3802 ( .A1(n7151), .A2(n481), .B1(n14664), .B2(n482), .ZN(n11551)
         );
  OAI22_X1 U3803 ( .A1(n7135), .A2(n483), .B1(n14965), .B2(n484), .ZN(n11552)
         );
  OAI22_X1 U3804 ( .A1(n7119), .A2(n483), .B1(n14904), .B2(n484), .ZN(n11553)
         );
  OAI22_X1 U3805 ( .A1(n7103), .A2(n483), .B1(n14864), .B2(n484), .ZN(n11554)
         );
  OAI22_X1 U3806 ( .A1(n7087), .A2(n483), .B1(n14824), .B2(n484), .ZN(n11555)
         );
  OAI22_X1 U3807 ( .A1(n7071), .A2(n483), .B1(n14784), .B2(n484), .ZN(n11556)
         );
  OAI22_X1 U3808 ( .A1(n7055), .A2(n483), .B1(n14744), .B2(n484), .ZN(n11557)
         );
  OAI22_X1 U3809 ( .A1(n7039), .A2(n483), .B1(n14704), .B2(n484), .ZN(n11558)
         );
  OAI22_X1 U3810 ( .A1(n7023), .A2(n483), .B1(n14664), .B2(n484), .ZN(n11559)
         );
  OAI22_X1 U3811 ( .A1(n7007), .A2(n485), .B1(n14965), .B2(n486), .ZN(n11560)
         );
  OAI22_X1 U3812 ( .A1(n6991), .A2(n485), .B1(n14904), .B2(n486), .ZN(n11561)
         );
  OAI22_X1 U3813 ( .A1(n6975), .A2(n485), .B1(n14864), .B2(n486), .ZN(n11562)
         );
  OAI22_X1 U3814 ( .A1(n6959), .A2(n485), .B1(n14824), .B2(n486), .ZN(n11563)
         );
  OAI22_X1 U3815 ( .A1(n6943), .A2(n485), .B1(n14784), .B2(n486), .ZN(n11564)
         );
  OAI22_X1 U3816 ( .A1(n6927), .A2(n485), .B1(n14744), .B2(n486), .ZN(n11565)
         );
  OAI22_X1 U3817 ( .A1(n6911), .A2(n485), .B1(n14704), .B2(n486), .ZN(n11566)
         );
  OAI22_X1 U3818 ( .A1(n6895), .A2(n485), .B1(n14664), .B2(n486), .ZN(n11567)
         );
  OAI22_X1 U3819 ( .A1(n6879), .A2(n487), .B1(n14964), .B2(n488), .ZN(n11568)
         );
  OAI22_X1 U3820 ( .A1(n6863), .A2(n487), .B1(n14904), .B2(n488), .ZN(n11569)
         );
  OAI22_X1 U3821 ( .A1(n6847), .A2(n487), .B1(n14864), .B2(n488), .ZN(n11570)
         );
  OAI22_X1 U3822 ( .A1(n6831), .A2(n487), .B1(n14824), .B2(n488), .ZN(n11571)
         );
  OAI22_X1 U3823 ( .A1(n6815), .A2(n487), .B1(n14784), .B2(n488), .ZN(n11572)
         );
  OAI22_X1 U3824 ( .A1(n6799), .A2(n487), .B1(n14744), .B2(n488), .ZN(n11573)
         );
  OAI22_X1 U3825 ( .A1(n6783), .A2(n487), .B1(n14704), .B2(n488), .ZN(n11574)
         );
  OAI22_X1 U3826 ( .A1(n6767), .A2(n487), .B1(n14664), .B2(n488), .ZN(n11575)
         );
  OAI22_X1 U3827 ( .A1(n6751), .A2(n489), .B1(n14964), .B2(n490), .ZN(n11576)
         );
  OAI22_X1 U3828 ( .A1(n6735), .A2(n489), .B1(n14904), .B2(n490), .ZN(n11577)
         );
  OAI22_X1 U3829 ( .A1(n6719), .A2(n489), .B1(n14864), .B2(n490), .ZN(n11578)
         );
  OAI22_X1 U3830 ( .A1(n6703), .A2(n489), .B1(n14824), .B2(n490), .ZN(n11579)
         );
  OAI22_X1 U3831 ( .A1(n6687), .A2(n489), .B1(n14784), .B2(n490), .ZN(n11580)
         );
  OAI22_X1 U3832 ( .A1(n6671), .A2(n489), .B1(n14744), .B2(n490), .ZN(n11581)
         );
  OAI22_X1 U3833 ( .A1(n6655), .A2(n489), .B1(n14704), .B2(n490), .ZN(n11582)
         );
  OAI22_X1 U3834 ( .A1(n6639), .A2(n489), .B1(n14664), .B2(n490), .ZN(n11583)
         );
  OAI22_X1 U3835 ( .A1(n6623), .A2(n491), .B1(n14964), .B2(n492), .ZN(n11584)
         );
  OAI22_X1 U3836 ( .A1(n6607), .A2(n491), .B1(n14904), .B2(n492), .ZN(n11585)
         );
  OAI22_X1 U3837 ( .A1(n6591), .A2(n491), .B1(n14864), .B2(n492), .ZN(n11586)
         );
  OAI22_X1 U3838 ( .A1(n6575), .A2(n491), .B1(n14824), .B2(n492), .ZN(n11587)
         );
  OAI22_X1 U3839 ( .A1(n6559), .A2(n491), .B1(n14784), .B2(n492), .ZN(n11588)
         );
  OAI22_X1 U3840 ( .A1(n6543), .A2(n491), .B1(n14744), .B2(n492), .ZN(n11589)
         );
  OAI22_X1 U3841 ( .A1(n6527), .A2(n491), .B1(n14704), .B2(n492), .ZN(n11590)
         );
  OAI22_X1 U3842 ( .A1(n6511), .A2(n491), .B1(n14664), .B2(n492), .ZN(n11591)
         );
  OAI22_X1 U3843 ( .A1(n6495), .A2(n493), .B1(n14964), .B2(n494), .ZN(n11592)
         );
  OAI22_X1 U3844 ( .A1(n6479), .A2(n493), .B1(n14904), .B2(n494), .ZN(n11593)
         );
  OAI22_X1 U3845 ( .A1(n6463), .A2(n493), .B1(n14864), .B2(n494), .ZN(n11594)
         );
  OAI22_X1 U3846 ( .A1(n6447), .A2(n493), .B1(n14824), .B2(n494), .ZN(n11595)
         );
  OAI22_X1 U3847 ( .A1(n6431), .A2(n493), .B1(n14784), .B2(n494), .ZN(n11596)
         );
  OAI22_X1 U3848 ( .A1(n6415), .A2(n493), .B1(n14744), .B2(n494), .ZN(n11597)
         );
  OAI22_X1 U3849 ( .A1(n6399), .A2(n493), .B1(n14704), .B2(n494), .ZN(n11598)
         );
  OAI22_X1 U3850 ( .A1(n6383), .A2(n493), .B1(n14664), .B2(n494), .ZN(n11599)
         );
  OAI22_X1 U3851 ( .A1(n6367), .A2(n495), .B1(n14964), .B2(n496), .ZN(n11600)
         );
  OAI22_X1 U3852 ( .A1(n6351), .A2(n495), .B1(n14904), .B2(n496), .ZN(n11601)
         );
  OAI22_X1 U3853 ( .A1(n6335), .A2(n495), .B1(n14864), .B2(n496), .ZN(n11602)
         );
  OAI22_X1 U3854 ( .A1(n6319), .A2(n495), .B1(n14824), .B2(n496), .ZN(n11603)
         );
  OAI22_X1 U3855 ( .A1(n6303), .A2(n495), .B1(n14784), .B2(n496), .ZN(n11604)
         );
  OAI22_X1 U3856 ( .A1(n6287), .A2(n495), .B1(n14744), .B2(n496), .ZN(n11605)
         );
  OAI22_X1 U3857 ( .A1(n6271), .A2(n495), .B1(n14704), .B2(n496), .ZN(n11606)
         );
  OAI22_X1 U3858 ( .A1(n6255), .A2(n495), .B1(n14664), .B2(n496), .ZN(n11607)
         );
  OAI22_X1 U3859 ( .A1(n6239), .A2(n497), .B1(n14964), .B2(n498), .ZN(n11608)
         );
  OAI22_X1 U3860 ( .A1(n6223), .A2(n497), .B1(n14904), .B2(n498), .ZN(n11609)
         );
  OAI22_X1 U3861 ( .A1(n6207), .A2(n497), .B1(n14864), .B2(n498), .ZN(n11610)
         );
  OAI22_X1 U3862 ( .A1(n6191), .A2(n497), .B1(n14824), .B2(n498), .ZN(n11611)
         );
  OAI22_X1 U3863 ( .A1(n6175), .A2(n497), .B1(n14784), .B2(n498), .ZN(n11612)
         );
  OAI22_X1 U3864 ( .A1(n6159), .A2(n497), .B1(n14744), .B2(n498), .ZN(n11613)
         );
  OAI22_X1 U3865 ( .A1(n6143), .A2(n497), .B1(n14704), .B2(n498), .ZN(n11614)
         );
  OAI22_X1 U3866 ( .A1(n6127), .A2(n497), .B1(n14664), .B2(n498), .ZN(n11615)
         );
  OAI22_X1 U3867 ( .A1(n6111), .A2(n499), .B1(n14964), .B2(n500), .ZN(n11616)
         );
  OAI22_X1 U3868 ( .A1(n6095), .A2(n499), .B1(n14904), .B2(n500), .ZN(n11617)
         );
  OAI22_X1 U3869 ( .A1(n6079), .A2(n499), .B1(n14864), .B2(n500), .ZN(n11618)
         );
  OAI22_X1 U3870 ( .A1(n6063), .A2(n499), .B1(n14824), .B2(n500), .ZN(n11619)
         );
  OAI22_X1 U3871 ( .A1(n6047), .A2(n499), .B1(n14784), .B2(n500), .ZN(n11620)
         );
  OAI22_X1 U3872 ( .A1(n6031), .A2(n499), .B1(n14744), .B2(n500), .ZN(n11621)
         );
  OAI22_X1 U3873 ( .A1(n6015), .A2(n499), .B1(n14704), .B2(n500), .ZN(n11622)
         );
  OAI22_X1 U3874 ( .A1(n5999), .A2(n499), .B1(n14664), .B2(n500), .ZN(n11623)
         );
  OAI22_X1 U3875 ( .A1(n7642), .A2(n933), .B1(n14948), .B2(n934), .ZN(n13312)
         );
  OAI22_X1 U3876 ( .A1(n7626), .A2(n933), .B1(n14921), .B2(n934), .ZN(n13313)
         );
  OAI22_X1 U3877 ( .A1(n7610), .A2(n933), .B1(n14881), .B2(n934), .ZN(n13314)
         );
  OAI22_X1 U3878 ( .A1(n7594), .A2(n933), .B1(n14841), .B2(n934), .ZN(n13315)
         );
  OAI22_X1 U3879 ( .A1(n7578), .A2(n933), .B1(n14801), .B2(n934), .ZN(n13316)
         );
  OAI22_X1 U3880 ( .A1(n7562), .A2(n933), .B1(n14761), .B2(n934), .ZN(n13317)
         );
  OAI22_X1 U3881 ( .A1(n7546), .A2(n933), .B1(n14721), .B2(n934), .ZN(n13318)
         );
  OAI22_X1 U3882 ( .A1(n7530), .A2(n933), .B1(n14681), .B2(n934), .ZN(n13319)
         );
  OAI22_X1 U3883 ( .A1(n7514), .A2(n935), .B1(n14948), .B2(n936), .ZN(n13320)
         );
  OAI22_X1 U3884 ( .A1(n7498), .A2(n935), .B1(n14921), .B2(n936), .ZN(n13321)
         );
  OAI22_X1 U3885 ( .A1(n7482), .A2(n935), .B1(n14881), .B2(n936), .ZN(n13322)
         );
  OAI22_X1 U3886 ( .A1(n7466), .A2(n935), .B1(n14841), .B2(n936), .ZN(n13323)
         );
  OAI22_X1 U3887 ( .A1(n7450), .A2(n935), .B1(n14801), .B2(n936), .ZN(n13324)
         );
  OAI22_X1 U3888 ( .A1(n7434), .A2(n935), .B1(n14761), .B2(n936), .ZN(n13325)
         );
  OAI22_X1 U3889 ( .A1(n7418), .A2(n935), .B1(n14721), .B2(n936), .ZN(n13326)
         );
  OAI22_X1 U3890 ( .A1(n7402), .A2(n935), .B1(n14681), .B2(n936), .ZN(n13327)
         );
  OAI22_X1 U3891 ( .A1(n7386), .A2(n937), .B1(n14948), .B2(n938), .ZN(n13328)
         );
  OAI22_X1 U3892 ( .A1(n7370), .A2(n937), .B1(n14921), .B2(n938), .ZN(n13329)
         );
  OAI22_X1 U3893 ( .A1(n7354), .A2(n937), .B1(n14881), .B2(n938), .ZN(n13330)
         );
  OAI22_X1 U3894 ( .A1(n7338), .A2(n937), .B1(n14841), .B2(n938), .ZN(n13331)
         );
  OAI22_X1 U3895 ( .A1(n7322), .A2(n937), .B1(n14801), .B2(n938), .ZN(n13332)
         );
  OAI22_X1 U3896 ( .A1(n7306), .A2(n937), .B1(n14761), .B2(n938), .ZN(n13333)
         );
  OAI22_X1 U3897 ( .A1(n7290), .A2(n937), .B1(n14721), .B2(n938), .ZN(n13334)
         );
  OAI22_X1 U3898 ( .A1(n7274), .A2(n937), .B1(n14681), .B2(n938), .ZN(n13335)
         );
  OAI22_X1 U3899 ( .A1(n7258), .A2(n939), .B1(n14947), .B2(n940), .ZN(n13336)
         );
  OAI22_X1 U3900 ( .A1(n7242), .A2(n939), .B1(n14921), .B2(n940), .ZN(n13337)
         );
  OAI22_X1 U3901 ( .A1(n7226), .A2(n939), .B1(n14881), .B2(n940), .ZN(n13338)
         );
  OAI22_X1 U3902 ( .A1(n7210), .A2(n939), .B1(n14841), .B2(n940), .ZN(n13339)
         );
  OAI22_X1 U3903 ( .A1(n7194), .A2(n939), .B1(n14801), .B2(n940), .ZN(n13340)
         );
  OAI22_X1 U3904 ( .A1(n7178), .A2(n939), .B1(n14761), .B2(n940), .ZN(n13341)
         );
  OAI22_X1 U3905 ( .A1(n7162), .A2(n939), .B1(n14721), .B2(n940), .ZN(n13342)
         );
  OAI22_X1 U3906 ( .A1(n7146), .A2(n939), .B1(n14681), .B2(n940), .ZN(n13343)
         );
  OAI22_X1 U3907 ( .A1(n7130), .A2(n941), .B1(n14947), .B2(n942), .ZN(n13344)
         );
  OAI22_X1 U3908 ( .A1(n7114), .A2(n941), .B1(n14921), .B2(n942), .ZN(n13345)
         );
  OAI22_X1 U3909 ( .A1(n7098), .A2(n941), .B1(n14881), .B2(n942), .ZN(n13346)
         );
  OAI22_X1 U3910 ( .A1(n7082), .A2(n941), .B1(n14841), .B2(n942), .ZN(n13347)
         );
  OAI22_X1 U3911 ( .A1(n7066), .A2(n941), .B1(n14801), .B2(n942), .ZN(n13348)
         );
  OAI22_X1 U3912 ( .A1(n7050), .A2(n941), .B1(n14761), .B2(n942), .ZN(n13349)
         );
  OAI22_X1 U3913 ( .A1(n7034), .A2(n941), .B1(n14721), .B2(n942), .ZN(n13350)
         );
  OAI22_X1 U3914 ( .A1(n7018), .A2(n941), .B1(n14681), .B2(n942), .ZN(n13351)
         );
  OAI22_X1 U3915 ( .A1(n7002), .A2(n943), .B1(n14947), .B2(n944), .ZN(n13352)
         );
  OAI22_X1 U3916 ( .A1(n6986), .A2(n943), .B1(n14921), .B2(n944), .ZN(n13353)
         );
  OAI22_X1 U3917 ( .A1(n6970), .A2(n943), .B1(n14881), .B2(n944), .ZN(n13354)
         );
  OAI22_X1 U3918 ( .A1(n6954), .A2(n943), .B1(n14841), .B2(n944), .ZN(n13355)
         );
  OAI22_X1 U3919 ( .A1(n6938), .A2(n943), .B1(n14801), .B2(n944), .ZN(n13356)
         );
  OAI22_X1 U3920 ( .A1(n6922), .A2(n943), .B1(n14761), .B2(n944), .ZN(n13357)
         );
  OAI22_X1 U3921 ( .A1(n6906), .A2(n943), .B1(n14721), .B2(n944), .ZN(n13358)
         );
  OAI22_X1 U3922 ( .A1(n6890), .A2(n943), .B1(n14681), .B2(n944), .ZN(n13359)
         );
  OAI22_X1 U3923 ( .A1(n6874), .A2(n945), .B1(n14947), .B2(n946), .ZN(n13360)
         );
  OAI22_X1 U3924 ( .A1(n6858), .A2(n945), .B1(n14921), .B2(n946), .ZN(n13361)
         );
  OAI22_X1 U3925 ( .A1(n6842), .A2(n945), .B1(n14881), .B2(n946), .ZN(n13362)
         );
  OAI22_X1 U3926 ( .A1(n6826), .A2(n945), .B1(n14841), .B2(n946), .ZN(n13363)
         );
  OAI22_X1 U3927 ( .A1(n6810), .A2(n945), .B1(n14801), .B2(n946), .ZN(n13364)
         );
  OAI22_X1 U3928 ( .A1(n6794), .A2(n945), .B1(n14761), .B2(n946), .ZN(n13365)
         );
  OAI22_X1 U3929 ( .A1(n6778), .A2(n945), .B1(n14721), .B2(n946), .ZN(n13366)
         );
  OAI22_X1 U3930 ( .A1(n6762), .A2(n945), .B1(n14681), .B2(n946), .ZN(n13367)
         );
  OAI22_X1 U3931 ( .A1(n6746), .A2(n947), .B1(n14947), .B2(n948), .ZN(n13368)
         );
  OAI22_X1 U3932 ( .A1(n6730), .A2(n947), .B1(n14921), .B2(n948), .ZN(n13369)
         );
  OAI22_X1 U3933 ( .A1(n6714), .A2(n947), .B1(n14881), .B2(n948), .ZN(n13370)
         );
  OAI22_X1 U3934 ( .A1(n6698), .A2(n947), .B1(n14841), .B2(n948), .ZN(n13371)
         );
  OAI22_X1 U3935 ( .A1(n6682), .A2(n947), .B1(n14801), .B2(n948), .ZN(n13372)
         );
  OAI22_X1 U3936 ( .A1(n6666), .A2(n947), .B1(n14761), .B2(n948), .ZN(n13373)
         );
  OAI22_X1 U3937 ( .A1(n6650), .A2(n947), .B1(n14721), .B2(n948), .ZN(n13374)
         );
  OAI22_X1 U3938 ( .A1(n6634), .A2(n947), .B1(n14681), .B2(n948), .ZN(n13375)
         );
  OAI22_X1 U3939 ( .A1(n6618), .A2(n949), .B1(n14947), .B2(n950), .ZN(n13376)
         );
  OAI22_X1 U3940 ( .A1(n6602), .A2(n949), .B1(n14921), .B2(n950), .ZN(n13377)
         );
  OAI22_X1 U3941 ( .A1(n6586), .A2(n949), .B1(n14881), .B2(n950), .ZN(n13378)
         );
  OAI22_X1 U3942 ( .A1(n6570), .A2(n949), .B1(n14841), .B2(n950), .ZN(n13379)
         );
  OAI22_X1 U3943 ( .A1(n6554), .A2(n949), .B1(n14801), .B2(n950), .ZN(n13380)
         );
  OAI22_X1 U3944 ( .A1(n6538), .A2(n949), .B1(n14761), .B2(n950), .ZN(n13381)
         );
  OAI22_X1 U3945 ( .A1(n6522), .A2(n949), .B1(n14721), .B2(n950), .ZN(n13382)
         );
  OAI22_X1 U3946 ( .A1(n6506), .A2(n949), .B1(n14681), .B2(n950), .ZN(n13383)
         );
  OAI22_X1 U3947 ( .A1(n6490), .A2(n951), .B1(n14947), .B2(n952), .ZN(n13384)
         );
  OAI22_X1 U3948 ( .A1(n6474), .A2(n951), .B1(n14921), .B2(n952), .ZN(n13385)
         );
  OAI22_X1 U3949 ( .A1(n6458), .A2(n951), .B1(n14881), .B2(n952), .ZN(n13386)
         );
  OAI22_X1 U3950 ( .A1(n6442), .A2(n951), .B1(n14841), .B2(n952), .ZN(n13387)
         );
  OAI22_X1 U3951 ( .A1(n6426), .A2(n951), .B1(n14801), .B2(n952), .ZN(n13388)
         );
  OAI22_X1 U3952 ( .A1(n6410), .A2(n951), .B1(n14761), .B2(n952), .ZN(n13389)
         );
  OAI22_X1 U3953 ( .A1(n6394), .A2(n951), .B1(n14721), .B2(n952), .ZN(n13390)
         );
  OAI22_X1 U3954 ( .A1(n6378), .A2(n951), .B1(n14681), .B2(n952), .ZN(n13391)
         );
  OAI22_X1 U3955 ( .A1(n6362), .A2(n953), .B1(n14947), .B2(n954), .ZN(n13392)
         );
  OAI22_X1 U3956 ( .A1(n6346), .A2(n953), .B1(n14921), .B2(n954), .ZN(n13393)
         );
  OAI22_X1 U3957 ( .A1(n6330), .A2(n953), .B1(n14881), .B2(n954), .ZN(n13394)
         );
  OAI22_X1 U3958 ( .A1(n6314), .A2(n953), .B1(n14841), .B2(n954), .ZN(n13395)
         );
  OAI22_X1 U3959 ( .A1(n6298), .A2(n953), .B1(n14801), .B2(n954), .ZN(n13396)
         );
  OAI22_X1 U3960 ( .A1(n6282), .A2(n953), .B1(n14761), .B2(n954), .ZN(n13397)
         );
  OAI22_X1 U3961 ( .A1(n6266), .A2(n953), .B1(n14721), .B2(n954), .ZN(n13398)
         );
  OAI22_X1 U3962 ( .A1(n6250), .A2(n953), .B1(n14681), .B2(n954), .ZN(n13399)
         );
  OAI22_X1 U3963 ( .A1(n6234), .A2(n955), .B1(n14947), .B2(n956), .ZN(n13400)
         );
  OAI22_X1 U3964 ( .A1(n6218), .A2(n955), .B1(n14921), .B2(n956), .ZN(n13401)
         );
  OAI22_X1 U3965 ( .A1(n6202), .A2(n955), .B1(n14881), .B2(n956), .ZN(n13402)
         );
  OAI22_X1 U3966 ( .A1(n6186), .A2(n955), .B1(n14841), .B2(n956), .ZN(n13403)
         );
  OAI22_X1 U3967 ( .A1(n6170), .A2(n955), .B1(n14801), .B2(n956), .ZN(n13404)
         );
  OAI22_X1 U3968 ( .A1(n6154), .A2(n955), .B1(n14761), .B2(n956), .ZN(n13405)
         );
  OAI22_X1 U3969 ( .A1(n6138), .A2(n955), .B1(n14721), .B2(n956), .ZN(n13406)
         );
  OAI22_X1 U3970 ( .A1(n6122), .A2(n955), .B1(n14681), .B2(n956), .ZN(n13407)
         );
  OAI22_X1 U3971 ( .A1(n6106), .A2(n957), .B1(n14947), .B2(n958), .ZN(n13408)
         );
  OAI22_X1 U3972 ( .A1(n6090), .A2(n957), .B1(n14921), .B2(n958), .ZN(n13409)
         );
  OAI22_X1 U3973 ( .A1(n6074), .A2(n957), .B1(n14881), .B2(n958), .ZN(n13410)
         );
  OAI22_X1 U3974 ( .A1(n6058), .A2(n957), .B1(n14841), .B2(n958), .ZN(n13411)
         );
  OAI22_X1 U3975 ( .A1(n6042), .A2(n957), .B1(n14801), .B2(n958), .ZN(n13412)
         );
  OAI22_X1 U3976 ( .A1(n6026), .A2(n957), .B1(n14761), .B2(n958), .ZN(n13413)
         );
  OAI22_X1 U3977 ( .A1(n6010), .A2(n957), .B1(n14721), .B2(n958), .ZN(n13414)
         );
  OAI22_X1 U3978 ( .A1(n5994), .A2(n957), .B1(n14681), .B2(n958), .ZN(n13415)
         );
  OAI22_X1 U3979 ( .A1(n9945), .A2(n78), .B1(n14930), .B2(n79), .ZN(n10096) );
  OAI22_X1 U3980 ( .A1(n9929), .A2(n78), .B1(n14890), .B2(n79), .ZN(n10097) );
  OAI22_X1 U3981 ( .A1(n9913), .A2(n78), .B1(n14850), .B2(n79), .ZN(n10098) );
  OAI22_X1 U3982 ( .A1(n9897), .A2(n78), .B1(n14810), .B2(n79), .ZN(n10099) );
  OAI22_X1 U3983 ( .A1(n9881), .A2(n78), .B1(n14770), .B2(n79), .ZN(n10100) );
  OAI22_X1 U3984 ( .A1(n9865), .A2(n78), .B1(n14730), .B2(n79), .ZN(n10101) );
  OAI22_X1 U3985 ( .A1(n9849), .A2(n78), .B1(n14690), .B2(n79), .ZN(n10102) );
  OAI22_X1 U3986 ( .A1(n9833), .A2(n78), .B1(n14650), .B2(n79), .ZN(n10103) );
  OAI22_X1 U3987 ( .A1(n9817), .A2(n81), .B1(n14959), .B2(n82), .ZN(n10104) );
  OAI22_X1 U3988 ( .A1(n9801), .A2(n81), .B1(n14890), .B2(n82), .ZN(n10105) );
  OAI22_X1 U3989 ( .A1(n9785), .A2(n81), .B1(n14850), .B2(n82), .ZN(n10106) );
  OAI22_X1 U3990 ( .A1(n9769), .A2(n81), .B1(n14810), .B2(n82), .ZN(n10107) );
  OAI22_X1 U3991 ( .A1(n9753), .A2(n81), .B1(n14770), .B2(n82), .ZN(n10108) );
  OAI22_X1 U3992 ( .A1(n9737), .A2(n81), .B1(n14730), .B2(n82), .ZN(n10109) );
  OAI22_X1 U3993 ( .A1(n9721), .A2(n81), .B1(n14690), .B2(n82), .ZN(n10110) );
  OAI22_X1 U3994 ( .A1(n9705), .A2(n81), .B1(n14650), .B2(n82), .ZN(n10111) );
  OAI22_X1 U3995 ( .A1(n9689), .A2(n84), .B1(n14959), .B2(n85), .ZN(n10112) );
  OAI22_X1 U3996 ( .A1(n9673), .A2(n84), .B1(n14890), .B2(n85), .ZN(n10113) );
  OAI22_X1 U3997 ( .A1(n9657), .A2(n84), .B1(n14850), .B2(n85), .ZN(n10114) );
  OAI22_X1 U3998 ( .A1(n9641), .A2(n84), .B1(n14810), .B2(n85), .ZN(n10115) );
  OAI22_X1 U3999 ( .A1(n9625), .A2(n84), .B1(n14770), .B2(n85), .ZN(n10116) );
  OAI22_X1 U4000 ( .A1(n9609), .A2(n84), .B1(n14730), .B2(n85), .ZN(n10117) );
  OAI22_X1 U4001 ( .A1(n9593), .A2(n84), .B1(n14690), .B2(n85), .ZN(n10118) );
  OAI22_X1 U4002 ( .A1(n9577), .A2(n84), .B1(n14650), .B2(n85), .ZN(n10119) );
  OAI22_X1 U4003 ( .A1(n9561), .A2(n87), .B1(n14959), .B2(n88), .ZN(n10120) );
  OAI22_X1 U4004 ( .A1(n9545), .A2(n87), .B1(n14890), .B2(n88), .ZN(n10121) );
  OAI22_X1 U4005 ( .A1(n9529), .A2(n87), .B1(n14850), .B2(n88), .ZN(n10122) );
  OAI22_X1 U4006 ( .A1(n9513), .A2(n87), .B1(n14810), .B2(n88), .ZN(n10123) );
  OAI22_X1 U4007 ( .A1(n9497), .A2(n87), .B1(n14770), .B2(n88), .ZN(n10124) );
  OAI22_X1 U4008 ( .A1(n9481), .A2(n87), .B1(n14730), .B2(n88), .ZN(n10125) );
  OAI22_X1 U4009 ( .A1(n9465), .A2(n87), .B1(n14690), .B2(n88), .ZN(n10126) );
  OAI22_X1 U4010 ( .A1(n9449), .A2(n87), .B1(n14650), .B2(n88), .ZN(n10127) );
  OAI22_X1 U4011 ( .A1(n9433), .A2(n90), .B1(n14959), .B2(n91), .ZN(n10128) );
  OAI22_X1 U4012 ( .A1(n9417), .A2(n90), .B1(n14890), .B2(n91), .ZN(n10129) );
  OAI22_X1 U4013 ( .A1(n9401), .A2(n90), .B1(n14850), .B2(n91), .ZN(n10130) );
  OAI22_X1 U4014 ( .A1(n9385), .A2(n90), .B1(n14810), .B2(n91), .ZN(n10131) );
  OAI22_X1 U4015 ( .A1(n9369), .A2(n90), .B1(n14770), .B2(n91), .ZN(n10132) );
  OAI22_X1 U4016 ( .A1(n9353), .A2(n90), .B1(n14730), .B2(n91), .ZN(n10133) );
  OAI22_X1 U4017 ( .A1(n9337), .A2(n90), .B1(n14690), .B2(n91), .ZN(n10134) );
  OAI22_X1 U4018 ( .A1(n9321), .A2(n90), .B1(n14650), .B2(n91), .ZN(n10135) );
  OAI22_X1 U4019 ( .A1(n10057), .A2(n66), .B1(n14890), .B2(n67), .ZN(n10089)
         );
  OAI22_X1 U4020 ( .A1(n10041), .A2(n66), .B1(n14850), .B2(n67), .ZN(n10090)
         );
  OAI22_X1 U4021 ( .A1(n10025), .A2(n66), .B1(n14810), .B2(n67), .ZN(n10091)
         );
  OAI22_X1 U4022 ( .A1(n10009), .A2(n66), .B1(n14770), .B2(n67), .ZN(n10092)
         );
  OAI22_X1 U4023 ( .A1(n9993), .A2(n66), .B1(n14730), .B2(n67), .ZN(n10093) );
  OAI22_X1 U4024 ( .A1(n9977), .A2(n66), .B1(n14690), .B2(n67), .ZN(n10094) );
  OAI22_X1 U4025 ( .A1(n9961), .A2(n66), .B1(n14650), .B2(n67), .ZN(n10095) );
  OAI22_X1 U4026 ( .A1(n7641), .A2(n132), .B1(n14958), .B2(n133), .ZN(n10240)
         );
  OAI22_X1 U4027 ( .A1(n7625), .A2(n132), .B1(n14891), .B2(n133), .ZN(n10241)
         );
  OAI22_X1 U4028 ( .A1(n7609), .A2(n132), .B1(n14851), .B2(n133), .ZN(n10242)
         );
  OAI22_X1 U4029 ( .A1(n7593), .A2(n132), .B1(n14811), .B2(n133), .ZN(n10243)
         );
  OAI22_X1 U4030 ( .A1(n7577), .A2(n132), .B1(n14771), .B2(n133), .ZN(n10244)
         );
  OAI22_X1 U4031 ( .A1(n7561), .A2(n132), .B1(n14731), .B2(n133), .ZN(n10245)
         );
  OAI22_X1 U4032 ( .A1(n7545), .A2(n132), .B1(n14691), .B2(n133), .ZN(n10246)
         );
  OAI22_X1 U4033 ( .A1(n7529), .A2(n132), .B1(n14651), .B2(n133), .ZN(n10247)
         );
  OAI22_X1 U4034 ( .A1(n7513), .A2(n135), .B1(n14958), .B2(n136), .ZN(n10248)
         );
  OAI22_X1 U4035 ( .A1(n7497), .A2(n135), .B1(n14891), .B2(n136), .ZN(n10249)
         );
  OAI22_X1 U4036 ( .A1(n7481), .A2(n135), .B1(n14851), .B2(n136), .ZN(n10250)
         );
  OAI22_X1 U4037 ( .A1(n7465), .A2(n135), .B1(n14811), .B2(n136), .ZN(n10251)
         );
  OAI22_X1 U4038 ( .A1(n7449), .A2(n135), .B1(n14771), .B2(n136), .ZN(n10252)
         );
  OAI22_X1 U4039 ( .A1(n7433), .A2(n135), .B1(n14731), .B2(n136), .ZN(n10253)
         );
  OAI22_X1 U4040 ( .A1(n7417), .A2(n135), .B1(n14691), .B2(n136), .ZN(n10254)
         );
  OAI22_X1 U4041 ( .A1(n7401), .A2(n135), .B1(n14651), .B2(n136), .ZN(n10255)
         );
  OAI22_X1 U4042 ( .A1(n7385), .A2(n138), .B1(n14957), .B2(n139), .ZN(n10256)
         );
  OAI22_X1 U4043 ( .A1(n7369), .A2(n138), .B1(n14891), .B2(n139), .ZN(n10257)
         );
  OAI22_X1 U4044 ( .A1(n7353), .A2(n138), .B1(n14851), .B2(n139), .ZN(n10258)
         );
  OAI22_X1 U4045 ( .A1(n7337), .A2(n138), .B1(n14811), .B2(n139), .ZN(n10259)
         );
  OAI22_X1 U4046 ( .A1(n7321), .A2(n138), .B1(n14771), .B2(n139), .ZN(n10260)
         );
  OAI22_X1 U4047 ( .A1(n7305), .A2(n138), .B1(n14731), .B2(n139), .ZN(n10261)
         );
  OAI22_X1 U4048 ( .A1(n7289), .A2(n138), .B1(n14691), .B2(n139), .ZN(n10262)
         );
  OAI22_X1 U4049 ( .A1(n7273), .A2(n138), .B1(n14651), .B2(n139), .ZN(n10263)
         );
  OAI22_X1 U4050 ( .A1(n7257), .A2(n141), .B1(n14957), .B2(n142), .ZN(n10264)
         );
  OAI22_X1 U4051 ( .A1(n7241), .A2(n141), .B1(n14891), .B2(n142), .ZN(n10265)
         );
  OAI22_X1 U4052 ( .A1(n7225), .A2(n141), .B1(n14851), .B2(n142), .ZN(n10266)
         );
  OAI22_X1 U4053 ( .A1(n7209), .A2(n141), .B1(n14811), .B2(n142), .ZN(n10267)
         );
  OAI22_X1 U4054 ( .A1(n7193), .A2(n141), .B1(n14771), .B2(n142), .ZN(n10268)
         );
  OAI22_X1 U4055 ( .A1(n7177), .A2(n141), .B1(n14731), .B2(n142), .ZN(n10269)
         );
  OAI22_X1 U4056 ( .A1(n7161), .A2(n141), .B1(n14691), .B2(n142), .ZN(n10270)
         );
  OAI22_X1 U4057 ( .A1(n7145), .A2(n141), .B1(n14651), .B2(n142), .ZN(n10271)
         );
  OAI22_X1 U4058 ( .A1(n7129), .A2(n144), .B1(n14957), .B2(n145), .ZN(n10272)
         );
  OAI22_X1 U4059 ( .A1(n7113), .A2(n144), .B1(n14891), .B2(n145), .ZN(n10273)
         );
  OAI22_X1 U4060 ( .A1(n7097), .A2(n144), .B1(n14851), .B2(n145), .ZN(n10274)
         );
  OAI22_X1 U4061 ( .A1(n7081), .A2(n144), .B1(n14811), .B2(n145), .ZN(n10275)
         );
  OAI22_X1 U4062 ( .A1(n7065), .A2(n144), .B1(n14771), .B2(n145), .ZN(n10276)
         );
  OAI22_X1 U4063 ( .A1(n7049), .A2(n144), .B1(n14731), .B2(n145), .ZN(n10277)
         );
  OAI22_X1 U4064 ( .A1(n7033), .A2(n144), .B1(n14691), .B2(n145), .ZN(n10278)
         );
  OAI22_X1 U4065 ( .A1(n7017), .A2(n144), .B1(n14651), .B2(n145), .ZN(n10279)
         );
  OAI22_X1 U4066 ( .A1(n7001), .A2(n147), .B1(n14957), .B2(n148), .ZN(n10280)
         );
  OAI22_X1 U4067 ( .A1(n6985), .A2(n147), .B1(n14891), .B2(n148), .ZN(n10281)
         );
  OAI22_X1 U4068 ( .A1(n6969), .A2(n147), .B1(n14851), .B2(n148), .ZN(n10282)
         );
  OAI22_X1 U4069 ( .A1(n6953), .A2(n147), .B1(n14811), .B2(n148), .ZN(n10283)
         );
  OAI22_X1 U4070 ( .A1(n6937), .A2(n147), .B1(n14771), .B2(n148), .ZN(n10284)
         );
  OAI22_X1 U4071 ( .A1(n6921), .A2(n147), .B1(n14731), .B2(n148), .ZN(n10285)
         );
  OAI22_X1 U4072 ( .A1(n6905), .A2(n147), .B1(n14691), .B2(n148), .ZN(n10286)
         );
  OAI22_X1 U4073 ( .A1(n6889), .A2(n147), .B1(n14651), .B2(n148), .ZN(n10287)
         );
  OAI22_X1 U4074 ( .A1(n6873), .A2(n150), .B1(n14957), .B2(n151), .ZN(n10288)
         );
  OAI22_X1 U4075 ( .A1(n6857), .A2(n150), .B1(n14891), .B2(n151), .ZN(n10289)
         );
  OAI22_X1 U4076 ( .A1(n6841), .A2(n150), .B1(n14851), .B2(n151), .ZN(n10290)
         );
  OAI22_X1 U4077 ( .A1(n6825), .A2(n150), .B1(n14811), .B2(n151), .ZN(n10291)
         );
  OAI22_X1 U4078 ( .A1(n6809), .A2(n150), .B1(n14771), .B2(n151), .ZN(n10292)
         );
  OAI22_X1 U4079 ( .A1(n6793), .A2(n150), .B1(n14731), .B2(n151), .ZN(n10293)
         );
  OAI22_X1 U4080 ( .A1(n6777), .A2(n150), .B1(n14691), .B2(n151), .ZN(n10294)
         );
  OAI22_X1 U4081 ( .A1(n6761), .A2(n150), .B1(n14651), .B2(n151), .ZN(n10295)
         );
  OAI22_X1 U4082 ( .A1(n6745), .A2(n153), .B1(n14957), .B2(n154), .ZN(n10296)
         );
  OAI22_X1 U4083 ( .A1(n6729), .A2(n153), .B1(n14892), .B2(n154), .ZN(n10297)
         );
  OAI22_X1 U4084 ( .A1(n6713), .A2(n153), .B1(n14852), .B2(n154), .ZN(n10298)
         );
  OAI22_X1 U4085 ( .A1(n6697), .A2(n153), .B1(n14812), .B2(n154), .ZN(n10299)
         );
  OAI22_X1 U4086 ( .A1(n6681), .A2(n153), .B1(n14772), .B2(n154), .ZN(n10300)
         );
  OAI22_X1 U4087 ( .A1(n6665), .A2(n153), .B1(n14732), .B2(n154), .ZN(n10301)
         );
  OAI22_X1 U4088 ( .A1(n6649), .A2(n153), .B1(n14692), .B2(n154), .ZN(n10302)
         );
  OAI22_X1 U4089 ( .A1(n6633), .A2(n153), .B1(n14652), .B2(n154), .ZN(n10303)
         );
  OAI22_X1 U4090 ( .A1(n6617), .A2(n156), .B1(n14957), .B2(n157), .ZN(n10304)
         );
  OAI22_X1 U4091 ( .A1(n6601), .A2(n156), .B1(n14892), .B2(n157), .ZN(n10305)
         );
  OAI22_X1 U4092 ( .A1(n6585), .A2(n156), .B1(n14852), .B2(n157), .ZN(n10306)
         );
  OAI22_X1 U4093 ( .A1(n6569), .A2(n156), .B1(n14812), .B2(n157), .ZN(n10307)
         );
  OAI22_X1 U4094 ( .A1(n6553), .A2(n156), .B1(n14772), .B2(n157), .ZN(n10308)
         );
  OAI22_X1 U4095 ( .A1(n6537), .A2(n156), .B1(n14732), .B2(n157), .ZN(n10309)
         );
  OAI22_X1 U4096 ( .A1(n6521), .A2(n156), .B1(n14692), .B2(n157), .ZN(n10310)
         );
  OAI22_X1 U4097 ( .A1(n6505), .A2(n156), .B1(n14652), .B2(n157), .ZN(n10311)
         );
  OAI22_X1 U4098 ( .A1(n6489), .A2(n159), .B1(n14957), .B2(n160), .ZN(n10312)
         );
  OAI22_X1 U4099 ( .A1(n6473), .A2(n159), .B1(n14892), .B2(n160), .ZN(n10313)
         );
  OAI22_X1 U4100 ( .A1(n6457), .A2(n159), .B1(n14852), .B2(n160), .ZN(n10314)
         );
  OAI22_X1 U4101 ( .A1(n6441), .A2(n159), .B1(n14812), .B2(n160), .ZN(n10315)
         );
  OAI22_X1 U4102 ( .A1(n6425), .A2(n159), .B1(n14772), .B2(n160), .ZN(n10316)
         );
  OAI22_X1 U4103 ( .A1(n6409), .A2(n159), .B1(n14732), .B2(n160), .ZN(n10317)
         );
  OAI22_X1 U4104 ( .A1(n6393), .A2(n159), .B1(n14692), .B2(n160), .ZN(n10318)
         );
  OAI22_X1 U4105 ( .A1(n6377), .A2(n159), .B1(n14652), .B2(n160), .ZN(n10319)
         );
  OAI22_X1 U4106 ( .A1(n6361), .A2(n162), .B1(n14957), .B2(n163), .ZN(n10320)
         );
  OAI22_X1 U4107 ( .A1(n6345), .A2(n162), .B1(n14892), .B2(n163), .ZN(n10321)
         );
  OAI22_X1 U4108 ( .A1(n6329), .A2(n162), .B1(n14852), .B2(n163), .ZN(n10322)
         );
  OAI22_X1 U4109 ( .A1(n6313), .A2(n162), .B1(n14812), .B2(n163), .ZN(n10323)
         );
  OAI22_X1 U4110 ( .A1(n6297), .A2(n162), .B1(n14772), .B2(n163), .ZN(n10324)
         );
  OAI22_X1 U4111 ( .A1(n6281), .A2(n162), .B1(n14732), .B2(n163), .ZN(n10325)
         );
  OAI22_X1 U4112 ( .A1(n6265), .A2(n162), .B1(n14692), .B2(n163), .ZN(n10326)
         );
  OAI22_X1 U4113 ( .A1(n6249), .A2(n162), .B1(n14652), .B2(n163), .ZN(n10327)
         );
  OAI22_X1 U4114 ( .A1(n6233), .A2(n165), .B1(n14957), .B2(n166), .ZN(n10328)
         );
  OAI22_X1 U4115 ( .A1(n6217), .A2(n165), .B1(n14892), .B2(n166), .ZN(n10329)
         );
  OAI22_X1 U4116 ( .A1(n6201), .A2(n165), .B1(n14852), .B2(n166), .ZN(n10330)
         );
  OAI22_X1 U4117 ( .A1(n6185), .A2(n165), .B1(n14812), .B2(n166), .ZN(n10331)
         );
  OAI22_X1 U4118 ( .A1(n6169), .A2(n165), .B1(n14772), .B2(n166), .ZN(n10332)
         );
  OAI22_X1 U4119 ( .A1(n6153), .A2(n165), .B1(n14732), .B2(n166), .ZN(n10333)
         );
  OAI22_X1 U4120 ( .A1(n6137), .A2(n165), .B1(n14692), .B2(n166), .ZN(n10334)
         );
  OAI22_X1 U4121 ( .A1(n6121), .A2(n165), .B1(n14652), .B2(n166), .ZN(n10335)
         );
  OAI22_X1 U4122 ( .A1(n6105), .A2(n168), .B1(n14957), .B2(n169), .ZN(n10336)
         );
  OAI22_X1 U4123 ( .A1(n6089), .A2(n168), .B1(n14892), .B2(n169), .ZN(n10337)
         );
  OAI22_X1 U4124 ( .A1(n6073), .A2(n168), .B1(n14852), .B2(n169), .ZN(n10338)
         );
  OAI22_X1 U4125 ( .A1(n6057), .A2(n168), .B1(n14812), .B2(n169), .ZN(n10339)
         );
  OAI22_X1 U4126 ( .A1(n6041), .A2(n168), .B1(n14772), .B2(n169), .ZN(n10340)
         );
  OAI22_X1 U4127 ( .A1(n6025), .A2(n168), .B1(n14732), .B2(n169), .ZN(n10341)
         );
  OAI22_X1 U4128 ( .A1(n6009), .A2(n168), .B1(n14692), .B2(n169), .ZN(n10342)
         );
  OAI22_X1 U4129 ( .A1(n5993), .A2(n168), .B1(n14652), .B2(n169), .ZN(n10343)
         );
  OAI22_X1 U4130 ( .A1(n9305), .A2(n93), .B1(n14959), .B2(n94), .ZN(n10136) );
  OAI22_X1 U4131 ( .A1(n9289), .A2(n93), .B1(n14890), .B2(n94), .ZN(n10137) );
  OAI22_X1 U4132 ( .A1(n9273), .A2(n93), .B1(n14850), .B2(n94), .ZN(n10138) );
  OAI22_X1 U4133 ( .A1(n9257), .A2(n93), .B1(n14810), .B2(n94), .ZN(n10139) );
  OAI22_X1 U4134 ( .A1(n9241), .A2(n93), .B1(n14770), .B2(n94), .ZN(n10140) );
  OAI22_X1 U4135 ( .A1(n9225), .A2(n93), .B1(n14730), .B2(n94), .ZN(n10141) );
  OAI22_X1 U4136 ( .A1(n9209), .A2(n93), .B1(n14690), .B2(n94), .ZN(n10142) );
  OAI22_X1 U4137 ( .A1(n9193), .A2(n93), .B1(n14650), .B2(n94), .ZN(n10143) );
  OAI22_X1 U4138 ( .A1(n9177), .A2(n96), .B1(n14959), .B2(n97), .ZN(n10144) );
  OAI22_X1 U4139 ( .A1(n9161), .A2(n96), .B1(n14890), .B2(n97), .ZN(n10145) );
  OAI22_X1 U4140 ( .A1(n9145), .A2(n96), .B1(n14850), .B2(n97), .ZN(n10146) );
  OAI22_X1 U4141 ( .A1(n9129), .A2(n96), .B1(n14810), .B2(n97), .ZN(n10147) );
  OAI22_X1 U4142 ( .A1(n9113), .A2(n96), .B1(n14770), .B2(n97), .ZN(n10148) );
  OAI22_X1 U4143 ( .A1(n9097), .A2(n96), .B1(n14730), .B2(n97), .ZN(n10149) );
  OAI22_X1 U4144 ( .A1(n9081), .A2(n96), .B1(n14690), .B2(n97), .ZN(n10150) );
  OAI22_X1 U4145 ( .A1(n9065), .A2(n96), .B1(n14650), .B2(n97), .ZN(n10151) );
  OAI22_X1 U4146 ( .A1(n9049), .A2(n99), .B1(n14958), .B2(n100), .ZN(n10152)
         );
  OAI22_X1 U4147 ( .A1(n9033), .A2(n99), .B1(n14890), .B2(n100), .ZN(n10153)
         );
  OAI22_X1 U4148 ( .A1(n9017), .A2(n99), .B1(n14850), .B2(n100), .ZN(n10154)
         );
  OAI22_X1 U4149 ( .A1(n9001), .A2(n99), .B1(n14810), .B2(n100), .ZN(n10155)
         );
  OAI22_X1 U4150 ( .A1(n8985), .A2(n99), .B1(n14770), .B2(n100), .ZN(n10156)
         );
  OAI22_X1 U4151 ( .A1(n8969), .A2(n99), .B1(n14730), .B2(n100), .ZN(n10157)
         );
  OAI22_X1 U4152 ( .A1(n8953), .A2(n99), .B1(n14690), .B2(n100), .ZN(n10158)
         );
  OAI22_X1 U4153 ( .A1(n8937), .A2(n99), .B1(n14650), .B2(n100), .ZN(n10159)
         );
  OAI22_X1 U4154 ( .A1(n8921), .A2(n102), .B1(n14958), .B2(n103), .ZN(n10160)
         );
  OAI22_X1 U4155 ( .A1(n8905), .A2(n102), .B1(n14890), .B2(n103), .ZN(n10161)
         );
  OAI22_X1 U4156 ( .A1(n8889), .A2(n102), .B1(n14850), .B2(n103), .ZN(n10162)
         );
  OAI22_X1 U4157 ( .A1(n8873), .A2(n102), .B1(n14810), .B2(n103), .ZN(n10163)
         );
  OAI22_X1 U4158 ( .A1(n8857), .A2(n102), .B1(n14770), .B2(n103), .ZN(n10164)
         );
  OAI22_X1 U4159 ( .A1(n8841), .A2(n102), .B1(n14730), .B2(n103), .ZN(n10165)
         );
  OAI22_X1 U4160 ( .A1(n8825), .A2(n102), .B1(n14690), .B2(n103), .ZN(n10166)
         );
  OAI22_X1 U4161 ( .A1(n8809), .A2(n102), .B1(n14650), .B2(n103), .ZN(n10167)
         );
  OAI22_X1 U4162 ( .A1(n8793), .A2(n105), .B1(n14958), .B2(n106), .ZN(n10168)
         );
  OAI22_X1 U4163 ( .A1(n8777), .A2(n105), .B1(n14890), .B2(n106), .ZN(n10169)
         );
  OAI22_X1 U4164 ( .A1(n8761), .A2(n105), .B1(n14850), .B2(n106), .ZN(n10170)
         );
  OAI22_X1 U4165 ( .A1(n8745), .A2(n105), .B1(n14810), .B2(n106), .ZN(n10171)
         );
  OAI22_X1 U4166 ( .A1(n8729), .A2(n105), .B1(n14770), .B2(n106), .ZN(n10172)
         );
  OAI22_X1 U4167 ( .A1(n8713), .A2(n105), .B1(n14730), .B2(n106), .ZN(n10173)
         );
  OAI22_X1 U4168 ( .A1(n8697), .A2(n105), .B1(n14690), .B2(n106), .ZN(n10174)
         );
  OAI22_X1 U4169 ( .A1(n8681), .A2(n105), .B1(n14650), .B2(n106), .ZN(n10175)
         );
  OAI22_X1 U4170 ( .A1(n8665), .A2(n108), .B1(n14958), .B2(n109), .ZN(n10176)
         );
  OAI22_X1 U4171 ( .A1(n8649), .A2(n108), .B1(n14890), .B2(n109), .ZN(n10177)
         );
  OAI22_X1 U4172 ( .A1(n8633), .A2(n108), .B1(n14850), .B2(n109), .ZN(n10178)
         );
  OAI22_X1 U4173 ( .A1(n8617), .A2(n108), .B1(n14810), .B2(n109), .ZN(n10179)
         );
  OAI22_X1 U4174 ( .A1(n8601), .A2(n108), .B1(n14770), .B2(n109), .ZN(n10180)
         );
  OAI22_X1 U4175 ( .A1(n8585), .A2(n108), .B1(n14730), .B2(n109), .ZN(n10181)
         );
  OAI22_X1 U4176 ( .A1(n8569), .A2(n108), .B1(n14690), .B2(n109), .ZN(n10182)
         );
  OAI22_X1 U4177 ( .A1(n8553), .A2(n108), .B1(n14650), .B2(n109), .ZN(n10183)
         );
  OAI22_X1 U4178 ( .A1(n8537), .A2(n111), .B1(n14958), .B2(n112), .ZN(n10184)
         );
  OAI22_X1 U4179 ( .A1(n8521), .A2(n111), .B1(n14890), .B2(n112), .ZN(n10185)
         );
  OAI22_X1 U4180 ( .A1(n8505), .A2(n111), .B1(n14850), .B2(n112), .ZN(n10186)
         );
  OAI22_X1 U4181 ( .A1(n8489), .A2(n111), .B1(n14810), .B2(n112), .ZN(n10187)
         );
  OAI22_X1 U4182 ( .A1(n8473), .A2(n111), .B1(n14770), .B2(n112), .ZN(n10188)
         );
  OAI22_X1 U4183 ( .A1(n8457), .A2(n111), .B1(n14730), .B2(n112), .ZN(n10189)
         );
  OAI22_X1 U4184 ( .A1(n8441), .A2(n111), .B1(n14690), .B2(n112), .ZN(n10190)
         );
  OAI22_X1 U4185 ( .A1(n8425), .A2(n111), .B1(n14650), .B2(n112), .ZN(n10191)
         );
  OAI22_X1 U4186 ( .A1(n8409), .A2(n114), .B1(n14958), .B2(n115), .ZN(n10192)
         );
  OAI22_X1 U4187 ( .A1(n8393), .A2(n114), .B1(n14891), .B2(n115), .ZN(n10193)
         );
  OAI22_X1 U4188 ( .A1(n8377), .A2(n114), .B1(n14851), .B2(n115), .ZN(n10194)
         );
  OAI22_X1 U4189 ( .A1(n8361), .A2(n114), .B1(n14811), .B2(n115), .ZN(n10195)
         );
  OAI22_X1 U4190 ( .A1(n8345), .A2(n114), .B1(n14771), .B2(n115), .ZN(n10196)
         );
  OAI22_X1 U4191 ( .A1(n8329), .A2(n114), .B1(n14731), .B2(n115), .ZN(n10197)
         );
  OAI22_X1 U4192 ( .A1(n8313), .A2(n114), .B1(n14691), .B2(n115), .ZN(n10198)
         );
  OAI22_X1 U4193 ( .A1(n8297), .A2(n114), .B1(n14651), .B2(n115), .ZN(n10199)
         );
  OAI22_X1 U4194 ( .A1(n8281), .A2(n117), .B1(n14958), .B2(n118), .ZN(n10200)
         );
  OAI22_X1 U4195 ( .A1(n8265), .A2(n117), .B1(n14891), .B2(n118), .ZN(n10201)
         );
  OAI22_X1 U4196 ( .A1(n8249), .A2(n117), .B1(n14851), .B2(n118), .ZN(n10202)
         );
  OAI22_X1 U4197 ( .A1(n8233), .A2(n117), .B1(n14811), .B2(n118), .ZN(n10203)
         );
  OAI22_X1 U4198 ( .A1(n8217), .A2(n117), .B1(n14771), .B2(n118), .ZN(n10204)
         );
  OAI22_X1 U4199 ( .A1(n8201), .A2(n117), .B1(n14731), .B2(n118), .ZN(n10205)
         );
  OAI22_X1 U4200 ( .A1(n8185), .A2(n117), .B1(n14691), .B2(n118), .ZN(n10206)
         );
  OAI22_X1 U4201 ( .A1(n8169), .A2(n117), .B1(n14651), .B2(n118), .ZN(n10207)
         );
  OAI22_X1 U4202 ( .A1(n8153), .A2(n120), .B1(n14958), .B2(n121), .ZN(n10208)
         );
  OAI22_X1 U4203 ( .A1(n8137), .A2(n120), .B1(n14891), .B2(n121), .ZN(n10209)
         );
  OAI22_X1 U4204 ( .A1(n8121), .A2(n120), .B1(n14851), .B2(n121), .ZN(n10210)
         );
  OAI22_X1 U4205 ( .A1(n8105), .A2(n120), .B1(n14811), .B2(n121), .ZN(n10211)
         );
  OAI22_X1 U4206 ( .A1(n8089), .A2(n120), .B1(n14771), .B2(n121), .ZN(n10212)
         );
  OAI22_X1 U4207 ( .A1(n8073), .A2(n120), .B1(n14731), .B2(n121), .ZN(n10213)
         );
  OAI22_X1 U4208 ( .A1(n8057), .A2(n120), .B1(n14691), .B2(n121), .ZN(n10214)
         );
  OAI22_X1 U4209 ( .A1(n8041), .A2(n120), .B1(n14651), .B2(n121), .ZN(n10215)
         );
  OAI22_X1 U4210 ( .A1(n8025), .A2(n123), .B1(n14958), .B2(n124), .ZN(n10216)
         );
  OAI22_X1 U4211 ( .A1(n8009), .A2(n123), .B1(n14891), .B2(n124), .ZN(n10217)
         );
  OAI22_X1 U4212 ( .A1(n7993), .A2(n123), .B1(n14851), .B2(n124), .ZN(n10218)
         );
  OAI22_X1 U4213 ( .A1(n7977), .A2(n123), .B1(n14811), .B2(n124), .ZN(n10219)
         );
  OAI22_X1 U4214 ( .A1(n7961), .A2(n123), .B1(n14771), .B2(n124), .ZN(n10220)
         );
  OAI22_X1 U4215 ( .A1(n7945), .A2(n123), .B1(n14731), .B2(n124), .ZN(n10221)
         );
  OAI22_X1 U4216 ( .A1(n7929), .A2(n123), .B1(n14691), .B2(n124), .ZN(n10222)
         );
  OAI22_X1 U4217 ( .A1(n7913), .A2(n123), .B1(n14651), .B2(n124), .ZN(n10223)
         );
  OAI22_X1 U4218 ( .A1(n7897), .A2(n126), .B1(n14958), .B2(n127), .ZN(n10224)
         );
  OAI22_X1 U4219 ( .A1(n7881), .A2(n126), .B1(n14891), .B2(n127), .ZN(n10225)
         );
  OAI22_X1 U4220 ( .A1(n7865), .A2(n126), .B1(n14851), .B2(n127), .ZN(n10226)
         );
  OAI22_X1 U4221 ( .A1(n7849), .A2(n126), .B1(n14811), .B2(n127), .ZN(n10227)
         );
  OAI22_X1 U4222 ( .A1(n7833), .A2(n126), .B1(n14771), .B2(n127), .ZN(n10228)
         );
  OAI22_X1 U4223 ( .A1(n7817), .A2(n126), .B1(n14731), .B2(n127), .ZN(n10229)
         );
  OAI22_X1 U4224 ( .A1(n7801), .A2(n126), .B1(n14691), .B2(n127), .ZN(n10230)
         );
  OAI22_X1 U4225 ( .A1(n7785), .A2(n126), .B1(n14651), .B2(n127), .ZN(n10231)
         );
  OAI22_X1 U4226 ( .A1(n7769), .A2(n129), .B1(n14958), .B2(n130), .ZN(n10232)
         );
  OAI22_X1 U4227 ( .A1(n7753), .A2(n129), .B1(n14891), .B2(n130), .ZN(n10233)
         );
  OAI22_X1 U4228 ( .A1(n7737), .A2(n129), .B1(n14851), .B2(n130), .ZN(n10234)
         );
  OAI22_X1 U4229 ( .A1(n7721), .A2(n129), .B1(n14811), .B2(n130), .ZN(n10235)
         );
  OAI22_X1 U4230 ( .A1(n7705), .A2(n129), .B1(n14771), .B2(n130), .ZN(n10236)
         );
  OAI22_X1 U4231 ( .A1(n7689), .A2(n129), .B1(n14731), .B2(n130), .ZN(n10237)
         );
  OAI22_X1 U4232 ( .A1(n7673), .A2(n129), .B1(n14691), .B2(n130), .ZN(n10238)
         );
  OAI22_X1 U4233 ( .A1(n7657), .A2(n129), .B1(n14651), .B2(n130), .ZN(n10239)
         );
  OAI22_X1 U4234 ( .A1(n10077), .A2(n173), .B1(n14957), .B2(n174), .ZN(n10344)
         );
  OAI22_X1 U4235 ( .A1(n10061), .A2(n173), .B1(n14892), .B2(n174), .ZN(n10345)
         );
  OAI22_X1 U4236 ( .A1(n10045), .A2(n173), .B1(n14852), .B2(n174), .ZN(n10346)
         );
  OAI22_X1 U4237 ( .A1(n10029), .A2(n173), .B1(n14812), .B2(n174), .ZN(n10347)
         );
  OAI22_X1 U4238 ( .A1(n10013), .A2(n173), .B1(n14772), .B2(n174), .ZN(n10348)
         );
  OAI22_X1 U4239 ( .A1(n9997), .A2(n173), .B1(n14732), .B2(n174), .ZN(n10349)
         );
  OAI22_X1 U4240 ( .A1(n9981), .A2(n173), .B1(n14692), .B2(n174), .ZN(n10350)
         );
  OAI22_X1 U4241 ( .A1(n9965), .A2(n173), .B1(n14652), .B2(n174), .ZN(n10351)
         );
  OAI22_X1 U4242 ( .A1(n9949), .A2(n176), .B1(n14957), .B2(n177), .ZN(n10352)
         );
  OAI22_X1 U4243 ( .A1(n9933), .A2(n176), .B1(n14892), .B2(n177), .ZN(n10353)
         );
  OAI22_X1 U4244 ( .A1(n9917), .A2(n176), .B1(n14852), .B2(n177), .ZN(n10354)
         );
  OAI22_X1 U4245 ( .A1(n9901), .A2(n176), .B1(n14812), .B2(n177), .ZN(n10355)
         );
  OAI22_X1 U4246 ( .A1(n9885), .A2(n176), .B1(n14772), .B2(n177), .ZN(n10356)
         );
  OAI22_X1 U4247 ( .A1(n9869), .A2(n176), .B1(n14732), .B2(n177), .ZN(n10357)
         );
  OAI22_X1 U4248 ( .A1(n9853), .A2(n176), .B1(n14692), .B2(n177), .ZN(n10358)
         );
  OAI22_X1 U4249 ( .A1(n9837), .A2(n176), .B1(n14652), .B2(n177), .ZN(n10359)
         );
  OAI22_X1 U4250 ( .A1(n9821), .A2(n178), .B1(n14956), .B2(n179), .ZN(n10360)
         );
  OAI22_X1 U4251 ( .A1(n9805), .A2(n178), .B1(n14892), .B2(n179), .ZN(n10361)
         );
  OAI22_X1 U4252 ( .A1(n9789), .A2(n178), .B1(n14852), .B2(n179), .ZN(n10362)
         );
  OAI22_X1 U4253 ( .A1(n9773), .A2(n178), .B1(n14812), .B2(n179), .ZN(n10363)
         );
  OAI22_X1 U4254 ( .A1(n9757), .A2(n178), .B1(n14772), .B2(n179), .ZN(n10364)
         );
  OAI22_X1 U4255 ( .A1(n9741), .A2(n178), .B1(n14732), .B2(n179), .ZN(n10365)
         );
  OAI22_X1 U4256 ( .A1(n9725), .A2(n178), .B1(n14692), .B2(n179), .ZN(n10366)
         );
  OAI22_X1 U4257 ( .A1(n9709), .A2(n178), .B1(n14652), .B2(n179), .ZN(n10367)
         );
  OAI22_X1 U4258 ( .A1(n9693), .A2(n180), .B1(n14956), .B2(n181), .ZN(n10368)
         );
  OAI22_X1 U4259 ( .A1(n9677), .A2(n180), .B1(n14892), .B2(n181), .ZN(n10369)
         );
  OAI22_X1 U4260 ( .A1(n9661), .A2(n180), .B1(n14852), .B2(n181), .ZN(n10370)
         );
  OAI22_X1 U4261 ( .A1(n9645), .A2(n180), .B1(n14812), .B2(n181), .ZN(n10371)
         );
  OAI22_X1 U4262 ( .A1(n9629), .A2(n180), .B1(n14772), .B2(n181), .ZN(n10372)
         );
  OAI22_X1 U4263 ( .A1(n9613), .A2(n180), .B1(n14732), .B2(n181), .ZN(n10373)
         );
  OAI22_X1 U4264 ( .A1(n9597), .A2(n180), .B1(n14692), .B2(n181), .ZN(n10374)
         );
  OAI22_X1 U4265 ( .A1(n9581), .A2(n180), .B1(n14652), .B2(n181), .ZN(n10375)
         );
  OAI22_X1 U4266 ( .A1(n9565), .A2(n182), .B1(n14956), .B2(n183), .ZN(n10376)
         );
  OAI22_X1 U4267 ( .A1(n9549), .A2(n182), .B1(n14892), .B2(n183), .ZN(n10377)
         );
  OAI22_X1 U4268 ( .A1(n9533), .A2(n182), .B1(n14852), .B2(n183), .ZN(n10378)
         );
  OAI22_X1 U4269 ( .A1(n9517), .A2(n182), .B1(n14812), .B2(n183), .ZN(n10379)
         );
  OAI22_X1 U4270 ( .A1(n9501), .A2(n182), .B1(n14772), .B2(n183), .ZN(n10380)
         );
  OAI22_X1 U4271 ( .A1(n9485), .A2(n182), .B1(n14732), .B2(n183), .ZN(n10381)
         );
  OAI22_X1 U4272 ( .A1(n9469), .A2(n182), .B1(n14692), .B2(n183), .ZN(n10382)
         );
  OAI22_X1 U4273 ( .A1(n9453), .A2(n182), .B1(n14652), .B2(n183), .ZN(n10383)
         );
  OAI22_X1 U4274 ( .A1(n9437), .A2(n184), .B1(n14956), .B2(n185), .ZN(n10384)
         );
  OAI22_X1 U4275 ( .A1(n9421), .A2(n184), .B1(n14892), .B2(n185), .ZN(n10385)
         );
  OAI22_X1 U4276 ( .A1(n9405), .A2(n184), .B1(n14852), .B2(n185), .ZN(n10386)
         );
  OAI22_X1 U4277 ( .A1(n9389), .A2(n184), .B1(n14812), .B2(n185), .ZN(n10387)
         );
  OAI22_X1 U4278 ( .A1(n9373), .A2(n184), .B1(n14772), .B2(n185), .ZN(n10388)
         );
  OAI22_X1 U4279 ( .A1(n9357), .A2(n184), .B1(n14732), .B2(n185), .ZN(n10389)
         );
  OAI22_X1 U4280 ( .A1(n9341), .A2(n184), .B1(n14692), .B2(n185), .ZN(n10390)
         );
  OAI22_X1 U4281 ( .A1(n9325), .A2(n184), .B1(n14652), .B2(n185), .ZN(n10391)
         );
  OAI22_X1 U4282 ( .A1(n9309), .A2(n186), .B1(n14956), .B2(n187), .ZN(n10392)
         );
  OAI22_X1 U4283 ( .A1(n9293), .A2(n186), .B1(n14892), .B2(n187), .ZN(n10393)
         );
  OAI22_X1 U4284 ( .A1(n9277), .A2(n186), .B1(n14852), .B2(n187), .ZN(n10394)
         );
  OAI22_X1 U4285 ( .A1(n9261), .A2(n186), .B1(n14812), .B2(n187), .ZN(n10395)
         );
  OAI22_X1 U4286 ( .A1(n9245), .A2(n186), .B1(n14772), .B2(n187), .ZN(n10396)
         );
  OAI22_X1 U4287 ( .A1(n9229), .A2(n186), .B1(n14732), .B2(n187), .ZN(n10397)
         );
  OAI22_X1 U4288 ( .A1(n9213), .A2(n186), .B1(n14692), .B2(n187), .ZN(n10398)
         );
  OAI22_X1 U4289 ( .A1(n9197), .A2(n186), .B1(n14652), .B2(n187), .ZN(n10399)
         );
  OAI22_X1 U4290 ( .A1(n9181), .A2(n188), .B1(n14956), .B2(n189), .ZN(n10400)
         );
  OAI22_X1 U4291 ( .A1(n9165), .A2(n188), .B1(n14893), .B2(n189), .ZN(n10401)
         );
  OAI22_X1 U4292 ( .A1(n9149), .A2(n188), .B1(n14853), .B2(n189), .ZN(n10402)
         );
  OAI22_X1 U4293 ( .A1(n9133), .A2(n188), .B1(n14813), .B2(n189), .ZN(n10403)
         );
  OAI22_X1 U4294 ( .A1(n9117), .A2(n188), .B1(n14773), .B2(n189), .ZN(n10404)
         );
  OAI22_X1 U4295 ( .A1(n9101), .A2(n188), .B1(n14733), .B2(n189), .ZN(n10405)
         );
  OAI22_X1 U4296 ( .A1(n9085), .A2(n188), .B1(n14693), .B2(n189), .ZN(n10406)
         );
  OAI22_X1 U4297 ( .A1(n9069), .A2(n188), .B1(n14653), .B2(n189), .ZN(n10407)
         );
  OAI22_X1 U4298 ( .A1(n9053), .A2(n190), .B1(n14956), .B2(n191), .ZN(n10408)
         );
  OAI22_X1 U4299 ( .A1(n9037), .A2(n190), .B1(n14893), .B2(n191), .ZN(n10409)
         );
  OAI22_X1 U4300 ( .A1(n9021), .A2(n190), .B1(n14853), .B2(n191), .ZN(n10410)
         );
  OAI22_X1 U4301 ( .A1(n9005), .A2(n190), .B1(n14813), .B2(n191), .ZN(n10411)
         );
  OAI22_X1 U4302 ( .A1(n8989), .A2(n190), .B1(n14773), .B2(n191), .ZN(n10412)
         );
  OAI22_X1 U4303 ( .A1(n8973), .A2(n190), .B1(n14733), .B2(n191), .ZN(n10413)
         );
  OAI22_X1 U4304 ( .A1(n8957), .A2(n190), .B1(n14693), .B2(n191), .ZN(n10414)
         );
  OAI22_X1 U4305 ( .A1(n8941), .A2(n190), .B1(n14653), .B2(n191), .ZN(n10415)
         );
  OAI22_X1 U4306 ( .A1(n8925), .A2(n192), .B1(n14956), .B2(n193), .ZN(n10416)
         );
  OAI22_X1 U4307 ( .A1(n8909), .A2(n192), .B1(n14893), .B2(n193), .ZN(n10417)
         );
  OAI22_X1 U4308 ( .A1(n8893), .A2(n192), .B1(n14853), .B2(n193), .ZN(n10418)
         );
  OAI22_X1 U4309 ( .A1(n8877), .A2(n192), .B1(n14813), .B2(n193), .ZN(n10419)
         );
  OAI22_X1 U4310 ( .A1(n8861), .A2(n192), .B1(n14773), .B2(n193), .ZN(n10420)
         );
  OAI22_X1 U4311 ( .A1(n8845), .A2(n192), .B1(n14733), .B2(n193), .ZN(n10421)
         );
  OAI22_X1 U4312 ( .A1(n8829), .A2(n192), .B1(n14693), .B2(n193), .ZN(n10422)
         );
  OAI22_X1 U4313 ( .A1(n8813), .A2(n192), .B1(n14653), .B2(n193), .ZN(n10423)
         );
  OAI22_X1 U4314 ( .A1(n8797), .A2(n194), .B1(n14956), .B2(n195), .ZN(n10424)
         );
  OAI22_X1 U4315 ( .A1(n8781), .A2(n194), .B1(n14893), .B2(n195), .ZN(n10425)
         );
  OAI22_X1 U4316 ( .A1(n8765), .A2(n194), .B1(n14853), .B2(n195), .ZN(n10426)
         );
  OAI22_X1 U4317 ( .A1(n8749), .A2(n194), .B1(n14813), .B2(n195), .ZN(n10427)
         );
  OAI22_X1 U4318 ( .A1(n8733), .A2(n194), .B1(n14773), .B2(n195), .ZN(n10428)
         );
  OAI22_X1 U4319 ( .A1(n8717), .A2(n194), .B1(n14733), .B2(n195), .ZN(n10429)
         );
  OAI22_X1 U4320 ( .A1(n8701), .A2(n194), .B1(n14693), .B2(n195), .ZN(n10430)
         );
  OAI22_X1 U4321 ( .A1(n8685), .A2(n194), .B1(n14653), .B2(n195), .ZN(n10431)
         );
  OAI22_X1 U4322 ( .A1(n8669), .A2(n196), .B1(n14956), .B2(n197), .ZN(n10432)
         );
  OAI22_X1 U4323 ( .A1(n8653), .A2(n196), .B1(n14893), .B2(n197), .ZN(n10433)
         );
  OAI22_X1 U4324 ( .A1(n8637), .A2(n196), .B1(n14853), .B2(n197), .ZN(n10434)
         );
  OAI22_X1 U4325 ( .A1(n8621), .A2(n196), .B1(n14813), .B2(n197), .ZN(n10435)
         );
  OAI22_X1 U4326 ( .A1(n8605), .A2(n196), .B1(n14773), .B2(n197), .ZN(n10436)
         );
  OAI22_X1 U4327 ( .A1(n8589), .A2(n196), .B1(n14733), .B2(n197), .ZN(n10437)
         );
  OAI22_X1 U4328 ( .A1(n8573), .A2(n196), .B1(n14693), .B2(n197), .ZN(n10438)
         );
  OAI22_X1 U4329 ( .A1(n8557), .A2(n196), .B1(n14653), .B2(n197), .ZN(n10439)
         );
  OAI22_X1 U4330 ( .A1(n8541), .A2(n198), .B1(n14956), .B2(n199), .ZN(n10440)
         );
  OAI22_X1 U4331 ( .A1(n8525), .A2(n198), .B1(n14893), .B2(n199), .ZN(n10441)
         );
  OAI22_X1 U4332 ( .A1(n8509), .A2(n198), .B1(n14853), .B2(n199), .ZN(n10442)
         );
  OAI22_X1 U4333 ( .A1(n8493), .A2(n198), .B1(n14813), .B2(n199), .ZN(n10443)
         );
  OAI22_X1 U4334 ( .A1(n8477), .A2(n198), .B1(n14773), .B2(n199), .ZN(n10444)
         );
  OAI22_X1 U4335 ( .A1(n8461), .A2(n198), .B1(n14733), .B2(n199), .ZN(n10445)
         );
  OAI22_X1 U4336 ( .A1(n8445), .A2(n198), .B1(n14693), .B2(n199), .ZN(n10446)
         );
  OAI22_X1 U4337 ( .A1(n8429), .A2(n198), .B1(n14653), .B2(n199), .ZN(n10447)
         );
  OAI22_X1 U4338 ( .A1(n8413), .A2(n200), .B1(n14956), .B2(n201), .ZN(n10448)
         );
  OAI22_X1 U4339 ( .A1(n8397), .A2(n200), .B1(n14893), .B2(n201), .ZN(n10449)
         );
  OAI22_X1 U4340 ( .A1(n8381), .A2(n200), .B1(n14853), .B2(n201), .ZN(n10450)
         );
  OAI22_X1 U4341 ( .A1(n8365), .A2(n200), .B1(n14813), .B2(n201), .ZN(n10451)
         );
  OAI22_X1 U4342 ( .A1(n8349), .A2(n200), .B1(n14773), .B2(n201), .ZN(n10452)
         );
  OAI22_X1 U4343 ( .A1(n8333), .A2(n200), .B1(n14733), .B2(n201), .ZN(n10453)
         );
  OAI22_X1 U4344 ( .A1(n8317), .A2(n200), .B1(n14693), .B2(n201), .ZN(n10454)
         );
  OAI22_X1 U4345 ( .A1(n8301), .A2(n200), .B1(n14653), .B2(n201), .ZN(n10455)
         );
  OAI22_X1 U4346 ( .A1(n8285), .A2(n202), .B1(n14956), .B2(n203), .ZN(n10456)
         );
  OAI22_X1 U4347 ( .A1(n8269), .A2(n202), .B1(n14893), .B2(n203), .ZN(n10457)
         );
  OAI22_X1 U4348 ( .A1(n8253), .A2(n202), .B1(n14853), .B2(n203), .ZN(n10458)
         );
  OAI22_X1 U4349 ( .A1(n8237), .A2(n202), .B1(n14813), .B2(n203), .ZN(n10459)
         );
  OAI22_X1 U4350 ( .A1(n8221), .A2(n202), .B1(n14773), .B2(n203), .ZN(n10460)
         );
  OAI22_X1 U4351 ( .A1(n8205), .A2(n202), .B1(n14733), .B2(n203), .ZN(n10461)
         );
  OAI22_X1 U4352 ( .A1(n8189), .A2(n202), .B1(n14693), .B2(n203), .ZN(n10462)
         );
  OAI22_X1 U4353 ( .A1(n8173), .A2(n202), .B1(n14653), .B2(n203), .ZN(n10463)
         );
  OAI22_X1 U4354 ( .A1(n8157), .A2(n204), .B1(n14955), .B2(n205), .ZN(n10464)
         );
  OAI22_X1 U4355 ( .A1(n8141), .A2(n204), .B1(n14893), .B2(n205), .ZN(n10465)
         );
  OAI22_X1 U4356 ( .A1(n8125), .A2(n204), .B1(n14853), .B2(n205), .ZN(n10466)
         );
  OAI22_X1 U4357 ( .A1(n8109), .A2(n204), .B1(n14813), .B2(n205), .ZN(n10467)
         );
  OAI22_X1 U4358 ( .A1(n8093), .A2(n204), .B1(n14773), .B2(n205), .ZN(n10468)
         );
  OAI22_X1 U4359 ( .A1(n8077), .A2(n204), .B1(n14733), .B2(n205), .ZN(n10469)
         );
  OAI22_X1 U4360 ( .A1(n8061), .A2(n204), .B1(n14693), .B2(n205), .ZN(n10470)
         );
  OAI22_X1 U4361 ( .A1(n8045), .A2(n204), .B1(n14653), .B2(n205), .ZN(n10471)
         );
  OAI22_X1 U4362 ( .A1(n8029), .A2(n206), .B1(n14955), .B2(n207), .ZN(n10472)
         );
  OAI22_X1 U4363 ( .A1(n8013), .A2(n206), .B1(n14893), .B2(n207), .ZN(n10473)
         );
  OAI22_X1 U4364 ( .A1(n7997), .A2(n206), .B1(n14853), .B2(n207), .ZN(n10474)
         );
  OAI22_X1 U4365 ( .A1(n7981), .A2(n206), .B1(n14813), .B2(n207), .ZN(n10475)
         );
  OAI22_X1 U4366 ( .A1(n7965), .A2(n206), .B1(n14773), .B2(n207), .ZN(n10476)
         );
  OAI22_X1 U4367 ( .A1(n7949), .A2(n206), .B1(n14733), .B2(n207), .ZN(n10477)
         );
  OAI22_X1 U4368 ( .A1(n7933), .A2(n206), .B1(n14693), .B2(n207), .ZN(n10478)
         );
  OAI22_X1 U4369 ( .A1(n7917), .A2(n206), .B1(n14653), .B2(n207), .ZN(n10479)
         );
  OAI22_X1 U4370 ( .A1(n7901), .A2(n208), .B1(n14955), .B2(n209), .ZN(n10480)
         );
  OAI22_X1 U4371 ( .A1(n7885), .A2(n208), .B1(n14893), .B2(n209), .ZN(n10481)
         );
  OAI22_X1 U4372 ( .A1(n7869), .A2(n208), .B1(n14853), .B2(n209), .ZN(n10482)
         );
  OAI22_X1 U4373 ( .A1(n7853), .A2(n208), .B1(n14813), .B2(n209), .ZN(n10483)
         );
  OAI22_X1 U4374 ( .A1(n7837), .A2(n208), .B1(n14773), .B2(n209), .ZN(n10484)
         );
  OAI22_X1 U4375 ( .A1(n7821), .A2(n208), .B1(n14733), .B2(n209), .ZN(n10485)
         );
  OAI22_X1 U4376 ( .A1(n7805), .A2(n208), .B1(n14693), .B2(n209), .ZN(n10486)
         );
  OAI22_X1 U4377 ( .A1(n7789), .A2(n208), .B1(n14653), .B2(n209), .ZN(n10487)
         );
  OAI22_X1 U4378 ( .A1(n7773), .A2(n210), .B1(n14955), .B2(n211), .ZN(n10488)
         );
  OAI22_X1 U4379 ( .A1(n7757), .A2(n210), .B1(n14893), .B2(n211), .ZN(n10489)
         );
  OAI22_X1 U4380 ( .A1(n7741), .A2(n210), .B1(n14853), .B2(n211), .ZN(n10490)
         );
  OAI22_X1 U4381 ( .A1(n7725), .A2(n210), .B1(n14813), .B2(n211), .ZN(n10491)
         );
  OAI22_X1 U4382 ( .A1(n7709), .A2(n210), .B1(n14773), .B2(n211), .ZN(n10492)
         );
  OAI22_X1 U4383 ( .A1(n7693), .A2(n210), .B1(n14733), .B2(n211), .ZN(n10493)
         );
  OAI22_X1 U4384 ( .A1(n7677), .A2(n210), .B1(n14693), .B2(n211), .ZN(n10494)
         );
  OAI22_X1 U4385 ( .A1(n7661), .A2(n210), .B1(n14653), .B2(n211), .ZN(n10495)
         );
  OAI22_X1 U4386 ( .A1(n7645), .A2(n212), .B1(n14955), .B2(n213), .ZN(n10496)
         );
  OAI22_X1 U4387 ( .A1(n7629), .A2(n212), .B1(n14893), .B2(n213), .ZN(n10497)
         );
  OAI22_X1 U4388 ( .A1(n7613), .A2(n212), .B1(n14853), .B2(n213), .ZN(n10498)
         );
  OAI22_X1 U4389 ( .A1(n7597), .A2(n212), .B1(n14813), .B2(n213), .ZN(n10499)
         );
  OAI22_X1 U4390 ( .A1(n7581), .A2(n212), .B1(n14773), .B2(n213), .ZN(n10500)
         );
  OAI22_X1 U4391 ( .A1(n7565), .A2(n212), .B1(n14733), .B2(n213), .ZN(n10501)
         );
  OAI22_X1 U4392 ( .A1(n7549), .A2(n212), .B1(n14693), .B2(n213), .ZN(n10502)
         );
  OAI22_X1 U4393 ( .A1(n7533), .A2(n212), .B1(n14653), .B2(n213), .ZN(n10503)
         );
  OAI22_X1 U4394 ( .A1(n7517), .A2(n214), .B1(n14955), .B2(n215), .ZN(n10504)
         );
  OAI22_X1 U4395 ( .A1(n7501), .A2(n214), .B1(n14894), .B2(n215), .ZN(n10505)
         );
  OAI22_X1 U4396 ( .A1(n7485), .A2(n214), .B1(n14854), .B2(n215), .ZN(n10506)
         );
  OAI22_X1 U4397 ( .A1(n7469), .A2(n214), .B1(n14814), .B2(n215), .ZN(n10507)
         );
  OAI22_X1 U4398 ( .A1(n7453), .A2(n214), .B1(n14774), .B2(n215), .ZN(n10508)
         );
  OAI22_X1 U4399 ( .A1(n7437), .A2(n214), .B1(n14734), .B2(n215), .ZN(n10509)
         );
  OAI22_X1 U4400 ( .A1(n7421), .A2(n214), .B1(n14694), .B2(n215), .ZN(n10510)
         );
  OAI22_X1 U4401 ( .A1(n7405), .A2(n214), .B1(n14654), .B2(n215), .ZN(n10511)
         );
  OAI22_X1 U4402 ( .A1(n7389), .A2(n216), .B1(n14955), .B2(n217), .ZN(n10512)
         );
  OAI22_X1 U4403 ( .A1(n7373), .A2(n216), .B1(n14894), .B2(n217), .ZN(n10513)
         );
  OAI22_X1 U4404 ( .A1(n7357), .A2(n216), .B1(n14854), .B2(n217), .ZN(n10514)
         );
  OAI22_X1 U4405 ( .A1(n7341), .A2(n216), .B1(n14814), .B2(n217), .ZN(n10515)
         );
  OAI22_X1 U4406 ( .A1(n7325), .A2(n216), .B1(n14774), .B2(n217), .ZN(n10516)
         );
  OAI22_X1 U4407 ( .A1(n7309), .A2(n216), .B1(n14734), .B2(n217), .ZN(n10517)
         );
  OAI22_X1 U4408 ( .A1(n7293), .A2(n216), .B1(n14694), .B2(n217), .ZN(n10518)
         );
  OAI22_X1 U4409 ( .A1(n7277), .A2(n216), .B1(n14654), .B2(n217), .ZN(n10519)
         );
  OAI22_X1 U4410 ( .A1(n7261), .A2(n218), .B1(n14955), .B2(n219), .ZN(n10520)
         );
  OAI22_X1 U4411 ( .A1(n7245), .A2(n218), .B1(n14894), .B2(n219), .ZN(n10521)
         );
  OAI22_X1 U4412 ( .A1(n7229), .A2(n218), .B1(n14854), .B2(n219), .ZN(n10522)
         );
  OAI22_X1 U4413 ( .A1(n7213), .A2(n218), .B1(n14814), .B2(n219), .ZN(n10523)
         );
  OAI22_X1 U4414 ( .A1(n7197), .A2(n218), .B1(n14774), .B2(n219), .ZN(n10524)
         );
  OAI22_X1 U4415 ( .A1(n7181), .A2(n218), .B1(n14734), .B2(n219), .ZN(n10525)
         );
  OAI22_X1 U4416 ( .A1(n7165), .A2(n218), .B1(n14694), .B2(n219), .ZN(n10526)
         );
  OAI22_X1 U4417 ( .A1(n7149), .A2(n218), .B1(n14654), .B2(n219), .ZN(n10527)
         );
  OAI22_X1 U4418 ( .A1(n7133), .A2(n220), .B1(n14955), .B2(n221), .ZN(n10528)
         );
  OAI22_X1 U4419 ( .A1(n7117), .A2(n220), .B1(n14894), .B2(n221), .ZN(n10529)
         );
  OAI22_X1 U4420 ( .A1(n7101), .A2(n220), .B1(n14854), .B2(n221), .ZN(n10530)
         );
  OAI22_X1 U4421 ( .A1(n7085), .A2(n220), .B1(n14814), .B2(n221), .ZN(n10531)
         );
  OAI22_X1 U4422 ( .A1(n7069), .A2(n220), .B1(n14774), .B2(n221), .ZN(n10532)
         );
  OAI22_X1 U4423 ( .A1(n7053), .A2(n220), .B1(n14734), .B2(n221), .ZN(n10533)
         );
  OAI22_X1 U4424 ( .A1(n7037), .A2(n220), .B1(n14694), .B2(n221), .ZN(n10534)
         );
  OAI22_X1 U4425 ( .A1(n7021), .A2(n220), .B1(n14654), .B2(n221), .ZN(n10535)
         );
  OAI22_X1 U4426 ( .A1(n7005), .A2(n222), .B1(n14955), .B2(n223), .ZN(n10536)
         );
  OAI22_X1 U4427 ( .A1(n6989), .A2(n222), .B1(n14894), .B2(n223), .ZN(n10537)
         );
  OAI22_X1 U4428 ( .A1(n6973), .A2(n222), .B1(n14854), .B2(n223), .ZN(n10538)
         );
  OAI22_X1 U4429 ( .A1(n6957), .A2(n222), .B1(n14814), .B2(n223), .ZN(n10539)
         );
  OAI22_X1 U4430 ( .A1(n6941), .A2(n222), .B1(n14774), .B2(n223), .ZN(n10540)
         );
  OAI22_X1 U4431 ( .A1(n6925), .A2(n222), .B1(n14734), .B2(n223), .ZN(n10541)
         );
  OAI22_X1 U4432 ( .A1(n6909), .A2(n222), .B1(n14694), .B2(n223), .ZN(n10542)
         );
  OAI22_X1 U4433 ( .A1(n6893), .A2(n222), .B1(n14654), .B2(n223), .ZN(n10543)
         );
  OAI22_X1 U4434 ( .A1(n6877), .A2(n224), .B1(n14955), .B2(n225), .ZN(n10544)
         );
  OAI22_X1 U4435 ( .A1(n6861), .A2(n224), .B1(n14894), .B2(n225), .ZN(n10545)
         );
  OAI22_X1 U4436 ( .A1(n6845), .A2(n224), .B1(n14854), .B2(n225), .ZN(n10546)
         );
  OAI22_X1 U4437 ( .A1(n6829), .A2(n224), .B1(n14814), .B2(n225), .ZN(n10547)
         );
  OAI22_X1 U4438 ( .A1(n6813), .A2(n224), .B1(n14774), .B2(n225), .ZN(n10548)
         );
  OAI22_X1 U4439 ( .A1(n6797), .A2(n224), .B1(n14734), .B2(n225), .ZN(n10549)
         );
  OAI22_X1 U4440 ( .A1(n6781), .A2(n224), .B1(n14694), .B2(n225), .ZN(n10550)
         );
  OAI22_X1 U4441 ( .A1(n6765), .A2(n224), .B1(n14654), .B2(n225), .ZN(n10551)
         );
  OAI22_X1 U4442 ( .A1(n10085), .A2(n305), .B1(n14952), .B2(n306), .ZN(n10856)
         );
  OAI22_X1 U4443 ( .A1(n10069), .A2(n305), .B1(n14897), .B2(n306), .ZN(n10857)
         );
  OAI22_X1 U4444 ( .A1(n10053), .A2(n305), .B1(n14857), .B2(n306), .ZN(n10858)
         );
  OAI22_X1 U4445 ( .A1(n10037), .A2(n305), .B1(n14817), .B2(n306), .ZN(n10859)
         );
  OAI22_X1 U4446 ( .A1(n10021), .A2(n305), .B1(n14777), .B2(n306), .ZN(n10860)
         );
  OAI22_X1 U4447 ( .A1(n10005), .A2(n305), .B1(n14737), .B2(n306), .ZN(n10861)
         );
  OAI22_X1 U4448 ( .A1(n9989), .A2(n305), .B1(n14697), .B2(n306), .ZN(n10862)
         );
  OAI22_X1 U4449 ( .A1(n9973), .A2(n305), .B1(n14657), .B2(n306), .ZN(n10863)
         );
  OAI22_X1 U4450 ( .A1(n9957), .A2(n308), .B1(n14952), .B2(n309), .ZN(n10864)
         );
  OAI22_X1 U4451 ( .A1(n9941), .A2(n308), .B1(n14897), .B2(n309), .ZN(n10865)
         );
  OAI22_X1 U4452 ( .A1(n9925), .A2(n308), .B1(n14857), .B2(n309), .ZN(n10866)
         );
  OAI22_X1 U4453 ( .A1(n9909), .A2(n308), .B1(n14817), .B2(n309), .ZN(n10867)
         );
  OAI22_X1 U4454 ( .A1(n9893), .A2(n308), .B1(n14777), .B2(n309), .ZN(n10868)
         );
  OAI22_X1 U4455 ( .A1(n9877), .A2(n308), .B1(n14737), .B2(n309), .ZN(n10869)
         );
  OAI22_X1 U4456 ( .A1(n9861), .A2(n308), .B1(n14697), .B2(n309), .ZN(n10870)
         );
  OAI22_X1 U4457 ( .A1(n9845), .A2(n308), .B1(n14657), .B2(n309), .ZN(n10871)
         );
  OAI22_X1 U4458 ( .A1(n9829), .A2(n310), .B1(n14951), .B2(n311), .ZN(n10872)
         );
  OAI22_X1 U4459 ( .A1(n9813), .A2(n310), .B1(n14897), .B2(n311), .ZN(n10873)
         );
  OAI22_X1 U4460 ( .A1(n9797), .A2(n310), .B1(n14857), .B2(n311), .ZN(n10874)
         );
  OAI22_X1 U4461 ( .A1(n9781), .A2(n310), .B1(n14817), .B2(n311), .ZN(n10875)
         );
  OAI22_X1 U4462 ( .A1(n9765), .A2(n310), .B1(n14777), .B2(n311), .ZN(n10876)
         );
  OAI22_X1 U4463 ( .A1(n9749), .A2(n310), .B1(n14737), .B2(n311), .ZN(n10877)
         );
  OAI22_X1 U4464 ( .A1(n9733), .A2(n310), .B1(n14697), .B2(n311), .ZN(n10878)
         );
  OAI22_X1 U4465 ( .A1(n9717), .A2(n310), .B1(n14657), .B2(n311), .ZN(n10879)
         );
  OAI22_X1 U4466 ( .A1(n9701), .A2(n312), .B1(n14951), .B2(n313), .ZN(n10880)
         );
  OAI22_X1 U4467 ( .A1(n9685), .A2(n312), .B1(n14897), .B2(n313), .ZN(n10881)
         );
  OAI22_X1 U4468 ( .A1(n9669), .A2(n312), .B1(n14857), .B2(n313), .ZN(n10882)
         );
  OAI22_X1 U4469 ( .A1(n9653), .A2(n312), .B1(n14817), .B2(n313), .ZN(n10883)
         );
  OAI22_X1 U4470 ( .A1(n9637), .A2(n312), .B1(n14777), .B2(n313), .ZN(n10884)
         );
  OAI22_X1 U4471 ( .A1(n9621), .A2(n312), .B1(n14737), .B2(n313), .ZN(n10885)
         );
  OAI22_X1 U4472 ( .A1(n9605), .A2(n312), .B1(n14697), .B2(n313), .ZN(n10886)
         );
  OAI22_X1 U4473 ( .A1(n9589), .A2(n312), .B1(n14657), .B2(n313), .ZN(n10887)
         );
  OAI22_X1 U4474 ( .A1(n9573), .A2(n314), .B1(n14951), .B2(n315), .ZN(n10888)
         );
  OAI22_X1 U4475 ( .A1(n9557), .A2(n314), .B1(n14897), .B2(n315), .ZN(n10889)
         );
  OAI22_X1 U4476 ( .A1(n9541), .A2(n314), .B1(n14857), .B2(n315), .ZN(n10890)
         );
  OAI22_X1 U4477 ( .A1(n9525), .A2(n314), .B1(n14817), .B2(n315), .ZN(n10891)
         );
  OAI22_X1 U4478 ( .A1(n9509), .A2(n314), .B1(n14777), .B2(n315), .ZN(n10892)
         );
  OAI22_X1 U4479 ( .A1(n9493), .A2(n314), .B1(n14737), .B2(n315), .ZN(n10893)
         );
  OAI22_X1 U4480 ( .A1(n9477), .A2(n314), .B1(n14697), .B2(n315), .ZN(n10894)
         );
  OAI22_X1 U4481 ( .A1(n9461), .A2(n314), .B1(n14657), .B2(n315), .ZN(n10895)
         );
  OAI22_X1 U4482 ( .A1(n9445), .A2(n316), .B1(n14951), .B2(n317), .ZN(n10896)
         );
  OAI22_X1 U4483 ( .A1(n9429), .A2(n316), .B1(n14897), .B2(n317), .ZN(n10897)
         );
  OAI22_X1 U4484 ( .A1(n9413), .A2(n316), .B1(n14857), .B2(n317), .ZN(n10898)
         );
  OAI22_X1 U4485 ( .A1(n9397), .A2(n316), .B1(n14817), .B2(n317), .ZN(n10899)
         );
  OAI22_X1 U4486 ( .A1(n9381), .A2(n316), .B1(n14777), .B2(n317), .ZN(n10900)
         );
  OAI22_X1 U4487 ( .A1(n9365), .A2(n316), .B1(n14737), .B2(n317), .ZN(n10901)
         );
  OAI22_X1 U4488 ( .A1(n9349), .A2(n316), .B1(n14697), .B2(n317), .ZN(n10902)
         );
  OAI22_X1 U4489 ( .A1(n9333), .A2(n316), .B1(n14657), .B2(n317), .ZN(n10903)
         );
  OAI22_X1 U4490 ( .A1(n9317), .A2(n318), .B1(n14951), .B2(n319), .ZN(n10904)
         );
  OAI22_X1 U4491 ( .A1(n9301), .A2(n318), .B1(n14897), .B2(n319), .ZN(n10905)
         );
  OAI22_X1 U4492 ( .A1(n9285), .A2(n318), .B1(n14857), .B2(n319), .ZN(n10906)
         );
  OAI22_X1 U4493 ( .A1(n9269), .A2(n318), .B1(n14817), .B2(n319), .ZN(n10907)
         );
  OAI22_X1 U4494 ( .A1(n9253), .A2(n318), .B1(n14777), .B2(n319), .ZN(n10908)
         );
  OAI22_X1 U4495 ( .A1(n9237), .A2(n318), .B1(n14737), .B2(n319), .ZN(n10909)
         );
  OAI22_X1 U4496 ( .A1(n9221), .A2(n318), .B1(n14697), .B2(n319), .ZN(n10910)
         );
  OAI22_X1 U4497 ( .A1(n9205), .A2(n318), .B1(n14657), .B2(n319), .ZN(n10911)
         );
  OAI22_X1 U4498 ( .A1(n9189), .A2(n320), .B1(n14951), .B2(n321), .ZN(n10912)
         );
  OAI22_X1 U4499 ( .A1(n9173), .A2(n320), .B1(n14897), .B2(n321), .ZN(n10913)
         );
  OAI22_X1 U4500 ( .A1(n9157), .A2(n320), .B1(n14857), .B2(n321), .ZN(n10914)
         );
  OAI22_X1 U4501 ( .A1(n9141), .A2(n320), .B1(n14817), .B2(n321), .ZN(n10915)
         );
  OAI22_X1 U4502 ( .A1(n9125), .A2(n320), .B1(n14777), .B2(n321), .ZN(n10916)
         );
  OAI22_X1 U4503 ( .A1(n9109), .A2(n320), .B1(n14737), .B2(n321), .ZN(n10917)
         );
  OAI22_X1 U4504 ( .A1(n9093), .A2(n320), .B1(n14697), .B2(n321), .ZN(n10918)
         );
  OAI22_X1 U4505 ( .A1(n9077), .A2(n320), .B1(n14657), .B2(n321), .ZN(n10919)
         );
  OAI22_X1 U4506 ( .A1(n9061), .A2(n322), .B1(n14951), .B2(n323), .ZN(n10920)
         );
  OAI22_X1 U4507 ( .A1(n9045), .A2(n322), .B1(n14898), .B2(n323), .ZN(n10921)
         );
  OAI22_X1 U4508 ( .A1(n9029), .A2(n322), .B1(n14858), .B2(n323), .ZN(n10922)
         );
  OAI22_X1 U4509 ( .A1(n9013), .A2(n322), .B1(n14818), .B2(n323), .ZN(n10923)
         );
  OAI22_X1 U4510 ( .A1(n8997), .A2(n322), .B1(n14778), .B2(n323), .ZN(n10924)
         );
  OAI22_X1 U4511 ( .A1(n8981), .A2(n322), .B1(n14738), .B2(n323), .ZN(n10925)
         );
  OAI22_X1 U4512 ( .A1(n8965), .A2(n322), .B1(n14698), .B2(n323), .ZN(n10926)
         );
  OAI22_X1 U4513 ( .A1(n8949), .A2(n322), .B1(n14658), .B2(n323), .ZN(n10927)
         );
  OAI22_X1 U4514 ( .A1(n8933), .A2(n324), .B1(n14951), .B2(n325), .ZN(n10928)
         );
  OAI22_X1 U4515 ( .A1(n8917), .A2(n324), .B1(n14898), .B2(n325), .ZN(n10929)
         );
  OAI22_X1 U4516 ( .A1(n8901), .A2(n324), .B1(n14858), .B2(n325), .ZN(n10930)
         );
  OAI22_X1 U4517 ( .A1(n8885), .A2(n324), .B1(n14818), .B2(n325), .ZN(n10931)
         );
  OAI22_X1 U4518 ( .A1(n8869), .A2(n324), .B1(n14778), .B2(n325), .ZN(n10932)
         );
  OAI22_X1 U4519 ( .A1(n8853), .A2(n324), .B1(n14738), .B2(n325), .ZN(n10933)
         );
  OAI22_X1 U4520 ( .A1(n8837), .A2(n324), .B1(n14698), .B2(n325), .ZN(n10934)
         );
  OAI22_X1 U4521 ( .A1(n8821), .A2(n324), .B1(n14658), .B2(n325), .ZN(n10935)
         );
  OAI22_X1 U4522 ( .A1(n8805), .A2(n326), .B1(n14951), .B2(n327), .ZN(n10936)
         );
  OAI22_X1 U4523 ( .A1(n8789), .A2(n326), .B1(n14898), .B2(n327), .ZN(n10937)
         );
  OAI22_X1 U4524 ( .A1(n8773), .A2(n326), .B1(n14858), .B2(n327), .ZN(n10938)
         );
  OAI22_X1 U4525 ( .A1(n8757), .A2(n326), .B1(n14818), .B2(n327), .ZN(n10939)
         );
  OAI22_X1 U4526 ( .A1(n8741), .A2(n326), .B1(n14778), .B2(n327), .ZN(n10940)
         );
  OAI22_X1 U4527 ( .A1(n8725), .A2(n326), .B1(n14738), .B2(n327), .ZN(n10941)
         );
  OAI22_X1 U4528 ( .A1(n8709), .A2(n326), .B1(n14698), .B2(n327), .ZN(n10942)
         );
  OAI22_X1 U4529 ( .A1(n8693), .A2(n326), .B1(n14658), .B2(n327), .ZN(n10943)
         );
  OAI22_X1 U4530 ( .A1(n8677), .A2(n328), .B1(n14951), .B2(n329), .ZN(n10944)
         );
  OAI22_X1 U4531 ( .A1(n8661), .A2(n328), .B1(n14898), .B2(n329), .ZN(n10945)
         );
  OAI22_X1 U4532 ( .A1(n8645), .A2(n328), .B1(n14858), .B2(n329), .ZN(n10946)
         );
  OAI22_X1 U4533 ( .A1(n8629), .A2(n328), .B1(n14818), .B2(n329), .ZN(n10947)
         );
  OAI22_X1 U4534 ( .A1(n8613), .A2(n328), .B1(n14778), .B2(n329), .ZN(n10948)
         );
  OAI22_X1 U4535 ( .A1(n8597), .A2(n328), .B1(n14738), .B2(n329), .ZN(n10949)
         );
  OAI22_X1 U4536 ( .A1(n8581), .A2(n328), .B1(n14698), .B2(n329), .ZN(n10950)
         );
  OAI22_X1 U4537 ( .A1(n8565), .A2(n328), .B1(n14658), .B2(n329), .ZN(n10951)
         );
  OAI22_X1 U4538 ( .A1(n8549), .A2(n330), .B1(n14951), .B2(n331), .ZN(n10952)
         );
  OAI22_X1 U4539 ( .A1(n8533), .A2(n330), .B1(n14898), .B2(n331), .ZN(n10953)
         );
  OAI22_X1 U4540 ( .A1(n8517), .A2(n330), .B1(n14858), .B2(n331), .ZN(n10954)
         );
  OAI22_X1 U4541 ( .A1(n8501), .A2(n330), .B1(n14818), .B2(n331), .ZN(n10955)
         );
  OAI22_X1 U4542 ( .A1(n8485), .A2(n330), .B1(n14778), .B2(n331), .ZN(n10956)
         );
  OAI22_X1 U4543 ( .A1(n8469), .A2(n330), .B1(n14738), .B2(n331), .ZN(n10957)
         );
  OAI22_X1 U4544 ( .A1(n8453), .A2(n330), .B1(n14698), .B2(n331), .ZN(n10958)
         );
  OAI22_X1 U4545 ( .A1(n8437), .A2(n330), .B1(n14658), .B2(n331), .ZN(n10959)
         );
  OAI22_X1 U4546 ( .A1(n8421), .A2(n332), .B1(n14951), .B2(n333), .ZN(n10960)
         );
  OAI22_X1 U4547 ( .A1(n8405), .A2(n332), .B1(n14898), .B2(n333), .ZN(n10961)
         );
  OAI22_X1 U4548 ( .A1(n8389), .A2(n332), .B1(n14858), .B2(n333), .ZN(n10962)
         );
  OAI22_X1 U4549 ( .A1(n8373), .A2(n332), .B1(n14818), .B2(n333), .ZN(n10963)
         );
  OAI22_X1 U4550 ( .A1(n8357), .A2(n332), .B1(n14778), .B2(n333), .ZN(n10964)
         );
  OAI22_X1 U4551 ( .A1(n8341), .A2(n332), .B1(n14738), .B2(n333), .ZN(n10965)
         );
  OAI22_X1 U4552 ( .A1(n8325), .A2(n332), .B1(n14698), .B2(n333), .ZN(n10966)
         );
  OAI22_X1 U4553 ( .A1(n8309), .A2(n332), .B1(n14658), .B2(n333), .ZN(n10967)
         );
  OAI22_X1 U4554 ( .A1(n8293), .A2(n334), .B1(n14951), .B2(n335), .ZN(n10968)
         );
  OAI22_X1 U4555 ( .A1(n8277), .A2(n334), .B1(n14898), .B2(n335), .ZN(n10969)
         );
  OAI22_X1 U4556 ( .A1(n8261), .A2(n334), .B1(n14858), .B2(n335), .ZN(n10970)
         );
  OAI22_X1 U4557 ( .A1(n8245), .A2(n334), .B1(n14818), .B2(n335), .ZN(n10971)
         );
  OAI22_X1 U4558 ( .A1(n8229), .A2(n334), .B1(n14778), .B2(n335), .ZN(n10972)
         );
  OAI22_X1 U4559 ( .A1(n8213), .A2(n334), .B1(n14738), .B2(n335), .ZN(n10973)
         );
  OAI22_X1 U4560 ( .A1(n8197), .A2(n334), .B1(n14698), .B2(n335), .ZN(n10974)
         );
  OAI22_X1 U4561 ( .A1(n8181), .A2(n334), .B1(n14658), .B2(n335), .ZN(n10975)
         );
  OAI22_X1 U4562 ( .A1(n8165), .A2(n336), .B1(n14950), .B2(n337), .ZN(n10976)
         );
  OAI22_X1 U4563 ( .A1(n8149), .A2(n336), .B1(n14898), .B2(n337), .ZN(n10977)
         );
  OAI22_X1 U4564 ( .A1(n8133), .A2(n336), .B1(n14858), .B2(n337), .ZN(n10978)
         );
  OAI22_X1 U4565 ( .A1(n8117), .A2(n336), .B1(n14818), .B2(n337), .ZN(n10979)
         );
  OAI22_X1 U4566 ( .A1(n8101), .A2(n336), .B1(n14778), .B2(n337), .ZN(n10980)
         );
  OAI22_X1 U4567 ( .A1(n8085), .A2(n336), .B1(n14738), .B2(n337), .ZN(n10981)
         );
  OAI22_X1 U4568 ( .A1(n8069), .A2(n336), .B1(n14698), .B2(n337), .ZN(n10982)
         );
  OAI22_X1 U4569 ( .A1(n8053), .A2(n336), .B1(n14658), .B2(n337), .ZN(n10983)
         );
  OAI22_X1 U4570 ( .A1(n8037), .A2(n338), .B1(n14950), .B2(n339), .ZN(n10984)
         );
  OAI22_X1 U4571 ( .A1(n8021), .A2(n338), .B1(n14898), .B2(n339), .ZN(n10985)
         );
  OAI22_X1 U4572 ( .A1(n8005), .A2(n338), .B1(n14858), .B2(n339), .ZN(n10986)
         );
  OAI22_X1 U4573 ( .A1(n7989), .A2(n338), .B1(n14818), .B2(n339), .ZN(n10987)
         );
  OAI22_X1 U4574 ( .A1(n7973), .A2(n338), .B1(n14778), .B2(n339), .ZN(n10988)
         );
  OAI22_X1 U4575 ( .A1(n7957), .A2(n338), .B1(n14738), .B2(n339), .ZN(n10989)
         );
  OAI22_X1 U4576 ( .A1(n7941), .A2(n338), .B1(n14698), .B2(n339), .ZN(n10990)
         );
  OAI22_X1 U4577 ( .A1(n7925), .A2(n338), .B1(n14658), .B2(n339), .ZN(n10991)
         );
  OAI22_X1 U4578 ( .A1(n7909), .A2(n340), .B1(n14950), .B2(n341), .ZN(n10992)
         );
  OAI22_X1 U4579 ( .A1(n7893), .A2(n340), .B1(n14898), .B2(n341), .ZN(n10993)
         );
  OAI22_X1 U4580 ( .A1(n7877), .A2(n340), .B1(n14858), .B2(n341), .ZN(n10994)
         );
  OAI22_X1 U4581 ( .A1(n7861), .A2(n340), .B1(n14818), .B2(n341), .ZN(n10995)
         );
  OAI22_X1 U4582 ( .A1(n7845), .A2(n340), .B1(n14778), .B2(n341), .ZN(n10996)
         );
  OAI22_X1 U4583 ( .A1(n7829), .A2(n340), .B1(n14738), .B2(n341), .ZN(n10997)
         );
  OAI22_X1 U4584 ( .A1(n7813), .A2(n340), .B1(n14698), .B2(n341), .ZN(n10998)
         );
  OAI22_X1 U4585 ( .A1(n7797), .A2(n340), .B1(n14658), .B2(n341), .ZN(n10999)
         );
  OAI22_X1 U4586 ( .A1(n7781), .A2(n342), .B1(n14950), .B2(n343), .ZN(n11000)
         );
  OAI22_X1 U4587 ( .A1(n7765), .A2(n342), .B1(n14898), .B2(n343), .ZN(n11001)
         );
  OAI22_X1 U4588 ( .A1(n7749), .A2(n342), .B1(n14858), .B2(n343), .ZN(n11002)
         );
  OAI22_X1 U4589 ( .A1(n7733), .A2(n342), .B1(n14818), .B2(n343), .ZN(n11003)
         );
  OAI22_X1 U4590 ( .A1(n7717), .A2(n342), .B1(n14778), .B2(n343), .ZN(n11004)
         );
  OAI22_X1 U4591 ( .A1(n7701), .A2(n342), .B1(n14738), .B2(n343), .ZN(n11005)
         );
  OAI22_X1 U4592 ( .A1(n7685), .A2(n342), .B1(n14698), .B2(n343), .ZN(n11006)
         );
  OAI22_X1 U4593 ( .A1(n7669), .A2(n342), .B1(n14658), .B2(n343), .ZN(n11007)
         );
  OAI22_X1 U4594 ( .A1(n7653), .A2(n344), .B1(n14950), .B2(n345), .ZN(n11008)
         );
  OAI22_X1 U4595 ( .A1(n7637), .A2(n344), .B1(n14898), .B2(n345), .ZN(n11009)
         );
  OAI22_X1 U4596 ( .A1(n7621), .A2(n344), .B1(n14858), .B2(n345), .ZN(n11010)
         );
  OAI22_X1 U4597 ( .A1(n7605), .A2(n344), .B1(n14818), .B2(n345), .ZN(n11011)
         );
  OAI22_X1 U4598 ( .A1(n7589), .A2(n344), .B1(n14778), .B2(n345), .ZN(n11012)
         );
  OAI22_X1 U4599 ( .A1(n7573), .A2(n344), .B1(n14738), .B2(n345), .ZN(n11013)
         );
  OAI22_X1 U4600 ( .A1(n7557), .A2(n344), .B1(n14698), .B2(n345), .ZN(n11014)
         );
  OAI22_X1 U4601 ( .A1(n7541), .A2(n344), .B1(n14658), .B2(n345), .ZN(n11015)
         );
  OAI22_X1 U4602 ( .A1(n7525), .A2(n346), .B1(n14950), .B2(n347), .ZN(n11016)
         );
  OAI22_X1 U4603 ( .A1(n7509), .A2(n346), .B1(n14898), .B2(n347), .ZN(n11017)
         );
  OAI22_X1 U4604 ( .A1(n7493), .A2(n346), .B1(n14858), .B2(n347), .ZN(n11018)
         );
  OAI22_X1 U4605 ( .A1(n7477), .A2(n346), .B1(n14818), .B2(n347), .ZN(n11019)
         );
  OAI22_X1 U4606 ( .A1(n7461), .A2(n346), .B1(n14778), .B2(n347), .ZN(n11020)
         );
  OAI22_X1 U4607 ( .A1(n7445), .A2(n346), .B1(n14738), .B2(n347), .ZN(n11021)
         );
  OAI22_X1 U4608 ( .A1(n7429), .A2(n346), .B1(n14698), .B2(n347), .ZN(n11022)
         );
  OAI22_X1 U4609 ( .A1(n7413), .A2(n346), .B1(n14658), .B2(n347), .ZN(n11023)
         );
  OAI22_X1 U4610 ( .A1(n7397), .A2(n348), .B1(n14950), .B2(n349), .ZN(n11024)
         );
  OAI22_X1 U4611 ( .A1(n7381), .A2(n348), .B1(n14899), .B2(n349), .ZN(n11025)
         );
  OAI22_X1 U4612 ( .A1(n7365), .A2(n348), .B1(n14859), .B2(n349), .ZN(n11026)
         );
  OAI22_X1 U4613 ( .A1(n7349), .A2(n348), .B1(n14819), .B2(n349), .ZN(n11027)
         );
  OAI22_X1 U4614 ( .A1(n7333), .A2(n348), .B1(n14779), .B2(n349), .ZN(n11028)
         );
  OAI22_X1 U4615 ( .A1(n7317), .A2(n348), .B1(n14739), .B2(n349), .ZN(n11029)
         );
  OAI22_X1 U4616 ( .A1(n7301), .A2(n348), .B1(n14699), .B2(n349), .ZN(n11030)
         );
  OAI22_X1 U4617 ( .A1(n7285), .A2(n348), .B1(n14659), .B2(n349), .ZN(n11031)
         );
  OAI22_X1 U4618 ( .A1(n7269), .A2(n350), .B1(n14950), .B2(n351), .ZN(n11032)
         );
  OAI22_X1 U4619 ( .A1(n7253), .A2(n350), .B1(n14899), .B2(n351), .ZN(n11033)
         );
  OAI22_X1 U4620 ( .A1(n7237), .A2(n350), .B1(n14859), .B2(n351), .ZN(n11034)
         );
  OAI22_X1 U4621 ( .A1(n7221), .A2(n350), .B1(n14819), .B2(n351), .ZN(n11035)
         );
  OAI22_X1 U4622 ( .A1(n7205), .A2(n350), .B1(n14779), .B2(n351), .ZN(n11036)
         );
  OAI22_X1 U4623 ( .A1(n7189), .A2(n350), .B1(n14739), .B2(n351), .ZN(n11037)
         );
  OAI22_X1 U4624 ( .A1(n7173), .A2(n350), .B1(n14699), .B2(n351), .ZN(n11038)
         );
  OAI22_X1 U4625 ( .A1(n7157), .A2(n350), .B1(n14659), .B2(n351), .ZN(n11039)
         );
  OAI22_X1 U4626 ( .A1(n7141), .A2(n352), .B1(n14950), .B2(n353), .ZN(n11040)
         );
  OAI22_X1 U4627 ( .A1(n7125), .A2(n352), .B1(n14899), .B2(n353), .ZN(n11041)
         );
  OAI22_X1 U4628 ( .A1(n7109), .A2(n352), .B1(n14859), .B2(n353), .ZN(n11042)
         );
  OAI22_X1 U4629 ( .A1(n7093), .A2(n352), .B1(n14819), .B2(n353), .ZN(n11043)
         );
  OAI22_X1 U4630 ( .A1(n7077), .A2(n352), .B1(n14779), .B2(n353), .ZN(n11044)
         );
  OAI22_X1 U4631 ( .A1(n7061), .A2(n352), .B1(n14739), .B2(n353), .ZN(n11045)
         );
  OAI22_X1 U4632 ( .A1(n7045), .A2(n352), .B1(n14699), .B2(n353), .ZN(n11046)
         );
  OAI22_X1 U4633 ( .A1(n7029), .A2(n352), .B1(n14659), .B2(n353), .ZN(n11047)
         );
  OAI22_X1 U4634 ( .A1(n7013), .A2(n354), .B1(n14950), .B2(n355), .ZN(n11048)
         );
  OAI22_X1 U4635 ( .A1(n6997), .A2(n354), .B1(n14899), .B2(n355), .ZN(n11049)
         );
  OAI22_X1 U4636 ( .A1(n6981), .A2(n354), .B1(n14859), .B2(n355), .ZN(n11050)
         );
  OAI22_X1 U4637 ( .A1(n6965), .A2(n354), .B1(n14819), .B2(n355), .ZN(n11051)
         );
  OAI22_X1 U4638 ( .A1(n6949), .A2(n354), .B1(n14779), .B2(n355), .ZN(n11052)
         );
  OAI22_X1 U4639 ( .A1(n6933), .A2(n354), .B1(n14739), .B2(n355), .ZN(n11053)
         );
  OAI22_X1 U4640 ( .A1(n6917), .A2(n354), .B1(n14699), .B2(n355), .ZN(n11054)
         );
  OAI22_X1 U4641 ( .A1(n6901), .A2(n354), .B1(n14659), .B2(n355), .ZN(n11055)
         );
  OAI22_X1 U4642 ( .A1(n6885), .A2(n356), .B1(n14950), .B2(n357), .ZN(n11056)
         );
  OAI22_X1 U4643 ( .A1(n6869), .A2(n356), .B1(n14899), .B2(n357), .ZN(n11057)
         );
  OAI22_X1 U4644 ( .A1(n6853), .A2(n356), .B1(n14859), .B2(n357), .ZN(n11058)
         );
  OAI22_X1 U4645 ( .A1(n6837), .A2(n356), .B1(n14819), .B2(n357), .ZN(n11059)
         );
  OAI22_X1 U4646 ( .A1(n6821), .A2(n356), .B1(n14779), .B2(n357), .ZN(n11060)
         );
  OAI22_X1 U4647 ( .A1(n6805), .A2(n356), .B1(n14739), .B2(n357), .ZN(n11061)
         );
  OAI22_X1 U4648 ( .A1(n6789), .A2(n356), .B1(n14699), .B2(n357), .ZN(n11062)
         );
  OAI22_X1 U4649 ( .A1(n6773), .A2(n356), .B1(n14659), .B2(n357), .ZN(n11063)
         );
  OAI22_X1 U4650 ( .A1(n9291), .A2(n384), .B1(n14900), .B2(n383), .ZN(n11161)
         );
  OAI22_X1 U4651 ( .A1(n9275), .A2(n384), .B1(n14860), .B2(n383), .ZN(n11162)
         );
  OAI22_X1 U4652 ( .A1(n9259), .A2(n384), .B1(n14820), .B2(n383), .ZN(n11163)
         );
  OAI22_X1 U4653 ( .A1(n9243), .A2(n384), .B1(n14780), .B2(n383), .ZN(n11164)
         );
  OAI22_X1 U4654 ( .A1(n9227), .A2(n384), .B1(n14740), .B2(n383), .ZN(n11165)
         );
  OAI22_X1 U4655 ( .A1(n9211), .A2(n384), .B1(n14700), .B2(n383), .ZN(n11166)
         );
  OAI22_X1 U4656 ( .A1(n9195), .A2(n384), .B1(n14660), .B2(n383), .ZN(n11167)
         );
  OAI22_X1 U4657 ( .A1(n9163), .A2(n386), .B1(n14900), .B2(n385), .ZN(n11169)
         );
  OAI22_X1 U4658 ( .A1(n9147), .A2(n386), .B1(n14860), .B2(n385), .ZN(n11170)
         );
  OAI22_X1 U4659 ( .A1(n9131), .A2(n386), .B1(n14820), .B2(n385), .ZN(n11171)
         );
  OAI22_X1 U4660 ( .A1(n9115), .A2(n386), .B1(n14780), .B2(n385), .ZN(n11172)
         );
  OAI22_X1 U4661 ( .A1(n9099), .A2(n386), .B1(n14740), .B2(n385), .ZN(n11173)
         );
  OAI22_X1 U4662 ( .A1(n9083), .A2(n386), .B1(n14700), .B2(n385), .ZN(n11174)
         );
  OAI22_X1 U4663 ( .A1(n9067), .A2(n386), .B1(n14660), .B2(n385), .ZN(n11175)
         );
  OAI22_X1 U4664 ( .A1(n9035), .A2(n388), .B1(n14900), .B2(n387), .ZN(n11177)
         );
  OAI22_X1 U4665 ( .A1(n9019), .A2(n388), .B1(n14860), .B2(n387), .ZN(n11178)
         );
  OAI22_X1 U4666 ( .A1(n9003), .A2(n388), .B1(n14820), .B2(n387), .ZN(n11179)
         );
  OAI22_X1 U4667 ( .A1(n8987), .A2(n388), .B1(n14780), .B2(n387), .ZN(n11180)
         );
  OAI22_X1 U4668 ( .A1(n8971), .A2(n388), .B1(n14740), .B2(n387), .ZN(n11181)
         );
  OAI22_X1 U4669 ( .A1(n8955), .A2(n388), .B1(n14700), .B2(n387), .ZN(n11182)
         );
  OAI22_X1 U4670 ( .A1(n8939), .A2(n388), .B1(n14660), .B2(n387), .ZN(n11183)
         );
  OAI22_X1 U4671 ( .A1(n8907), .A2(n390), .B1(n14900), .B2(n389), .ZN(n11185)
         );
  OAI22_X1 U4672 ( .A1(n8891), .A2(n390), .B1(n14860), .B2(n389), .ZN(n11186)
         );
  OAI22_X1 U4673 ( .A1(n8875), .A2(n390), .B1(n14820), .B2(n389), .ZN(n11187)
         );
  OAI22_X1 U4674 ( .A1(n8859), .A2(n390), .B1(n14780), .B2(n389), .ZN(n11188)
         );
  OAI22_X1 U4675 ( .A1(n8843), .A2(n390), .B1(n14740), .B2(n389), .ZN(n11189)
         );
  OAI22_X1 U4676 ( .A1(n8827), .A2(n390), .B1(n14700), .B2(n389), .ZN(n11190)
         );
  OAI22_X1 U4677 ( .A1(n8811), .A2(n390), .B1(n14660), .B2(n389), .ZN(n11191)
         );
  OAI22_X1 U4678 ( .A1(n8779), .A2(n392), .B1(n14900), .B2(n391), .ZN(n11193)
         );
  OAI22_X1 U4679 ( .A1(n8763), .A2(n392), .B1(n14860), .B2(n391), .ZN(n11194)
         );
  OAI22_X1 U4680 ( .A1(n8747), .A2(n392), .B1(n14820), .B2(n391), .ZN(n11195)
         );
  OAI22_X1 U4681 ( .A1(n8731), .A2(n392), .B1(n14780), .B2(n391), .ZN(n11196)
         );
  OAI22_X1 U4682 ( .A1(n8715), .A2(n392), .B1(n14740), .B2(n391), .ZN(n11197)
         );
  OAI22_X1 U4683 ( .A1(n8699), .A2(n392), .B1(n14700), .B2(n391), .ZN(n11198)
         );
  OAI22_X1 U4684 ( .A1(n8683), .A2(n392), .B1(n14660), .B2(n391), .ZN(n11199)
         );
  OAI22_X1 U4685 ( .A1(n8651), .A2(n394), .B1(n14900), .B2(n393), .ZN(n11201)
         );
  OAI22_X1 U4686 ( .A1(n8635), .A2(n394), .B1(n14860), .B2(n393), .ZN(n11202)
         );
  OAI22_X1 U4687 ( .A1(n8619), .A2(n394), .B1(n14820), .B2(n393), .ZN(n11203)
         );
  OAI22_X1 U4688 ( .A1(n8603), .A2(n394), .B1(n14780), .B2(n393), .ZN(n11204)
         );
  OAI22_X1 U4689 ( .A1(n8587), .A2(n394), .B1(n14740), .B2(n393), .ZN(n11205)
         );
  OAI22_X1 U4690 ( .A1(n8571), .A2(n394), .B1(n14700), .B2(n393), .ZN(n11206)
         );
  OAI22_X1 U4691 ( .A1(n8555), .A2(n394), .B1(n14660), .B2(n393), .ZN(n11207)
         );
  OAI22_X1 U4692 ( .A1(n8523), .A2(n396), .B1(n14900), .B2(n395), .ZN(n11209)
         );
  OAI22_X1 U4693 ( .A1(n8507), .A2(n396), .B1(n14860), .B2(n395), .ZN(n11210)
         );
  OAI22_X1 U4694 ( .A1(n8491), .A2(n396), .B1(n14820), .B2(n395), .ZN(n11211)
         );
  OAI22_X1 U4695 ( .A1(n8475), .A2(n396), .B1(n14780), .B2(n395), .ZN(n11212)
         );
  OAI22_X1 U4696 ( .A1(n8459), .A2(n396), .B1(n14740), .B2(n395), .ZN(n11213)
         );
  OAI22_X1 U4697 ( .A1(n8443), .A2(n396), .B1(n14700), .B2(n395), .ZN(n11214)
         );
  OAI22_X1 U4698 ( .A1(n8427), .A2(n396), .B1(n14660), .B2(n395), .ZN(n11215)
         );
  OAI22_X1 U4699 ( .A1(n8411), .A2(n397), .B1(n14968), .B2(n398), .ZN(n11216)
         );
  OAI22_X1 U4700 ( .A1(n8395), .A2(n397), .B1(n14900), .B2(n398), .ZN(n11217)
         );
  OAI22_X1 U4701 ( .A1(n8379), .A2(n397), .B1(n14860), .B2(n398), .ZN(n11218)
         );
  OAI22_X1 U4702 ( .A1(n8363), .A2(n397), .B1(n14820), .B2(n398), .ZN(n11219)
         );
  OAI22_X1 U4703 ( .A1(n8347), .A2(n397), .B1(n14780), .B2(n398), .ZN(n11220)
         );
  OAI22_X1 U4704 ( .A1(n8331), .A2(n397), .B1(n14740), .B2(n398), .ZN(n11221)
         );
  OAI22_X1 U4705 ( .A1(n8315), .A2(n397), .B1(n14700), .B2(n398), .ZN(n11222)
         );
  OAI22_X1 U4706 ( .A1(n8299), .A2(n397), .B1(n14660), .B2(n398), .ZN(n11223)
         );
  OAI22_X1 U4707 ( .A1(n8283), .A2(n399), .B1(n14968), .B2(n400), .ZN(n11224)
         );
  OAI22_X1 U4708 ( .A1(n8267), .A2(n399), .B1(n14900), .B2(n400), .ZN(n11225)
         );
  OAI22_X1 U4709 ( .A1(n8251), .A2(n399), .B1(n14860), .B2(n400), .ZN(n11226)
         );
  OAI22_X1 U4710 ( .A1(n8235), .A2(n399), .B1(n14820), .B2(n400), .ZN(n11227)
         );
  OAI22_X1 U4711 ( .A1(n8219), .A2(n399), .B1(n14780), .B2(n400), .ZN(n11228)
         );
  OAI22_X1 U4712 ( .A1(n8203), .A2(n399), .B1(n14740), .B2(n400), .ZN(n11229)
         );
  OAI22_X1 U4713 ( .A1(n8187), .A2(n399), .B1(n14700), .B2(n400), .ZN(n11230)
         );
  OAI22_X1 U4714 ( .A1(n8171), .A2(n399), .B1(n14660), .B2(n400), .ZN(n11231)
         );
  OAI22_X1 U4715 ( .A1(n8155), .A2(n401), .B1(n14968), .B2(n402), .ZN(n11232)
         );
  OAI22_X1 U4716 ( .A1(n8139), .A2(n401), .B1(n14901), .B2(n402), .ZN(n11233)
         );
  OAI22_X1 U4717 ( .A1(n8123), .A2(n401), .B1(n14861), .B2(n402), .ZN(n11234)
         );
  OAI22_X1 U4718 ( .A1(n8107), .A2(n401), .B1(n14821), .B2(n402), .ZN(n11235)
         );
  OAI22_X1 U4719 ( .A1(n8091), .A2(n401), .B1(n14781), .B2(n402), .ZN(n11236)
         );
  OAI22_X1 U4720 ( .A1(n8075), .A2(n401), .B1(n14741), .B2(n402), .ZN(n11237)
         );
  OAI22_X1 U4721 ( .A1(n8059), .A2(n401), .B1(n14701), .B2(n402), .ZN(n11238)
         );
  OAI22_X1 U4722 ( .A1(n8043), .A2(n401), .B1(n14661), .B2(n402), .ZN(n11239)
         );
  OAI22_X1 U4723 ( .A1(n8027), .A2(n403), .B1(n14968), .B2(n404), .ZN(n11240)
         );
  OAI22_X1 U4724 ( .A1(n8011), .A2(n403), .B1(n14901), .B2(n404), .ZN(n11241)
         );
  OAI22_X1 U4725 ( .A1(n7995), .A2(n403), .B1(n14861), .B2(n404), .ZN(n11242)
         );
  OAI22_X1 U4726 ( .A1(n7979), .A2(n403), .B1(n14821), .B2(n404), .ZN(n11243)
         );
  OAI22_X1 U4727 ( .A1(n7963), .A2(n403), .B1(n14781), .B2(n404), .ZN(n11244)
         );
  OAI22_X1 U4728 ( .A1(n7947), .A2(n403), .B1(n14741), .B2(n404), .ZN(n11245)
         );
  OAI22_X1 U4729 ( .A1(n7931), .A2(n403), .B1(n14701), .B2(n404), .ZN(n11246)
         );
  OAI22_X1 U4730 ( .A1(n7915), .A2(n403), .B1(n14661), .B2(n404), .ZN(n11247)
         );
  OAI22_X1 U4731 ( .A1(n7899), .A2(n405), .B1(n14968), .B2(n406), .ZN(n11248)
         );
  OAI22_X1 U4732 ( .A1(n7883), .A2(n405), .B1(n14901), .B2(n406), .ZN(n11249)
         );
  OAI22_X1 U4733 ( .A1(n7867), .A2(n405), .B1(n14861), .B2(n406), .ZN(n11250)
         );
  OAI22_X1 U4734 ( .A1(n7851), .A2(n405), .B1(n14821), .B2(n406), .ZN(n11251)
         );
  OAI22_X1 U4735 ( .A1(n7835), .A2(n405), .B1(n14781), .B2(n406), .ZN(n11252)
         );
  OAI22_X1 U4736 ( .A1(n7819), .A2(n405), .B1(n14741), .B2(n406), .ZN(n11253)
         );
  OAI22_X1 U4737 ( .A1(n7803), .A2(n405), .B1(n14701), .B2(n406), .ZN(n11254)
         );
  OAI22_X1 U4738 ( .A1(n7787), .A2(n405), .B1(n14661), .B2(n406), .ZN(n11255)
         );
  OAI22_X1 U4739 ( .A1(n7771), .A2(n407), .B1(n14967), .B2(n408), .ZN(n11256)
         );
  OAI22_X1 U4740 ( .A1(n7755), .A2(n407), .B1(n14901), .B2(n408), .ZN(n11257)
         );
  OAI22_X1 U4741 ( .A1(n7739), .A2(n407), .B1(n14861), .B2(n408), .ZN(n11258)
         );
  OAI22_X1 U4742 ( .A1(n7723), .A2(n407), .B1(n14821), .B2(n408), .ZN(n11259)
         );
  OAI22_X1 U4743 ( .A1(n7707), .A2(n407), .B1(n14781), .B2(n408), .ZN(n11260)
         );
  OAI22_X1 U4744 ( .A1(n7691), .A2(n407), .B1(n14741), .B2(n408), .ZN(n11261)
         );
  OAI22_X1 U4745 ( .A1(n7675), .A2(n407), .B1(n14701), .B2(n408), .ZN(n11262)
         );
  OAI22_X1 U4746 ( .A1(n7659), .A2(n407), .B1(n14661), .B2(n408), .ZN(n11263)
         );
  OAI22_X1 U4747 ( .A1(n9311), .A2(n449), .B1(n14966), .B2(n450), .ZN(n11416)
         );
  OAI22_X1 U4748 ( .A1(n9295), .A2(n449), .B1(n14902), .B2(n450), .ZN(n11417)
         );
  OAI22_X1 U4749 ( .A1(n9279), .A2(n449), .B1(n14862), .B2(n450), .ZN(n11418)
         );
  OAI22_X1 U4750 ( .A1(n9263), .A2(n449), .B1(n14822), .B2(n450), .ZN(n11419)
         );
  OAI22_X1 U4751 ( .A1(n9247), .A2(n449), .B1(n14782), .B2(n450), .ZN(n11420)
         );
  OAI22_X1 U4752 ( .A1(n9231), .A2(n449), .B1(n14742), .B2(n450), .ZN(n11421)
         );
  OAI22_X1 U4753 ( .A1(n9215), .A2(n449), .B1(n14702), .B2(n450), .ZN(n11422)
         );
  OAI22_X1 U4754 ( .A1(n9199), .A2(n449), .B1(n14662), .B2(n450), .ZN(n11423)
         );
  OAI22_X1 U4755 ( .A1(n9183), .A2(n451), .B1(n14966), .B2(n452), .ZN(n11424)
         );
  OAI22_X1 U4756 ( .A1(n9167), .A2(n451), .B1(n14902), .B2(n452), .ZN(n11425)
         );
  OAI22_X1 U4757 ( .A1(n9151), .A2(n451), .B1(n14862), .B2(n452), .ZN(n11426)
         );
  OAI22_X1 U4758 ( .A1(n9135), .A2(n451), .B1(n14822), .B2(n452), .ZN(n11427)
         );
  OAI22_X1 U4759 ( .A1(n9119), .A2(n451), .B1(n14782), .B2(n452), .ZN(n11428)
         );
  OAI22_X1 U4760 ( .A1(n9103), .A2(n451), .B1(n14742), .B2(n452), .ZN(n11429)
         );
  OAI22_X1 U4761 ( .A1(n9087), .A2(n451), .B1(n14702), .B2(n452), .ZN(n11430)
         );
  OAI22_X1 U4762 ( .A1(n9071), .A2(n451), .B1(n14662), .B2(n452), .ZN(n11431)
         );
  OAI22_X1 U4763 ( .A1(n9055), .A2(n453), .B1(n14966), .B2(n454), .ZN(n11432)
         );
  OAI22_X1 U4764 ( .A1(n9039), .A2(n453), .B1(n14902), .B2(n454), .ZN(n11433)
         );
  OAI22_X1 U4765 ( .A1(n9023), .A2(n453), .B1(n14862), .B2(n454), .ZN(n11434)
         );
  OAI22_X1 U4766 ( .A1(n9007), .A2(n453), .B1(n14822), .B2(n454), .ZN(n11435)
         );
  OAI22_X1 U4767 ( .A1(n8991), .A2(n453), .B1(n14782), .B2(n454), .ZN(n11436)
         );
  OAI22_X1 U4768 ( .A1(n8975), .A2(n453), .B1(n14742), .B2(n454), .ZN(n11437)
         );
  OAI22_X1 U4769 ( .A1(n8959), .A2(n453), .B1(n14702), .B2(n454), .ZN(n11438)
         );
  OAI22_X1 U4770 ( .A1(n8943), .A2(n453), .B1(n14662), .B2(n454), .ZN(n11439)
         );
  OAI22_X1 U4771 ( .A1(n8927), .A2(n455), .B1(n14966), .B2(n456), .ZN(n11440)
         );
  OAI22_X1 U4772 ( .A1(n8911), .A2(n455), .B1(n14903), .B2(n456), .ZN(n11441)
         );
  OAI22_X1 U4773 ( .A1(n8895), .A2(n455), .B1(n14863), .B2(n456), .ZN(n11442)
         );
  OAI22_X1 U4774 ( .A1(n8879), .A2(n455), .B1(n14823), .B2(n456), .ZN(n11443)
         );
  OAI22_X1 U4775 ( .A1(n8863), .A2(n455), .B1(n14783), .B2(n456), .ZN(n11444)
         );
  OAI22_X1 U4776 ( .A1(n8847), .A2(n455), .B1(n14743), .B2(n456), .ZN(n11445)
         );
  OAI22_X1 U4777 ( .A1(n8831), .A2(n455), .B1(n14703), .B2(n456), .ZN(n11446)
         );
  OAI22_X1 U4778 ( .A1(n8815), .A2(n455), .B1(n14663), .B2(n456), .ZN(n11447)
         );
  OAI22_X1 U4779 ( .A1(n8799), .A2(n457), .B1(n14966), .B2(n458), .ZN(n11448)
         );
  OAI22_X1 U4780 ( .A1(n8783), .A2(n457), .B1(n14903), .B2(n458), .ZN(n11449)
         );
  OAI22_X1 U4781 ( .A1(n8767), .A2(n457), .B1(n14863), .B2(n458), .ZN(n11450)
         );
  OAI22_X1 U4782 ( .A1(n8751), .A2(n457), .B1(n14823), .B2(n458), .ZN(n11451)
         );
  OAI22_X1 U4783 ( .A1(n8735), .A2(n457), .B1(n14783), .B2(n458), .ZN(n11452)
         );
  OAI22_X1 U4784 ( .A1(n8719), .A2(n457), .B1(n14743), .B2(n458), .ZN(n11453)
         );
  OAI22_X1 U4785 ( .A1(n8703), .A2(n457), .B1(n14703), .B2(n458), .ZN(n11454)
         );
  OAI22_X1 U4786 ( .A1(n8687), .A2(n457), .B1(n14663), .B2(n458), .ZN(n11455)
         );
  OAI22_X1 U4787 ( .A1(n8671), .A2(n459), .B1(n14966), .B2(n460), .ZN(n11456)
         );
  OAI22_X1 U4788 ( .A1(n8655), .A2(n459), .B1(n14903), .B2(n460), .ZN(n11457)
         );
  OAI22_X1 U4789 ( .A1(n8639), .A2(n459), .B1(n14863), .B2(n460), .ZN(n11458)
         );
  OAI22_X1 U4790 ( .A1(n8623), .A2(n459), .B1(n14823), .B2(n460), .ZN(n11459)
         );
  OAI22_X1 U4791 ( .A1(n8607), .A2(n459), .B1(n14783), .B2(n460), .ZN(n11460)
         );
  OAI22_X1 U4792 ( .A1(n8591), .A2(n459), .B1(n14743), .B2(n460), .ZN(n11461)
         );
  OAI22_X1 U4793 ( .A1(n8575), .A2(n459), .B1(n14703), .B2(n460), .ZN(n11462)
         );
  OAI22_X1 U4794 ( .A1(n8559), .A2(n459), .B1(n14663), .B2(n460), .ZN(n11463)
         );
  OAI22_X1 U4795 ( .A1(n8543), .A2(n461), .B1(n14965), .B2(n462), .ZN(n11464)
         );
  OAI22_X1 U4796 ( .A1(n8527), .A2(n461), .B1(n14903), .B2(n462), .ZN(n11465)
         );
  OAI22_X1 U4797 ( .A1(n8511), .A2(n461), .B1(n14863), .B2(n462), .ZN(n11466)
         );
  OAI22_X1 U4798 ( .A1(n8495), .A2(n461), .B1(n14823), .B2(n462), .ZN(n11467)
         );
  OAI22_X1 U4799 ( .A1(n8479), .A2(n461), .B1(n14783), .B2(n462), .ZN(n11468)
         );
  OAI22_X1 U4800 ( .A1(n8463), .A2(n461), .B1(n14743), .B2(n462), .ZN(n11469)
         );
  OAI22_X1 U4801 ( .A1(n8447), .A2(n461), .B1(n14703), .B2(n462), .ZN(n11470)
         );
  OAI22_X1 U4802 ( .A1(n8431), .A2(n461), .B1(n14663), .B2(n462), .ZN(n11471)
         );
  OAI22_X1 U4803 ( .A1(n8415), .A2(n463), .B1(n14965), .B2(n464), .ZN(n11472)
         );
  OAI22_X1 U4804 ( .A1(n8399), .A2(n463), .B1(n14903), .B2(n464), .ZN(n11473)
         );
  OAI22_X1 U4805 ( .A1(n8383), .A2(n463), .B1(n14863), .B2(n464), .ZN(n11474)
         );
  OAI22_X1 U4806 ( .A1(n8367), .A2(n463), .B1(n14823), .B2(n464), .ZN(n11475)
         );
  OAI22_X1 U4807 ( .A1(n8351), .A2(n463), .B1(n14783), .B2(n464), .ZN(n11476)
         );
  OAI22_X1 U4808 ( .A1(n8335), .A2(n463), .B1(n14743), .B2(n464), .ZN(n11477)
         );
  OAI22_X1 U4809 ( .A1(n8319), .A2(n463), .B1(n14703), .B2(n464), .ZN(n11478)
         );
  OAI22_X1 U4810 ( .A1(n8303), .A2(n463), .B1(n14663), .B2(n464), .ZN(n11479)
         );
  OAI22_X1 U4811 ( .A1(n8287), .A2(n465), .B1(n14965), .B2(n466), .ZN(n11480)
         );
  OAI22_X1 U4812 ( .A1(n8271), .A2(n465), .B1(n14903), .B2(n466), .ZN(n11481)
         );
  OAI22_X1 U4813 ( .A1(n8255), .A2(n465), .B1(n14863), .B2(n466), .ZN(n11482)
         );
  OAI22_X1 U4814 ( .A1(n8239), .A2(n465), .B1(n14823), .B2(n466), .ZN(n11483)
         );
  OAI22_X1 U4815 ( .A1(n8223), .A2(n465), .B1(n14783), .B2(n466), .ZN(n11484)
         );
  OAI22_X1 U4816 ( .A1(n8207), .A2(n465), .B1(n14743), .B2(n466), .ZN(n11485)
         );
  OAI22_X1 U4817 ( .A1(n8191), .A2(n465), .B1(n14703), .B2(n466), .ZN(n11486)
         );
  OAI22_X1 U4818 ( .A1(n8175), .A2(n465), .B1(n14663), .B2(n466), .ZN(n11487)
         );
  OAI22_X1 U4819 ( .A1(n8159), .A2(n467), .B1(n14965), .B2(n468), .ZN(n11488)
         );
  OAI22_X1 U4820 ( .A1(n8143), .A2(n467), .B1(n14903), .B2(n468), .ZN(n11489)
         );
  OAI22_X1 U4821 ( .A1(n8127), .A2(n467), .B1(n14863), .B2(n468), .ZN(n11490)
         );
  OAI22_X1 U4822 ( .A1(n8111), .A2(n467), .B1(n14823), .B2(n468), .ZN(n11491)
         );
  OAI22_X1 U4823 ( .A1(n8095), .A2(n467), .B1(n14783), .B2(n468), .ZN(n11492)
         );
  OAI22_X1 U4824 ( .A1(n8079), .A2(n467), .B1(n14743), .B2(n468), .ZN(n11493)
         );
  OAI22_X1 U4825 ( .A1(n8063), .A2(n467), .B1(n14703), .B2(n468), .ZN(n11494)
         );
  OAI22_X1 U4826 ( .A1(n8047), .A2(n467), .B1(n14663), .B2(n468), .ZN(n11495)
         );
  OAI22_X1 U4827 ( .A1(n8031), .A2(n469), .B1(n14965), .B2(n470), .ZN(n11496)
         );
  OAI22_X1 U4828 ( .A1(n8015), .A2(n469), .B1(n14903), .B2(n470), .ZN(n11497)
         );
  OAI22_X1 U4829 ( .A1(n7999), .A2(n469), .B1(n14863), .B2(n470), .ZN(n11498)
         );
  OAI22_X1 U4830 ( .A1(n7983), .A2(n469), .B1(n14823), .B2(n470), .ZN(n11499)
         );
  OAI22_X1 U4831 ( .A1(n7967), .A2(n469), .B1(n14783), .B2(n470), .ZN(n11500)
         );
  OAI22_X1 U4832 ( .A1(n7951), .A2(n469), .B1(n14743), .B2(n470), .ZN(n11501)
         );
  OAI22_X1 U4833 ( .A1(n7935), .A2(n469), .B1(n14703), .B2(n470), .ZN(n11502)
         );
  OAI22_X1 U4834 ( .A1(n7919), .A2(n469), .B1(n14663), .B2(n470), .ZN(n11503)
         );
  OAI22_X1 U4835 ( .A1(n7903), .A2(n471), .B1(n14965), .B2(n472), .ZN(n11504)
         );
  OAI22_X1 U4836 ( .A1(n7887), .A2(n471), .B1(n14903), .B2(n472), .ZN(n11505)
         );
  OAI22_X1 U4837 ( .A1(n7871), .A2(n471), .B1(n14863), .B2(n472), .ZN(n11506)
         );
  OAI22_X1 U4838 ( .A1(n7855), .A2(n471), .B1(n14823), .B2(n472), .ZN(n11507)
         );
  OAI22_X1 U4839 ( .A1(n7839), .A2(n471), .B1(n14783), .B2(n472), .ZN(n11508)
         );
  OAI22_X1 U4840 ( .A1(n7823), .A2(n471), .B1(n14743), .B2(n472), .ZN(n11509)
         );
  OAI22_X1 U4841 ( .A1(n7807), .A2(n471), .B1(n14703), .B2(n472), .ZN(n11510)
         );
  OAI22_X1 U4842 ( .A1(n7791), .A2(n471), .B1(n14663), .B2(n472), .ZN(n11511)
         );
  OAI22_X1 U4843 ( .A1(n7775), .A2(n473), .B1(n14965), .B2(n474), .ZN(n11512)
         );
  OAI22_X1 U4844 ( .A1(n7759), .A2(n473), .B1(n14903), .B2(n474), .ZN(n11513)
         );
  OAI22_X1 U4845 ( .A1(n7743), .A2(n473), .B1(n14863), .B2(n474), .ZN(n11514)
         );
  OAI22_X1 U4846 ( .A1(n7727), .A2(n473), .B1(n14823), .B2(n474), .ZN(n11515)
         );
  OAI22_X1 U4847 ( .A1(n7711), .A2(n473), .B1(n14783), .B2(n474), .ZN(n11516)
         );
  OAI22_X1 U4848 ( .A1(n7695), .A2(n473), .B1(n14743), .B2(n474), .ZN(n11517)
         );
  OAI22_X1 U4849 ( .A1(n7679), .A2(n473), .B1(n14703), .B2(n474), .ZN(n11518)
         );
  OAI22_X1 U4850 ( .A1(n7663), .A2(n473), .B1(n14663), .B2(n474), .ZN(n11519)
         );
  OAI22_X1 U4851 ( .A1(n10072), .A2(n632), .B1(n14964), .B2(n633), .ZN(n12136)
         );
  OAI22_X1 U4852 ( .A1(n10056), .A2(n632), .B1(n14909), .B2(n633), .ZN(n12137)
         );
  OAI22_X1 U4853 ( .A1(n10040), .A2(n632), .B1(n14869), .B2(n633), .ZN(n12138)
         );
  OAI22_X1 U4854 ( .A1(n10024), .A2(n632), .B1(n14829), .B2(n633), .ZN(n12139)
         );
  OAI22_X1 U4855 ( .A1(n10008), .A2(n632), .B1(n14789), .B2(n633), .ZN(n12140)
         );
  OAI22_X1 U4856 ( .A1(n9992), .A2(n632), .B1(n14749), .B2(n633), .ZN(n12141)
         );
  OAI22_X1 U4857 ( .A1(n9976), .A2(n632), .B1(n14709), .B2(n633), .ZN(n12142)
         );
  OAI22_X1 U4858 ( .A1(n9960), .A2(n632), .B1(n14669), .B2(n633), .ZN(n12143)
         );
  OAI22_X1 U4859 ( .A1(n9944), .A2(n635), .B1(n14939), .B2(n636), .ZN(n12144)
         );
  OAI22_X1 U4860 ( .A1(n9928), .A2(n635), .B1(n14909), .B2(n636), .ZN(n12145)
         );
  OAI22_X1 U4861 ( .A1(n9912), .A2(n635), .B1(n14869), .B2(n636), .ZN(n12146)
         );
  OAI22_X1 U4862 ( .A1(n9896), .A2(n635), .B1(n14829), .B2(n636), .ZN(n12147)
         );
  OAI22_X1 U4863 ( .A1(n9880), .A2(n635), .B1(n14789), .B2(n636), .ZN(n12148)
         );
  OAI22_X1 U4864 ( .A1(n9864), .A2(n635), .B1(n14749), .B2(n636), .ZN(n12149)
         );
  OAI22_X1 U4865 ( .A1(n9848), .A2(n635), .B1(n14709), .B2(n636), .ZN(n12150)
         );
  OAI22_X1 U4866 ( .A1(n9832), .A2(n635), .B1(n14669), .B2(n636), .ZN(n12151)
         );
  OAI22_X1 U4867 ( .A1(n9816), .A2(n637), .B1(n14939), .B2(n638), .ZN(n12152)
         );
  OAI22_X1 U4868 ( .A1(n9800), .A2(n637), .B1(n14909), .B2(n638), .ZN(n12153)
         );
  OAI22_X1 U4869 ( .A1(n9784), .A2(n637), .B1(n14869), .B2(n638), .ZN(n12154)
         );
  OAI22_X1 U4870 ( .A1(n9768), .A2(n637), .B1(n14829), .B2(n638), .ZN(n12155)
         );
  OAI22_X1 U4871 ( .A1(n9752), .A2(n637), .B1(n14789), .B2(n638), .ZN(n12156)
         );
  OAI22_X1 U4872 ( .A1(n9736), .A2(n637), .B1(n14749), .B2(n638), .ZN(n12157)
         );
  OAI22_X1 U4873 ( .A1(n9720), .A2(n637), .B1(n14709), .B2(n638), .ZN(n12158)
         );
  OAI22_X1 U4874 ( .A1(n9704), .A2(n637), .B1(n14669), .B2(n638), .ZN(n12159)
         );
  OAI22_X1 U4875 ( .A1(n9688), .A2(n639), .B1(n14939), .B2(n640), .ZN(n12160)
         );
  OAI22_X1 U4876 ( .A1(n9672), .A2(n639), .B1(n14909), .B2(n640), .ZN(n12161)
         );
  OAI22_X1 U4877 ( .A1(n9656), .A2(n639), .B1(n14869), .B2(n640), .ZN(n12162)
         );
  OAI22_X1 U4878 ( .A1(n9640), .A2(n639), .B1(n14829), .B2(n640), .ZN(n12163)
         );
  OAI22_X1 U4879 ( .A1(n9624), .A2(n639), .B1(n14789), .B2(n640), .ZN(n12164)
         );
  OAI22_X1 U4880 ( .A1(n9608), .A2(n639), .B1(n14749), .B2(n640), .ZN(n12165)
         );
  OAI22_X1 U4881 ( .A1(n9592), .A2(n639), .B1(n14709), .B2(n640), .ZN(n12166)
         );
  OAI22_X1 U4882 ( .A1(n9576), .A2(n639), .B1(n14669), .B2(n640), .ZN(n12167)
         );
  OAI22_X1 U4883 ( .A1(n9560), .A2(n641), .B1(n14939), .B2(n642), .ZN(n12168)
         );
  OAI22_X1 U4884 ( .A1(n9544), .A2(n641), .B1(n14910), .B2(n642), .ZN(n12169)
         );
  OAI22_X1 U4885 ( .A1(n9528), .A2(n641), .B1(n14870), .B2(n642), .ZN(n12170)
         );
  OAI22_X1 U4886 ( .A1(n9512), .A2(n641), .B1(n14830), .B2(n642), .ZN(n12171)
         );
  OAI22_X1 U4887 ( .A1(n9496), .A2(n641), .B1(n14790), .B2(n642), .ZN(n12172)
         );
  OAI22_X1 U4888 ( .A1(n9480), .A2(n641), .B1(n14750), .B2(n642), .ZN(n12173)
         );
  OAI22_X1 U4889 ( .A1(n9464), .A2(n641), .B1(n14710), .B2(n642), .ZN(n12174)
         );
  OAI22_X1 U4890 ( .A1(n9448), .A2(n641), .B1(n14670), .B2(n642), .ZN(n12175)
         );
  OAI22_X1 U4891 ( .A1(n9432), .A2(n643), .B1(n14939), .B2(n644), .ZN(n12176)
         );
  OAI22_X1 U4892 ( .A1(n9416), .A2(n643), .B1(n14910), .B2(n644), .ZN(n12177)
         );
  OAI22_X1 U4893 ( .A1(n9400), .A2(n643), .B1(n14870), .B2(n644), .ZN(n12178)
         );
  OAI22_X1 U4894 ( .A1(n9384), .A2(n643), .B1(n14830), .B2(n644), .ZN(n12179)
         );
  OAI22_X1 U4895 ( .A1(n9368), .A2(n643), .B1(n14790), .B2(n644), .ZN(n12180)
         );
  OAI22_X1 U4896 ( .A1(n9352), .A2(n643), .B1(n14750), .B2(n644), .ZN(n12181)
         );
  OAI22_X1 U4897 ( .A1(n9336), .A2(n643), .B1(n14710), .B2(n644), .ZN(n12182)
         );
  OAI22_X1 U4898 ( .A1(n9320), .A2(n643), .B1(n14670), .B2(n644), .ZN(n12183)
         );
  OAI22_X1 U4899 ( .A1(n9304), .A2(n645), .B1(n14939), .B2(n646), .ZN(n12184)
         );
  OAI22_X1 U4900 ( .A1(n9288), .A2(n645), .B1(n14910), .B2(n646), .ZN(n12185)
         );
  OAI22_X1 U4901 ( .A1(n9272), .A2(n645), .B1(n14870), .B2(n646), .ZN(n12186)
         );
  OAI22_X1 U4902 ( .A1(n9256), .A2(n645), .B1(n14830), .B2(n646), .ZN(n12187)
         );
  OAI22_X1 U4903 ( .A1(n9240), .A2(n645), .B1(n14790), .B2(n646), .ZN(n12188)
         );
  OAI22_X1 U4904 ( .A1(n9224), .A2(n645), .B1(n14750), .B2(n646), .ZN(n12189)
         );
  OAI22_X1 U4905 ( .A1(n9208), .A2(n645), .B1(n14710), .B2(n646), .ZN(n12190)
         );
  OAI22_X1 U4906 ( .A1(n9192), .A2(n645), .B1(n14670), .B2(n646), .ZN(n12191)
         );
  OAI22_X1 U4907 ( .A1(n9176), .A2(n647), .B1(n14939), .B2(n648), .ZN(n12192)
         );
  OAI22_X1 U4908 ( .A1(n9160), .A2(n647), .B1(n14910), .B2(n648), .ZN(n12193)
         );
  OAI22_X1 U4909 ( .A1(n9144), .A2(n647), .B1(n14870), .B2(n648), .ZN(n12194)
         );
  OAI22_X1 U4910 ( .A1(n9128), .A2(n647), .B1(n14830), .B2(n648), .ZN(n12195)
         );
  OAI22_X1 U4911 ( .A1(n9112), .A2(n647), .B1(n14790), .B2(n648), .ZN(n12196)
         );
  OAI22_X1 U4912 ( .A1(n9096), .A2(n647), .B1(n14750), .B2(n648), .ZN(n12197)
         );
  OAI22_X1 U4913 ( .A1(n9080), .A2(n647), .B1(n14710), .B2(n648), .ZN(n12198)
         );
  OAI22_X1 U4914 ( .A1(n9064), .A2(n647), .B1(n14670), .B2(n648), .ZN(n12199)
         );
  OAI22_X1 U4915 ( .A1(n9048), .A2(n649), .B1(n14939), .B2(n650), .ZN(n12200)
         );
  OAI22_X1 U4916 ( .A1(n9032), .A2(n649), .B1(n14910), .B2(n650), .ZN(n12201)
         );
  OAI22_X1 U4917 ( .A1(n9016), .A2(n649), .B1(n14870), .B2(n650), .ZN(n12202)
         );
  OAI22_X1 U4918 ( .A1(n9000), .A2(n649), .B1(n14830), .B2(n650), .ZN(n12203)
         );
  OAI22_X1 U4919 ( .A1(n8984), .A2(n649), .B1(n14790), .B2(n650), .ZN(n12204)
         );
  OAI22_X1 U4920 ( .A1(n8968), .A2(n649), .B1(n14750), .B2(n650), .ZN(n12205)
         );
  OAI22_X1 U4921 ( .A1(n8952), .A2(n649), .B1(n14710), .B2(n650), .ZN(n12206)
         );
  OAI22_X1 U4922 ( .A1(n8936), .A2(n649), .B1(n14670), .B2(n650), .ZN(n12207)
         );
  OAI22_X1 U4923 ( .A1(n8920), .A2(n651), .B1(n14939), .B2(n652), .ZN(n12208)
         );
  OAI22_X1 U4924 ( .A1(n8904), .A2(n651), .B1(n14910), .B2(n652), .ZN(n12209)
         );
  OAI22_X1 U4925 ( .A1(n8888), .A2(n651), .B1(n14870), .B2(n652), .ZN(n12210)
         );
  OAI22_X1 U4926 ( .A1(n8872), .A2(n651), .B1(n14830), .B2(n652), .ZN(n12211)
         );
  OAI22_X1 U4927 ( .A1(n8856), .A2(n651), .B1(n14790), .B2(n652), .ZN(n12212)
         );
  OAI22_X1 U4928 ( .A1(n8840), .A2(n651), .B1(n14750), .B2(n652), .ZN(n12213)
         );
  OAI22_X1 U4929 ( .A1(n8824), .A2(n651), .B1(n14710), .B2(n652), .ZN(n12214)
         );
  OAI22_X1 U4930 ( .A1(n8808), .A2(n651), .B1(n14670), .B2(n652), .ZN(n12215)
         );
  OAI22_X1 U4931 ( .A1(n8792), .A2(n653), .B1(n14939), .B2(n654), .ZN(n12216)
         );
  OAI22_X1 U4932 ( .A1(n8776), .A2(n653), .B1(n14910), .B2(n654), .ZN(n12217)
         );
  OAI22_X1 U4933 ( .A1(n8760), .A2(n653), .B1(n14870), .B2(n654), .ZN(n12218)
         );
  OAI22_X1 U4934 ( .A1(n8744), .A2(n653), .B1(n14830), .B2(n654), .ZN(n12219)
         );
  OAI22_X1 U4935 ( .A1(n8728), .A2(n653), .B1(n14790), .B2(n654), .ZN(n12220)
         );
  OAI22_X1 U4936 ( .A1(n8712), .A2(n653), .B1(n14750), .B2(n654), .ZN(n12221)
         );
  OAI22_X1 U4937 ( .A1(n8696), .A2(n653), .B1(n14710), .B2(n654), .ZN(n12222)
         );
  OAI22_X1 U4938 ( .A1(n8680), .A2(n653), .B1(n14670), .B2(n654), .ZN(n12223)
         );
  OAI22_X1 U4939 ( .A1(n8664), .A2(n655), .B1(n14939), .B2(n656), .ZN(n12224)
         );
  OAI22_X1 U4940 ( .A1(n8648), .A2(n655), .B1(n14910), .B2(n656), .ZN(n12225)
         );
  OAI22_X1 U4941 ( .A1(n8632), .A2(n655), .B1(n14870), .B2(n656), .ZN(n12226)
         );
  OAI22_X1 U4942 ( .A1(n8616), .A2(n655), .B1(n14830), .B2(n656), .ZN(n12227)
         );
  OAI22_X1 U4943 ( .A1(n8600), .A2(n655), .B1(n14790), .B2(n656), .ZN(n12228)
         );
  OAI22_X1 U4944 ( .A1(n8584), .A2(n655), .B1(n14750), .B2(n656), .ZN(n12229)
         );
  OAI22_X1 U4945 ( .A1(n8568), .A2(n655), .B1(n14710), .B2(n656), .ZN(n12230)
         );
  OAI22_X1 U4946 ( .A1(n8552), .A2(n655), .B1(n14670), .B2(n656), .ZN(n12231)
         );
  OAI22_X1 U4947 ( .A1(n8536), .A2(n657), .B1(n14939), .B2(n658), .ZN(n12232)
         );
  OAI22_X1 U4948 ( .A1(n8520), .A2(n657), .B1(n14910), .B2(n658), .ZN(n12233)
         );
  OAI22_X1 U4949 ( .A1(n8504), .A2(n657), .B1(n14870), .B2(n658), .ZN(n12234)
         );
  OAI22_X1 U4950 ( .A1(n8488), .A2(n657), .B1(n14830), .B2(n658), .ZN(n12235)
         );
  OAI22_X1 U4951 ( .A1(n8472), .A2(n657), .B1(n14790), .B2(n658), .ZN(n12236)
         );
  OAI22_X1 U4952 ( .A1(n8456), .A2(n657), .B1(n14750), .B2(n658), .ZN(n12237)
         );
  OAI22_X1 U4953 ( .A1(n8440), .A2(n657), .B1(n14710), .B2(n658), .ZN(n12238)
         );
  OAI22_X1 U4954 ( .A1(n8424), .A2(n657), .B1(n14670), .B2(n658), .ZN(n12239)
         );
  OAI22_X1 U4955 ( .A1(n8408), .A2(n659), .B1(n14938), .B2(n660), .ZN(n12240)
         );
  OAI22_X1 U4956 ( .A1(n8392), .A2(n659), .B1(n14910), .B2(n660), .ZN(n12241)
         );
  OAI22_X1 U4957 ( .A1(n8376), .A2(n659), .B1(n14870), .B2(n660), .ZN(n12242)
         );
  OAI22_X1 U4958 ( .A1(n8360), .A2(n659), .B1(n14830), .B2(n660), .ZN(n12243)
         );
  OAI22_X1 U4959 ( .A1(n8344), .A2(n659), .B1(n14790), .B2(n660), .ZN(n12244)
         );
  OAI22_X1 U4960 ( .A1(n8328), .A2(n659), .B1(n14750), .B2(n660), .ZN(n12245)
         );
  OAI22_X1 U4961 ( .A1(n8312), .A2(n659), .B1(n14710), .B2(n660), .ZN(n12246)
         );
  OAI22_X1 U4962 ( .A1(n8296), .A2(n659), .B1(n14670), .B2(n660), .ZN(n12247)
         );
  OAI22_X1 U4963 ( .A1(n8280), .A2(n661), .B1(n14938), .B2(n662), .ZN(n12248)
         );
  OAI22_X1 U4964 ( .A1(n8264), .A2(n661), .B1(n14910), .B2(n662), .ZN(n12249)
         );
  OAI22_X1 U4965 ( .A1(n8248), .A2(n661), .B1(n14870), .B2(n662), .ZN(n12250)
         );
  OAI22_X1 U4966 ( .A1(n8232), .A2(n661), .B1(n14830), .B2(n662), .ZN(n12251)
         );
  OAI22_X1 U4967 ( .A1(n8216), .A2(n661), .B1(n14790), .B2(n662), .ZN(n12252)
         );
  OAI22_X1 U4968 ( .A1(n8200), .A2(n661), .B1(n14750), .B2(n662), .ZN(n12253)
         );
  OAI22_X1 U4969 ( .A1(n8184), .A2(n661), .B1(n14710), .B2(n662), .ZN(n12254)
         );
  OAI22_X1 U4970 ( .A1(n8168), .A2(n661), .B1(n14670), .B2(n662), .ZN(n12255)
         );
  OAI22_X1 U4971 ( .A1(n8152), .A2(n663), .B1(n14938), .B2(n664), .ZN(n12256)
         );
  OAI22_X1 U4972 ( .A1(n8136), .A2(n663), .B1(n14910), .B2(n664), .ZN(n12257)
         );
  OAI22_X1 U4973 ( .A1(n8120), .A2(n663), .B1(n14870), .B2(n664), .ZN(n12258)
         );
  OAI22_X1 U4974 ( .A1(n8104), .A2(n663), .B1(n14830), .B2(n664), .ZN(n12259)
         );
  OAI22_X1 U4975 ( .A1(n8088), .A2(n663), .B1(n14790), .B2(n664), .ZN(n12260)
         );
  OAI22_X1 U4976 ( .A1(n8072), .A2(n663), .B1(n14750), .B2(n664), .ZN(n12261)
         );
  OAI22_X1 U4977 ( .A1(n8056), .A2(n663), .B1(n14710), .B2(n664), .ZN(n12262)
         );
  OAI22_X1 U4978 ( .A1(n8040), .A2(n663), .B1(n14670), .B2(n664), .ZN(n12263)
         );
  OAI22_X1 U4979 ( .A1(n8024), .A2(n665), .B1(n14938), .B2(n666), .ZN(n12264)
         );
  OAI22_X1 U4980 ( .A1(n8008), .A2(n665), .B1(n14910), .B2(n666), .ZN(n12265)
         );
  OAI22_X1 U4981 ( .A1(n7992), .A2(n665), .B1(n14870), .B2(n666), .ZN(n12266)
         );
  OAI22_X1 U4982 ( .A1(n7976), .A2(n665), .B1(n14830), .B2(n666), .ZN(n12267)
         );
  OAI22_X1 U4983 ( .A1(n7960), .A2(n665), .B1(n14790), .B2(n666), .ZN(n12268)
         );
  OAI22_X1 U4984 ( .A1(n7944), .A2(n665), .B1(n14750), .B2(n666), .ZN(n12269)
         );
  OAI22_X1 U4985 ( .A1(n7928), .A2(n665), .B1(n14710), .B2(n666), .ZN(n12270)
         );
  OAI22_X1 U4986 ( .A1(n7912), .A2(n665), .B1(n14670), .B2(n666), .ZN(n12271)
         );
  OAI22_X1 U4987 ( .A1(n7896), .A2(n667), .B1(n14938), .B2(n668), .ZN(n12272)
         );
  OAI22_X1 U4988 ( .A1(n7880), .A2(n667), .B1(n14911), .B2(n668), .ZN(n12273)
         );
  OAI22_X1 U4989 ( .A1(n7864), .A2(n667), .B1(n14871), .B2(n668), .ZN(n12274)
         );
  OAI22_X1 U4990 ( .A1(n7848), .A2(n667), .B1(n14831), .B2(n668), .ZN(n12275)
         );
  OAI22_X1 U4991 ( .A1(n7832), .A2(n667), .B1(n14791), .B2(n668), .ZN(n12276)
         );
  OAI22_X1 U4992 ( .A1(n7816), .A2(n667), .B1(n14751), .B2(n668), .ZN(n12277)
         );
  OAI22_X1 U4993 ( .A1(n7800), .A2(n667), .B1(n14711), .B2(n668), .ZN(n12278)
         );
  OAI22_X1 U4994 ( .A1(n7784), .A2(n667), .B1(n14671), .B2(n668), .ZN(n12279)
         );
  OAI22_X1 U4995 ( .A1(n7768), .A2(n669), .B1(n14938), .B2(n670), .ZN(n12280)
         );
  OAI22_X1 U4996 ( .A1(n7752), .A2(n669), .B1(n14911), .B2(n670), .ZN(n12281)
         );
  OAI22_X1 U4997 ( .A1(n7736), .A2(n669), .B1(n14871), .B2(n670), .ZN(n12282)
         );
  OAI22_X1 U4998 ( .A1(n7720), .A2(n669), .B1(n14831), .B2(n670), .ZN(n12283)
         );
  OAI22_X1 U4999 ( .A1(n7704), .A2(n669), .B1(n14791), .B2(n670), .ZN(n12284)
         );
  OAI22_X1 U5000 ( .A1(n7688), .A2(n669), .B1(n14751), .B2(n670), .ZN(n12285)
         );
  OAI22_X1 U5001 ( .A1(n7672), .A2(n669), .B1(n14711), .B2(n670), .ZN(n12286)
         );
  OAI22_X1 U5002 ( .A1(n7656), .A2(n669), .B1(n14671), .B2(n670), .ZN(n12287)
         );
  OAI22_X1 U5003 ( .A1(n7640), .A2(n671), .B1(n14938), .B2(n672), .ZN(n12288)
         );
  OAI22_X1 U5004 ( .A1(n7624), .A2(n671), .B1(n14911), .B2(n672), .ZN(n12289)
         );
  OAI22_X1 U5005 ( .A1(n7608), .A2(n671), .B1(n14871), .B2(n672), .ZN(n12290)
         );
  OAI22_X1 U5006 ( .A1(n7592), .A2(n671), .B1(n14831), .B2(n672), .ZN(n12291)
         );
  OAI22_X1 U5007 ( .A1(n7576), .A2(n671), .B1(n14791), .B2(n672), .ZN(n12292)
         );
  OAI22_X1 U5008 ( .A1(n7560), .A2(n671), .B1(n14751), .B2(n672), .ZN(n12293)
         );
  OAI22_X1 U5009 ( .A1(n7544), .A2(n671), .B1(n14711), .B2(n672), .ZN(n12294)
         );
  OAI22_X1 U5010 ( .A1(n7528), .A2(n671), .B1(n14671), .B2(n672), .ZN(n12295)
         );
  OAI22_X1 U5011 ( .A1(n7512), .A2(n673), .B1(n14938), .B2(n674), .ZN(n12296)
         );
  OAI22_X1 U5012 ( .A1(n7496), .A2(n673), .B1(n14911), .B2(n674), .ZN(n12297)
         );
  OAI22_X1 U5013 ( .A1(n7480), .A2(n673), .B1(n14871), .B2(n674), .ZN(n12298)
         );
  OAI22_X1 U5014 ( .A1(n7464), .A2(n673), .B1(n14831), .B2(n674), .ZN(n12299)
         );
  OAI22_X1 U5015 ( .A1(n7448), .A2(n673), .B1(n14791), .B2(n674), .ZN(n12300)
         );
  OAI22_X1 U5016 ( .A1(n7432), .A2(n673), .B1(n14751), .B2(n674), .ZN(n12301)
         );
  OAI22_X1 U5017 ( .A1(n7416), .A2(n673), .B1(n14711), .B2(n674), .ZN(n12302)
         );
  OAI22_X1 U5018 ( .A1(n7400), .A2(n673), .B1(n14671), .B2(n674), .ZN(n12303)
         );
  OAI22_X1 U5019 ( .A1(n7384), .A2(n675), .B1(n14938), .B2(n676), .ZN(n12304)
         );
  OAI22_X1 U5020 ( .A1(n7368), .A2(n675), .B1(n14911), .B2(n676), .ZN(n12305)
         );
  OAI22_X1 U5021 ( .A1(n7352), .A2(n675), .B1(n14871), .B2(n676), .ZN(n12306)
         );
  OAI22_X1 U5022 ( .A1(n7336), .A2(n675), .B1(n14831), .B2(n676), .ZN(n12307)
         );
  OAI22_X1 U5023 ( .A1(n7320), .A2(n675), .B1(n14791), .B2(n676), .ZN(n12308)
         );
  OAI22_X1 U5024 ( .A1(n7304), .A2(n675), .B1(n14751), .B2(n676), .ZN(n12309)
         );
  OAI22_X1 U5025 ( .A1(n7288), .A2(n675), .B1(n14711), .B2(n676), .ZN(n12310)
         );
  OAI22_X1 U5026 ( .A1(n7272), .A2(n675), .B1(n14671), .B2(n676), .ZN(n12311)
         );
  OAI22_X1 U5027 ( .A1(n7256), .A2(n677), .B1(n14938), .B2(n678), .ZN(n12312)
         );
  OAI22_X1 U5028 ( .A1(n7240), .A2(n677), .B1(n14911), .B2(n678), .ZN(n12313)
         );
  OAI22_X1 U5029 ( .A1(n7224), .A2(n677), .B1(n14871), .B2(n678), .ZN(n12314)
         );
  OAI22_X1 U5030 ( .A1(n7208), .A2(n677), .B1(n14831), .B2(n678), .ZN(n12315)
         );
  OAI22_X1 U5031 ( .A1(n7192), .A2(n677), .B1(n14791), .B2(n678), .ZN(n12316)
         );
  OAI22_X1 U5032 ( .A1(n7176), .A2(n677), .B1(n14751), .B2(n678), .ZN(n12317)
         );
  OAI22_X1 U5033 ( .A1(n7160), .A2(n677), .B1(n14711), .B2(n678), .ZN(n12318)
         );
  OAI22_X1 U5034 ( .A1(n7144), .A2(n677), .B1(n14671), .B2(n678), .ZN(n12319)
         );
  OAI22_X1 U5035 ( .A1(n7128), .A2(n679), .B1(n14938), .B2(n680), .ZN(n12320)
         );
  OAI22_X1 U5036 ( .A1(n7112), .A2(n679), .B1(n14911), .B2(n680), .ZN(n12321)
         );
  OAI22_X1 U5037 ( .A1(n7096), .A2(n679), .B1(n14871), .B2(n680), .ZN(n12322)
         );
  OAI22_X1 U5038 ( .A1(n7080), .A2(n679), .B1(n14831), .B2(n680), .ZN(n12323)
         );
  OAI22_X1 U5039 ( .A1(n7064), .A2(n679), .B1(n14791), .B2(n680), .ZN(n12324)
         );
  OAI22_X1 U5040 ( .A1(n7048), .A2(n679), .B1(n14751), .B2(n680), .ZN(n12325)
         );
  OAI22_X1 U5041 ( .A1(n7032), .A2(n679), .B1(n14711), .B2(n680), .ZN(n12326)
         );
  OAI22_X1 U5042 ( .A1(n7016), .A2(n679), .B1(n14671), .B2(n680), .ZN(n12327)
         );
  OAI22_X1 U5043 ( .A1(n7000), .A2(n681), .B1(n14938), .B2(n682), .ZN(n12328)
         );
  OAI22_X1 U5044 ( .A1(n6984), .A2(n681), .B1(n14911), .B2(n682), .ZN(n12329)
         );
  OAI22_X1 U5045 ( .A1(n6968), .A2(n681), .B1(n14871), .B2(n682), .ZN(n12330)
         );
  OAI22_X1 U5046 ( .A1(n6952), .A2(n681), .B1(n14831), .B2(n682), .ZN(n12331)
         );
  OAI22_X1 U5047 ( .A1(n6936), .A2(n681), .B1(n14791), .B2(n682), .ZN(n12332)
         );
  OAI22_X1 U5048 ( .A1(n6920), .A2(n681), .B1(n14751), .B2(n682), .ZN(n12333)
         );
  OAI22_X1 U5049 ( .A1(n6904), .A2(n681), .B1(n14711), .B2(n682), .ZN(n12334)
         );
  OAI22_X1 U5050 ( .A1(n6888), .A2(n681), .B1(n14671), .B2(n682), .ZN(n12335)
         );
  OAI22_X1 U5051 ( .A1(n6872), .A2(n683), .B1(n14938), .B2(n684), .ZN(n12336)
         );
  OAI22_X1 U5052 ( .A1(n6856), .A2(n683), .B1(n14911), .B2(n684), .ZN(n12337)
         );
  OAI22_X1 U5053 ( .A1(n6840), .A2(n683), .B1(n14871), .B2(n684), .ZN(n12338)
         );
  OAI22_X1 U5054 ( .A1(n6824), .A2(n683), .B1(n14831), .B2(n684), .ZN(n12339)
         );
  OAI22_X1 U5055 ( .A1(n6808), .A2(n683), .B1(n14791), .B2(n684), .ZN(n12340)
         );
  OAI22_X1 U5056 ( .A1(n6792), .A2(n683), .B1(n14751), .B2(n684), .ZN(n12341)
         );
  OAI22_X1 U5057 ( .A1(n6776), .A2(n683), .B1(n14711), .B2(n684), .ZN(n12342)
         );
  OAI22_X1 U5058 ( .A1(n6760), .A2(n683), .B1(n14671), .B2(n684), .ZN(n12343)
         );
  OAI22_X1 U5059 ( .A1(n10076), .A2(n698), .B1(n14937), .B2(n699), .ZN(n12392)
         );
  OAI22_X1 U5060 ( .A1(n10060), .A2(n698), .B1(n14912), .B2(n699), .ZN(n12393)
         );
  OAI22_X1 U5061 ( .A1(n10044), .A2(n698), .B1(n14872), .B2(n699), .ZN(n12394)
         );
  OAI22_X1 U5062 ( .A1(n10028), .A2(n698), .B1(n14832), .B2(n699), .ZN(n12395)
         );
  OAI22_X1 U5063 ( .A1(n10012), .A2(n698), .B1(n14792), .B2(n699), .ZN(n12396)
         );
  OAI22_X1 U5064 ( .A1(n9996), .A2(n698), .B1(n14752), .B2(n699), .ZN(n12397)
         );
  OAI22_X1 U5065 ( .A1(n9980), .A2(n698), .B1(n14712), .B2(n699), .ZN(n12398)
         );
  OAI22_X1 U5066 ( .A1(n9964), .A2(n698), .B1(n14672), .B2(n699), .ZN(n12399)
         );
  OAI22_X1 U5067 ( .A1(n9948), .A2(n701), .B1(n14937), .B2(n702), .ZN(n12400)
         );
  OAI22_X1 U5068 ( .A1(n9932), .A2(n701), .B1(n14912), .B2(n702), .ZN(n12401)
         );
  OAI22_X1 U5069 ( .A1(n9916), .A2(n701), .B1(n14872), .B2(n702), .ZN(n12402)
         );
  OAI22_X1 U5070 ( .A1(n9900), .A2(n701), .B1(n14832), .B2(n702), .ZN(n12403)
         );
  OAI22_X1 U5071 ( .A1(n9884), .A2(n701), .B1(n14792), .B2(n702), .ZN(n12404)
         );
  OAI22_X1 U5072 ( .A1(n9868), .A2(n701), .B1(n14752), .B2(n702), .ZN(n12405)
         );
  OAI22_X1 U5073 ( .A1(n9852), .A2(n701), .B1(n14712), .B2(n702), .ZN(n12406)
         );
  OAI22_X1 U5074 ( .A1(n9836), .A2(n701), .B1(n14672), .B2(n702), .ZN(n12407)
         );
  OAI22_X1 U5075 ( .A1(n9820), .A2(n703), .B1(n14937), .B2(n704), .ZN(n12408)
         );
  OAI22_X1 U5076 ( .A1(n9804), .A2(n703), .B1(n14912), .B2(n704), .ZN(n12409)
         );
  OAI22_X1 U5077 ( .A1(n9788), .A2(n703), .B1(n14872), .B2(n704), .ZN(n12410)
         );
  OAI22_X1 U5078 ( .A1(n9772), .A2(n703), .B1(n14832), .B2(n704), .ZN(n12411)
         );
  OAI22_X1 U5079 ( .A1(n9756), .A2(n703), .B1(n14792), .B2(n704), .ZN(n12412)
         );
  OAI22_X1 U5080 ( .A1(n9740), .A2(n703), .B1(n14752), .B2(n704), .ZN(n12413)
         );
  OAI22_X1 U5081 ( .A1(n9724), .A2(n703), .B1(n14712), .B2(n704), .ZN(n12414)
         );
  OAI22_X1 U5082 ( .A1(n9708), .A2(n703), .B1(n14672), .B2(n704), .ZN(n12415)
         );
  OAI22_X1 U5083 ( .A1(n9692), .A2(n705), .B1(n14937), .B2(n706), .ZN(n12416)
         );
  OAI22_X1 U5084 ( .A1(n9676), .A2(n705), .B1(n14912), .B2(n706), .ZN(n12417)
         );
  OAI22_X1 U5085 ( .A1(n9660), .A2(n705), .B1(n14872), .B2(n706), .ZN(n12418)
         );
  OAI22_X1 U5086 ( .A1(n9644), .A2(n705), .B1(n14832), .B2(n706), .ZN(n12419)
         );
  OAI22_X1 U5087 ( .A1(n9628), .A2(n705), .B1(n14792), .B2(n706), .ZN(n12420)
         );
  OAI22_X1 U5088 ( .A1(n9612), .A2(n705), .B1(n14752), .B2(n706), .ZN(n12421)
         );
  OAI22_X1 U5089 ( .A1(n9596), .A2(n705), .B1(n14712), .B2(n706), .ZN(n12422)
         );
  OAI22_X1 U5090 ( .A1(n9580), .A2(n705), .B1(n14672), .B2(n706), .ZN(n12423)
         );
  OAI22_X1 U5091 ( .A1(n9564), .A2(n707), .B1(n14937), .B2(n708), .ZN(n12424)
         );
  OAI22_X1 U5092 ( .A1(n9548), .A2(n707), .B1(n14912), .B2(n708), .ZN(n12425)
         );
  OAI22_X1 U5093 ( .A1(n9532), .A2(n707), .B1(n14872), .B2(n708), .ZN(n12426)
         );
  OAI22_X1 U5094 ( .A1(n9516), .A2(n707), .B1(n14832), .B2(n708), .ZN(n12427)
         );
  OAI22_X1 U5095 ( .A1(n9500), .A2(n707), .B1(n14792), .B2(n708), .ZN(n12428)
         );
  OAI22_X1 U5096 ( .A1(n9484), .A2(n707), .B1(n14752), .B2(n708), .ZN(n12429)
         );
  OAI22_X1 U5097 ( .A1(n9468), .A2(n707), .B1(n14712), .B2(n708), .ZN(n12430)
         );
  OAI22_X1 U5098 ( .A1(n9452), .A2(n707), .B1(n14672), .B2(n708), .ZN(n12431)
         );
  OAI22_X1 U5099 ( .A1(n9436), .A2(n709), .B1(n14937), .B2(n710), .ZN(n12432)
         );
  OAI22_X1 U5100 ( .A1(n9420), .A2(n709), .B1(n14912), .B2(n710), .ZN(n12433)
         );
  OAI22_X1 U5101 ( .A1(n9404), .A2(n709), .B1(n14872), .B2(n710), .ZN(n12434)
         );
  OAI22_X1 U5102 ( .A1(n9388), .A2(n709), .B1(n14832), .B2(n710), .ZN(n12435)
         );
  OAI22_X1 U5103 ( .A1(n9372), .A2(n709), .B1(n14792), .B2(n710), .ZN(n12436)
         );
  OAI22_X1 U5104 ( .A1(n9356), .A2(n709), .B1(n14752), .B2(n710), .ZN(n12437)
         );
  OAI22_X1 U5105 ( .A1(n9340), .A2(n709), .B1(n14712), .B2(n710), .ZN(n12438)
         );
  OAI22_X1 U5106 ( .A1(n9324), .A2(n709), .B1(n14672), .B2(n710), .ZN(n12439)
         );
  OAI22_X1 U5107 ( .A1(n9308), .A2(n711), .B1(n14937), .B2(n712), .ZN(n12440)
         );
  OAI22_X1 U5108 ( .A1(n9292), .A2(n711), .B1(n14912), .B2(n712), .ZN(n12441)
         );
  OAI22_X1 U5109 ( .A1(n9276), .A2(n711), .B1(n14872), .B2(n712), .ZN(n12442)
         );
  OAI22_X1 U5110 ( .A1(n9260), .A2(n711), .B1(n14832), .B2(n712), .ZN(n12443)
         );
  OAI22_X1 U5111 ( .A1(n9244), .A2(n711), .B1(n14792), .B2(n712), .ZN(n12444)
         );
  OAI22_X1 U5112 ( .A1(n9228), .A2(n711), .B1(n14752), .B2(n712), .ZN(n12445)
         );
  OAI22_X1 U5113 ( .A1(n9212), .A2(n711), .B1(n14712), .B2(n712), .ZN(n12446)
         );
  OAI22_X1 U5114 ( .A1(n9196), .A2(n711), .B1(n14672), .B2(n712), .ZN(n12447)
         );
  OAI22_X1 U5115 ( .A1(n9180), .A2(n713), .B1(n14936), .B2(n714), .ZN(n12448)
         );
  OAI22_X1 U5116 ( .A1(n9164), .A2(n713), .B1(n14912), .B2(n714), .ZN(n12449)
         );
  OAI22_X1 U5117 ( .A1(n9148), .A2(n713), .B1(n14872), .B2(n714), .ZN(n12450)
         );
  OAI22_X1 U5118 ( .A1(n9132), .A2(n713), .B1(n14832), .B2(n714), .ZN(n12451)
         );
  OAI22_X1 U5119 ( .A1(n9116), .A2(n713), .B1(n14792), .B2(n714), .ZN(n12452)
         );
  OAI22_X1 U5120 ( .A1(n9100), .A2(n713), .B1(n14752), .B2(n714), .ZN(n12453)
         );
  OAI22_X1 U5121 ( .A1(n9084), .A2(n713), .B1(n14712), .B2(n714), .ZN(n12454)
         );
  OAI22_X1 U5122 ( .A1(n9068), .A2(n713), .B1(n14672), .B2(n714), .ZN(n12455)
         );
  OAI22_X1 U5123 ( .A1(n9052), .A2(n715), .B1(n14936), .B2(n716), .ZN(n12456)
         );
  OAI22_X1 U5124 ( .A1(n9036), .A2(n715), .B1(n14912), .B2(n716), .ZN(n12457)
         );
  OAI22_X1 U5125 ( .A1(n9020), .A2(n715), .B1(n14872), .B2(n716), .ZN(n12458)
         );
  OAI22_X1 U5126 ( .A1(n9004), .A2(n715), .B1(n14832), .B2(n716), .ZN(n12459)
         );
  OAI22_X1 U5127 ( .A1(n8988), .A2(n715), .B1(n14792), .B2(n716), .ZN(n12460)
         );
  OAI22_X1 U5128 ( .A1(n8972), .A2(n715), .B1(n14752), .B2(n716), .ZN(n12461)
         );
  OAI22_X1 U5129 ( .A1(n8956), .A2(n715), .B1(n14712), .B2(n716), .ZN(n12462)
         );
  OAI22_X1 U5130 ( .A1(n8940), .A2(n715), .B1(n14672), .B2(n716), .ZN(n12463)
         );
  OAI22_X1 U5131 ( .A1(n8924), .A2(n717), .B1(n14936), .B2(n718), .ZN(n12464)
         );
  OAI22_X1 U5132 ( .A1(n8908), .A2(n717), .B1(n14912), .B2(n718), .ZN(n12465)
         );
  OAI22_X1 U5133 ( .A1(n8892), .A2(n717), .B1(n14872), .B2(n718), .ZN(n12466)
         );
  OAI22_X1 U5134 ( .A1(n8876), .A2(n717), .B1(n14832), .B2(n718), .ZN(n12467)
         );
  OAI22_X1 U5135 ( .A1(n8860), .A2(n717), .B1(n14792), .B2(n718), .ZN(n12468)
         );
  OAI22_X1 U5136 ( .A1(n8844), .A2(n717), .B1(n14752), .B2(n718), .ZN(n12469)
         );
  OAI22_X1 U5137 ( .A1(n8828), .A2(n717), .B1(n14712), .B2(n718), .ZN(n12470)
         );
  OAI22_X1 U5138 ( .A1(n8812), .A2(n717), .B1(n14672), .B2(n718), .ZN(n12471)
         );
  OAI22_X1 U5139 ( .A1(n8796), .A2(n719), .B1(n14936), .B2(n720), .ZN(n12472)
         );
  OAI22_X1 U5140 ( .A1(n8780), .A2(n719), .B1(n14912), .B2(n720), .ZN(n12473)
         );
  OAI22_X1 U5141 ( .A1(n8764), .A2(n719), .B1(n14872), .B2(n720), .ZN(n12474)
         );
  OAI22_X1 U5142 ( .A1(n8748), .A2(n719), .B1(n14832), .B2(n720), .ZN(n12475)
         );
  OAI22_X1 U5143 ( .A1(n8732), .A2(n719), .B1(n14792), .B2(n720), .ZN(n12476)
         );
  OAI22_X1 U5144 ( .A1(n8716), .A2(n719), .B1(n14752), .B2(n720), .ZN(n12477)
         );
  OAI22_X1 U5145 ( .A1(n8700), .A2(n719), .B1(n14712), .B2(n720), .ZN(n12478)
         );
  OAI22_X1 U5146 ( .A1(n8684), .A2(n719), .B1(n14672), .B2(n720), .ZN(n12479)
         );
  OAI22_X1 U5147 ( .A1(n8668), .A2(n721), .B1(n14936), .B2(n722), .ZN(n12480)
         );
  OAI22_X1 U5148 ( .A1(n8652), .A2(n721), .B1(n14913), .B2(n722), .ZN(n12481)
         );
  OAI22_X1 U5149 ( .A1(n8636), .A2(n721), .B1(n14873), .B2(n722), .ZN(n12482)
         );
  OAI22_X1 U5150 ( .A1(n8620), .A2(n721), .B1(n14833), .B2(n722), .ZN(n12483)
         );
  OAI22_X1 U5151 ( .A1(n8604), .A2(n721), .B1(n14793), .B2(n722), .ZN(n12484)
         );
  OAI22_X1 U5152 ( .A1(n8588), .A2(n721), .B1(n14753), .B2(n722), .ZN(n12485)
         );
  OAI22_X1 U5153 ( .A1(n8572), .A2(n721), .B1(n14713), .B2(n722), .ZN(n12486)
         );
  OAI22_X1 U5154 ( .A1(n8556), .A2(n721), .B1(n14673), .B2(n722), .ZN(n12487)
         );
  OAI22_X1 U5155 ( .A1(n8540), .A2(n723), .B1(n14936), .B2(n724), .ZN(n12488)
         );
  OAI22_X1 U5156 ( .A1(n8524), .A2(n723), .B1(n14913), .B2(n724), .ZN(n12489)
         );
  OAI22_X1 U5157 ( .A1(n8508), .A2(n723), .B1(n14873), .B2(n724), .ZN(n12490)
         );
  OAI22_X1 U5158 ( .A1(n8492), .A2(n723), .B1(n14833), .B2(n724), .ZN(n12491)
         );
  OAI22_X1 U5159 ( .A1(n8476), .A2(n723), .B1(n14793), .B2(n724), .ZN(n12492)
         );
  OAI22_X1 U5160 ( .A1(n8460), .A2(n723), .B1(n14753), .B2(n724), .ZN(n12493)
         );
  OAI22_X1 U5161 ( .A1(n8444), .A2(n723), .B1(n14713), .B2(n724), .ZN(n12494)
         );
  OAI22_X1 U5162 ( .A1(n8428), .A2(n723), .B1(n14673), .B2(n724), .ZN(n12495)
         );
  OAI22_X1 U5163 ( .A1(n8412), .A2(n725), .B1(n14936), .B2(n726), .ZN(n12496)
         );
  OAI22_X1 U5164 ( .A1(n8396), .A2(n725), .B1(n14913), .B2(n726), .ZN(n12497)
         );
  OAI22_X1 U5165 ( .A1(n8380), .A2(n725), .B1(n14873), .B2(n726), .ZN(n12498)
         );
  OAI22_X1 U5166 ( .A1(n8364), .A2(n725), .B1(n14833), .B2(n726), .ZN(n12499)
         );
  OAI22_X1 U5167 ( .A1(n8348), .A2(n725), .B1(n14793), .B2(n726), .ZN(n12500)
         );
  OAI22_X1 U5168 ( .A1(n8332), .A2(n725), .B1(n14753), .B2(n726), .ZN(n12501)
         );
  OAI22_X1 U5169 ( .A1(n8316), .A2(n725), .B1(n14713), .B2(n726), .ZN(n12502)
         );
  OAI22_X1 U5170 ( .A1(n8300), .A2(n725), .B1(n14673), .B2(n726), .ZN(n12503)
         );
  OAI22_X1 U5171 ( .A1(n8284), .A2(n727), .B1(n14936), .B2(n728), .ZN(n12504)
         );
  OAI22_X1 U5172 ( .A1(n8268), .A2(n727), .B1(n14913), .B2(n728), .ZN(n12505)
         );
  OAI22_X1 U5173 ( .A1(n8252), .A2(n727), .B1(n14873), .B2(n728), .ZN(n12506)
         );
  OAI22_X1 U5174 ( .A1(n8236), .A2(n727), .B1(n14833), .B2(n728), .ZN(n12507)
         );
  OAI22_X1 U5175 ( .A1(n8220), .A2(n727), .B1(n14793), .B2(n728), .ZN(n12508)
         );
  OAI22_X1 U5176 ( .A1(n8204), .A2(n727), .B1(n14753), .B2(n728), .ZN(n12509)
         );
  OAI22_X1 U5177 ( .A1(n8188), .A2(n727), .B1(n14713), .B2(n728), .ZN(n12510)
         );
  OAI22_X1 U5178 ( .A1(n8172), .A2(n727), .B1(n14673), .B2(n728), .ZN(n12511)
         );
  OAI22_X1 U5179 ( .A1(n8156), .A2(n729), .B1(n14936), .B2(n730), .ZN(n12512)
         );
  OAI22_X1 U5180 ( .A1(n8140), .A2(n729), .B1(n14913), .B2(n730), .ZN(n12513)
         );
  OAI22_X1 U5181 ( .A1(n8124), .A2(n729), .B1(n14873), .B2(n730), .ZN(n12514)
         );
  OAI22_X1 U5182 ( .A1(n8108), .A2(n729), .B1(n14833), .B2(n730), .ZN(n12515)
         );
  OAI22_X1 U5183 ( .A1(n8092), .A2(n729), .B1(n14793), .B2(n730), .ZN(n12516)
         );
  OAI22_X1 U5185 ( .A1(n8076), .A2(n729), .B1(n14753), .B2(n730), .ZN(n12517)
         );
  OAI22_X1 U5186 ( .A1(n8060), .A2(n729), .B1(n14713), .B2(n730), .ZN(n12518)
         );
  OAI22_X1 U5187 ( .A1(n8044), .A2(n729), .B1(n14673), .B2(n730), .ZN(n12519)
         );
  OAI22_X1 U5188 ( .A1(n8028), .A2(n731), .B1(n14936), .B2(n732), .ZN(n12520)
         );
  OAI22_X1 U5189 ( .A1(n8012), .A2(n731), .B1(n14913), .B2(n732), .ZN(n12521)
         );
  OAI22_X1 U5190 ( .A1(n7996), .A2(n731), .B1(n14873), .B2(n732), .ZN(n12522)
         );
  OAI22_X1 U5191 ( .A1(n7980), .A2(n731), .B1(n14833), .B2(n732), .ZN(n12523)
         );
  OAI22_X1 U5192 ( .A1(n7964), .A2(n731), .B1(n14793), .B2(n732), .ZN(n12524)
         );
  OAI22_X1 U5193 ( .A1(n7948), .A2(n731), .B1(n14753), .B2(n732), .ZN(n12525)
         );
  OAI22_X1 U5194 ( .A1(n7932), .A2(n731), .B1(n14713), .B2(n732), .ZN(n12526)
         );
  OAI22_X1 U5195 ( .A1(n7916), .A2(n731), .B1(n14673), .B2(n732), .ZN(n12527)
         );
  OAI22_X1 U5196 ( .A1(n7900), .A2(n733), .B1(n14936), .B2(n734), .ZN(n12528)
         );
  OAI22_X1 U5197 ( .A1(n7884), .A2(n733), .B1(n14913), .B2(n734), .ZN(n12529)
         );
  OAI22_X1 U5198 ( .A1(n7868), .A2(n733), .B1(n14873), .B2(n734), .ZN(n12530)
         );
  OAI22_X1 U5199 ( .A1(n7852), .A2(n733), .B1(n14833), .B2(n734), .ZN(n12531)
         );
  OAI22_X1 U5200 ( .A1(n7836), .A2(n733), .B1(n14793), .B2(n734), .ZN(n12532)
         );
  OAI22_X1 U5201 ( .A1(n7820), .A2(n733), .B1(n14753), .B2(n734), .ZN(n12533)
         );
  OAI22_X1 U5202 ( .A1(n7804), .A2(n733), .B1(n14713), .B2(n734), .ZN(n12534)
         );
  OAI22_X1 U5203 ( .A1(n7788), .A2(n733), .B1(n14673), .B2(n734), .ZN(n12535)
         );
  OAI22_X1 U5204 ( .A1(n7772), .A2(n735), .B1(n14936), .B2(n736), .ZN(n12536)
         );
  OAI22_X1 U5205 ( .A1(n7756), .A2(n735), .B1(n14913), .B2(n736), .ZN(n12537)
         );
  OAI22_X1 U5206 ( .A1(n7740), .A2(n735), .B1(n14873), .B2(n736), .ZN(n12538)
         );
  OAI22_X1 U5207 ( .A1(n7724), .A2(n735), .B1(n14833), .B2(n736), .ZN(n12539)
         );
  OAI22_X1 U5208 ( .A1(n7708), .A2(n735), .B1(n14793), .B2(n736), .ZN(n12540)
         );
  OAI22_X1 U5209 ( .A1(n7692), .A2(n735), .B1(n14753), .B2(n736), .ZN(n12541)
         );
  OAI22_X1 U5210 ( .A1(n7676), .A2(n735), .B1(n14713), .B2(n736), .ZN(n12542)
         );
  OAI22_X1 U5211 ( .A1(n7660), .A2(n735), .B1(n14673), .B2(n736), .ZN(n12543)
         );
  OAI22_X1 U5212 ( .A1(n7644), .A2(n737), .B1(n14936), .B2(n738), .ZN(n12544)
         );
  OAI22_X1 U5213 ( .A1(n7628), .A2(n737), .B1(n14913), .B2(n738), .ZN(n12545)
         );
  OAI22_X1 U5214 ( .A1(n7612), .A2(n737), .B1(n14873), .B2(n738), .ZN(n12546)
         );
  OAI22_X1 U5215 ( .A1(n7596), .A2(n737), .B1(n14833), .B2(n738), .ZN(n12547)
         );
  OAI22_X1 U5216 ( .A1(n7580), .A2(n737), .B1(n14793), .B2(n738), .ZN(n12548)
         );
  OAI22_X1 U5217 ( .A1(n7564), .A2(n737), .B1(n14753), .B2(n738), .ZN(n12549)
         );
  OAI22_X1 U5218 ( .A1(n7548), .A2(n737), .B1(n14713), .B2(n738), .ZN(n12550)
         );
  OAI22_X1 U5219 ( .A1(n7532), .A2(n737), .B1(n14673), .B2(n738), .ZN(n12551)
         );
  OAI22_X1 U5220 ( .A1(n7516), .A2(n739), .B1(n14935), .B2(n740), .ZN(n12552)
         );
  OAI22_X1 U5221 ( .A1(n7500), .A2(n739), .B1(n14913), .B2(n740), .ZN(n12553)
         );
  OAI22_X1 U5222 ( .A1(n7484), .A2(n739), .B1(n14873), .B2(n740), .ZN(n12554)
         );
  OAI22_X1 U5223 ( .A1(n7468), .A2(n739), .B1(n14833), .B2(n740), .ZN(n12555)
         );
  OAI22_X1 U5224 ( .A1(n7452), .A2(n739), .B1(n14793), .B2(n740), .ZN(n12556)
         );
  OAI22_X1 U5225 ( .A1(n7436), .A2(n739), .B1(n14753), .B2(n740), .ZN(n12557)
         );
  OAI22_X1 U5226 ( .A1(n7420), .A2(n739), .B1(n14713), .B2(n740), .ZN(n12558)
         );
  OAI22_X1 U5227 ( .A1(n7404), .A2(n739), .B1(n14673), .B2(n740), .ZN(n12559)
         );
  OAI22_X1 U5228 ( .A1(n7388), .A2(n741), .B1(n14935), .B2(n742), .ZN(n12560)
         );
  OAI22_X1 U5229 ( .A1(n7372), .A2(n741), .B1(n14913), .B2(n742), .ZN(n12561)
         );
  OAI22_X1 U5230 ( .A1(n7356), .A2(n741), .B1(n14873), .B2(n742), .ZN(n12562)
         );
  OAI22_X1 U5231 ( .A1(n7340), .A2(n741), .B1(n14833), .B2(n742), .ZN(n12563)
         );
  OAI22_X1 U5232 ( .A1(n7324), .A2(n741), .B1(n14793), .B2(n742), .ZN(n12564)
         );
  OAI22_X1 U5233 ( .A1(n7308), .A2(n741), .B1(n14753), .B2(n742), .ZN(n12565)
         );
  OAI22_X1 U5234 ( .A1(n7292), .A2(n741), .B1(n14713), .B2(n742), .ZN(n12566)
         );
  OAI22_X1 U5235 ( .A1(n7276), .A2(n741), .B1(n14673), .B2(n742), .ZN(n12567)
         );
  OAI22_X1 U5236 ( .A1(n7260), .A2(n743), .B1(n14935), .B2(n744), .ZN(n12568)
         );
  OAI22_X1 U5237 ( .A1(n7244), .A2(n743), .B1(n14913), .B2(n744), .ZN(n12569)
         );
  OAI22_X1 U5238 ( .A1(n7228), .A2(n743), .B1(n14873), .B2(n744), .ZN(n12570)
         );
  OAI22_X1 U5239 ( .A1(n7212), .A2(n743), .B1(n14833), .B2(n744), .ZN(n12571)
         );
  OAI22_X1 U5240 ( .A1(n7196), .A2(n743), .B1(n14793), .B2(n744), .ZN(n12572)
         );
  OAI22_X1 U5241 ( .A1(n7180), .A2(n743), .B1(n14753), .B2(n744), .ZN(n12573)
         );
  OAI22_X1 U5242 ( .A1(n7164), .A2(n743), .B1(n14713), .B2(n744), .ZN(n12574)
         );
  OAI22_X1 U5243 ( .A1(n7148), .A2(n743), .B1(n14673), .B2(n744), .ZN(n12575)
         );
  OAI22_X1 U5244 ( .A1(n7132), .A2(n745), .B1(n14935), .B2(n746), .ZN(n12576)
         );
  OAI22_X1 U5245 ( .A1(n7116), .A2(n745), .B1(n14913), .B2(n746), .ZN(n12577)
         );
  OAI22_X1 U5246 ( .A1(n7100), .A2(n745), .B1(n14873), .B2(n746), .ZN(n12578)
         );
  OAI22_X1 U5247 ( .A1(n7084), .A2(n745), .B1(n14833), .B2(n746), .ZN(n12579)
         );
  OAI22_X1 U5248 ( .A1(n7068), .A2(n745), .B1(n14793), .B2(n746), .ZN(n12580)
         );
  OAI22_X1 U5249 ( .A1(n7052), .A2(n745), .B1(n14753), .B2(n746), .ZN(n12581)
         );
  OAI22_X1 U5250 ( .A1(n7036), .A2(n745), .B1(n14713), .B2(n746), .ZN(n12582)
         );
  OAI22_X1 U5251 ( .A1(n7020), .A2(n745), .B1(n14673), .B2(n746), .ZN(n12583)
         );
  OAI22_X1 U5252 ( .A1(n7004), .A2(n747), .B1(n14935), .B2(n748), .ZN(n12584)
         );
  OAI22_X1 U5253 ( .A1(n6988), .A2(n747), .B1(n14914), .B2(n748), .ZN(n12585)
         );
  OAI22_X1 U5254 ( .A1(n6972), .A2(n747), .B1(n14874), .B2(n748), .ZN(n12586)
         );
  OAI22_X1 U5255 ( .A1(n6956), .A2(n747), .B1(n14834), .B2(n748), .ZN(n12587)
         );
  OAI22_X1 U5256 ( .A1(n6940), .A2(n747), .B1(n14794), .B2(n748), .ZN(n12588)
         );
  OAI22_X1 U5257 ( .A1(n6924), .A2(n747), .B1(n14754), .B2(n748), .ZN(n12589)
         );
  OAI22_X1 U5258 ( .A1(n6908), .A2(n747), .B1(n14714), .B2(n748), .ZN(n12590)
         );
  OAI22_X1 U5259 ( .A1(n6892), .A2(n747), .B1(n14674), .B2(n748), .ZN(n12591)
         );
  OAI22_X1 U5260 ( .A1(n6876), .A2(n749), .B1(n14935), .B2(n750), .ZN(n12592)
         );
  OAI22_X1 U5261 ( .A1(n6860), .A2(n749), .B1(n14914), .B2(n750), .ZN(n12593)
         );
  OAI22_X1 U5262 ( .A1(n6844), .A2(n749), .B1(n14874), .B2(n750), .ZN(n12594)
         );
  OAI22_X1 U5263 ( .A1(n6828), .A2(n749), .B1(n14834), .B2(n750), .ZN(n12595)
         );
  OAI22_X1 U5264 ( .A1(n6812), .A2(n749), .B1(n14794), .B2(n750), .ZN(n12596)
         );
  OAI22_X1 U5265 ( .A1(n6796), .A2(n749), .B1(n14754), .B2(n750), .ZN(n12597)
         );
  OAI22_X1 U5266 ( .A1(n6780), .A2(n749), .B1(n14714), .B2(n750), .ZN(n12598)
         );
  OAI22_X1 U5267 ( .A1(n6764), .A2(n749), .B1(n14674), .B2(n750), .ZN(n12599)
         );
  OAI22_X1 U5268 ( .A1(n10080), .A2(n764), .B1(n14935), .B2(n765), .ZN(n12648)
         );
  OAI22_X1 U5269 ( .A1(n10064), .A2(n764), .B1(n14914), .B2(n765), .ZN(n12649)
         );
  OAI22_X1 U5270 ( .A1(n10048), .A2(n764), .B1(n14874), .B2(n765), .ZN(n12650)
         );
  OAI22_X1 U5271 ( .A1(n10032), .A2(n764), .B1(n14834), .B2(n765), .ZN(n12651)
         );
  OAI22_X1 U5272 ( .A1(n10016), .A2(n764), .B1(n14794), .B2(n765), .ZN(n12652)
         );
  OAI22_X1 U5273 ( .A1(n10000), .A2(n764), .B1(n14754), .B2(n765), .ZN(n12653)
         );
  OAI22_X1 U5274 ( .A1(n9984), .A2(n764), .B1(n14714), .B2(n765), .ZN(n12654)
         );
  OAI22_X1 U5275 ( .A1(n9968), .A2(n764), .B1(n14674), .B2(n765), .ZN(n12655)
         );
  OAI22_X1 U5276 ( .A1(n9952), .A2(n767), .B1(n14934), .B2(n768), .ZN(n12656)
         );
  OAI22_X1 U5277 ( .A1(n9936), .A2(n767), .B1(n14914), .B2(n768), .ZN(n12657)
         );
  OAI22_X1 U5278 ( .A1(n9920), .A2(n767), .B1(n14874), .B2(n768), .ZN(n12658)
         );
  OAI22_X1 U5279 ( .A1(n9904), .A2(n767), .B1(n14834), .B2(n768), .ZN(n12659)
         );
  OAI22_X1 U5280 ( .A1(n9888), .A2(n767), .B1(n14794), .B2(n768), .ZN(n12660)
         );
  OAI22_X1 U5281 ( .A1(n9872), .A2(n767), .B1(n14754), .B2(n768), .ZN(n12661)
         );
  OAI22_X1 U5282 ( .A1(n9856), .A2(n767), .B1(n14714), .B2(n768), .ZN(n12662)
         );
  OAI22_X1 U5283 ( .A1(n9840), .A2(n767), .B1(n14674), .B2(n768), .ZN(n12663)
         );
  OAI22_X1 U5284 ( .A1(n9824), .A2(n769), .B1(n14934), .B2(n770), .ZN(n12664)
         );
  OAI22_X1 U5285 ( .A1(n9808), .A2(n769), .B1(n14914), .B2(n770), .ZN(n12665)
         );
  OAI22_X1 U5286 ( .A1(n9792), .A2(n769), .B1(n14874), .B2(n770), .ZN(n12666)
         );
  OAI22_X1 U5287 ( .A1(n9776), .A2(n769), .B1(n14834), .B2(n770), .ZN(n12667)
         );
  OAI22_X1 U5288 ( .A1(n9760), .A2(n769), .B1(n14794), .B2(n770), .ZN(n12668)
         );
  OAI22_X1 U5289 ( .A1(n9744), .A2(n769), .B1(n14754), .B2(n770), .ZN(n12669)
         );
  OAI22_X1 U5290 ( .A1(n9728), .A2(n769), .B1(n14714), .B2(n770), .ZN(n12670)
         );
  OAI22_X1 U5291 ( .A1(n9712), .A2(n769), .B1(n14674), .B2(n770), .ZN(n12671)
         );
  OAI22_X1 U5292 ( .A1(n9696), .A2(n771), .B1(n14934), .B2(n772), .ZN(n12672)
         );
  OAI22_X1 U5293 ( .A1(n9680), .A2(n771), .B1(n14914), .B2(n772), .ZN(n12673)
         );
  OAI22_X1 U5294 ( .A1(n9664), .A2(n771), .B1(n14874), .B2(n772), .ZN(n12674)
         );
  OAI22_X1 U5295 ( .A1(n9648), .A2(n771), .B1(n14834), .B2(n772), .ZN(n12675)
         );
  OAI22_X1 U5296 ( .A1(n9632), .A2(n771), .B1(n14794), .B2(n772), .ZN(n12676)
         );
  OAI22_X1 U5297 ( .A1(n9616), .A2(n771), .B1(n14754), .B2(n772), .ZN(n12677)
         );
  OAI22_X1 U5298 ( .A1(n9600), .A2(n771), .B1(n14714), .B2(n772), .ZN(n12678)
         );
  OAI22_X1 U5299 ( .A1(n9584), .A2(n771), .B1(n14674), .B2(n772), .ZN(n12679)
         );
  OAI22_X1 U5300 ( .A1(n9568), .A2(n773), .B1(n14934), .B2(n774), .ZN(n12680)
         );
  OAI22_X1 U5301 ( .A1(n9552), .A2(n773), .B1(n14914), .B2(n774), .ZN(n12681)
         );
  OAI22_X1 U5302 ( .A1(n9536), .A2(n773), .B1(n14874), .B2(n774), .ZN(n12682)
         );
  OAI22_X1 U5303 ( .A1(n9520), .A2(n773), .B1(n14834), .B2(n774), .ZN(n12683)
         );
  OAI22_X1 U5304 ( .A1(n9504), .A2(n773), .B1(n14794), .B2(n774), .ZN(n12684)
         );
  OAI22_X1 U5305 ( .A1(n9488), .A2(n773), .B1(n14754), .B2(n774), .ZN(n12685)
         );
  OAI22_X1 U5306 ( .A1(n9472), .A2(n773), .B1(n14714), .B2(n774), .ZN(n12686)
         );
  OAI22_X1 U5307 ( .A1(n9456), .A2(n773), .B1(n14674), .B2(n774), .ZN(n12687)
         );
  OAI22_X1 U5308 ( .A1(n9440), .A2(n775), .B1(n14934), .B2(n776), .ZN(n12688)
         );
  OAI22_X1 U5309 ( .A1(n9424), .A2(n775), .B1(n14915), .B2(n776), .ZN(n12689)
         );
  OAI22_X1 U5310 ( .A1(n9408), .A2(n775), .B1(n14875), .B2(n776), .ZN(n12690)
         );
  OAI22_X1 U5311 ( .A1(n9392), .A2(n775), .B1(n14835), .B2(n776), .ZN(n12691)
         );
  OAI22_X1 U5312 ( .A1(n9376), .A2(n775), .B1(n14795), .B2(n776), .ZN(n12692)
         );
  OAI22_X1 U5313 ( .A1(n9360), .A2(n775), .B1(n14755), .B2(n776), .ZN(n12693)
         );
  OAI22_X1 U5314 ( .A1(n9344), .A2(n775), .B1(n14715), .B2(n776), .ZN(n12694)
         );
  OAI22_X1 U5315 ( .A1(n9328), .A2(n775), .B1(n14675), .B2(n776), .ZN(n12695)
         );
  OAI22_X1 U5316 ( .A1(n9312), .A2(n777), .B1(n14934), .B2(n778), .ZN(n12696)
         );
  OAI22_X1 U5317 ( .A1(n9296), .A2(n777), .B1(n14915), .B2(n778), .ZN(n12697)
         );
  OAI22_X1 U5318 ( .A1(n9280), .A2(n777), .B1(n14875), .B2(n778), .ZN(n12698)
         );
  OAI22_X1 U5319 ( .A1(n9264), .A2(n777), .B1(n14835), .B2(n778), .ZN(n12699)
         );
  OAI22_X1 U5320 ( .A1(n9248), .A2(n777), .B1(n14795), .B2(n778), .ZN(n12700)
         );
  OAI22_X1 U5321 ( .A1(n9232), .A2(n777), .B1(n14755), .B2(n778), .ZN(n12701)
         );
  OAI22_X1 U5322 ( .A1(n9216), .A2(n777), .B1(n14715), .B2(n778), .ZN(n12702)
         );
  OAI22_X1 U5323 ( .A1(n9200), .A2(n777), .B1(n14675), .B2(n778), .ZN(n12703)
         );
  OAI22_X1 U5324 ( .A1(n9184), .A2(n779), .B1(n14934), .B2(n780), .ZN(n12704)
         );
  OAI22_X1 U5325 ( .A1(n9168), .A2(n779), .B1(n14915), .B2(n780), .ZN(n12705)
         );
  OAI22_X1 U5326 ( .A1(n9152), .A2(n779), .B1(n14875), .B2(n780), .ZN(n12706)
         );
  OAI22_X1 U5327 ( .A1(n9136), .A2(n779), .B1(n14835), .B2(n780), .ZN(n12707)
         );
  OAI22_X1 U5328 ( .A1(n9120), .A2(n779), .B1(n14795), .B2(n780), .ZN(n12708)
         );
  OAI22_X1 U5329 ( .A1(n9104), .A2(n779), .B1(n14755), .B2(n780), .ZN(n12709)
         );
  OAI22_X1 U5330 ( .A1(n9088), .A2(n779), .B1(n14715), .B2(n780), .ZN(n12710)
         );
  OAI22_X1 U5331 ( .A1(n9072), .A2(n779), .B1(n14675), .B2(n780), .ZN(n12711)
         );
  OAI22_X1 U5332 ( .A1(n9056), .A2(n781), .B1(n14934), .B2(n782), .ZN(n12712)
         );
  OAI22_X1 U5333 ( .A1(n9040), .A2(n781), .B1(n14915), .B2(n782), .ZN(n12713)
         );
  OAI22_X1 U5334 ( .A1(n9024), .A2(n781), .B1(n14875), .B2(n782), .ZN(n12714)
         );
  OAI22_X1 U5335 ( .A1(n9008), .A2(n781), .B1(n14835), .B2(n782), .ZN(n12715)
         );
  OAI22_X1 U5337 ( .A1(n8992), .A2(n781), .B1(n14795), .B2(n782), .ZN(n12716)
         );
  OAI22_X1 U5338 ( .A1(n8976), .A2(n781), .B1(n14755), .B2(n782), .ZN(n12717)
         );
  OAI22_X1 U5339 ( .A1(n8960), .A2(n781), .B1(n14715), .B2(n782), .ZN(n12718)
         );
  OAI22_X1 U5340 ( .A1(n8944), .A2(n781), .B1(n14675), .B2(n782), .ZN(n12719)
         );
  OAI22_X1 U5341 ( .A1(n8928), .A2(n783), .B1(n14934), .B2(n784), .ZN(n12720)
         );
  OAI22_X1 U5342 ( .A1(n8912), .A2(n783), .B1(n14915), .B2(n784), .ZN(n12721)
         );
  OAI22_X1 U5343 ( .A1(n8896), .A2(n783), .B1(n14875), .B2(n784), .ZN(n12722)
         );
  OAI22_X1 U5344 ( .A1(n8880), .A2(n783), .B1(n14835), .B2(n784), .ZN(n12723)
         );
  OAI22_X1 U5345 ( .A1(n8864), .A2(n783), .B1(n14795), .B2(n784), .ZN(n12724)
         );
  OAI22_X1 U5346 ( .A1(n8848), .A2(n783), .B1(n14755), .B2(n784), .ZN(n12725)
         );
  OAI22_X1 U5347 ( .A1(n8832), .A2(n783), .B1(n14715), .B2(n784), .ZN(n12726)
         );
  OAI22_X1 U5348 ( .A1(n8816), .A2(n783), .B1(n14675), .B2(n784), .ZN(n12727)
         );
  OAI22_X1 U5349 ( .A1(n8800), .A2(n785), .B1(n14934), .B2(n786), .ZN(n12728)
         );
  OAI22_X1 U5350 ( .A1(n8784), .A2(n785), .B1(n14915), .B2(n786), .ZN(n12729)
         );
  OAI22_X1 U5351 ( .A1(n8768), .A2(n785), .B1(n14875), .B2(n786), .ZN(n12730)
         );
  OAI22_X1 U5352 ( .A1(n8752), .A2(n785), .B1(n14835), .B2(n786), .ZN(n12731)
         );
  OAI22_X1 U5353 ( .A1(n8736), .A2(n785), .B1(n14795), .B2(n786), .ZN(n12732)
         );
  OAI22_X1 U5354 ( .A1(n8720), .A2(n785), .B1(n14755), .B2(n786), .ZN(n12733)
         );
  OAI22_X1 U5355 ( .A1(n8704), .A2(n785), .B1(n14715), .B2(n786), .ZN(n12734)
         );
  OAI22_X1 U5356 ( .A1(n8688), .A2(n785), .B1(n14675), .B2(n786), .ZN(n12735)
         );
  OAI22_X1 U5357 ( .A1(n8672), .A2(n787), .B1(n14934), .B2(n788), .ZN(n12736)
         );
  OAI22_X1 U5358 ( .A1(n8656), .A2(n787), .B1(n14915), .B2(n788), .ZN(n12737)
         );
  OAI22_X1 U5359 ( .A1(n8640), .A2(n787), .B1(n14875), .B2(n788), .ZN(n12738)
         );
  OAI22_X1 U5360 ( .A1(n8624), .A2(n787), .B1(n14835), .B2(n788), .ZN(n12739)
         );
  OAI22_X1 U5361 ( .A1(n8608), .A2(n787), .B1(n14795), .B2(n788), .ZN(n12740)
         );
  OAI22_X1 U5362 ( .A1(n8592), .A2(n787), .B1(n14755), .B2(n788), .ZN(n12741)
         );
  OAI22_X1 U5363 ( .A1(n8576), .A2(n787), .B1(n14715), .B2(n788), .ZN(n12742)
         );
  OAI22_X1 U5364 ( .A1(n8560), .A2(n787), .B1(n14675), .B2(n788), .ZN(n12743)
         );
  OAI22_X1 U5365 ( .A1(n8544), .A2(n789), .B1(n14934), .B2(n790), .ZN(n12744)
         );
  OAI22_X1 U5366 ( .A1(n8528), .A2(n789), .B1(n14915), .B2(n790), .ZN(n12745)
         );
  OAI22_X1 U5367 ( .A1(n8512), .A2(n789), .B1(n14875), .B2(n790), .ZN(n12746)
         );
  OAI22_X1 U5368 ( .A1(n8496), .A2(n789), .B1(n14835), .B2(n790), .ZN(n12747)
         );
  OAI22_X1 U5369 ( .A1(n8480), .A2(n789), .B1(n14795), .B2(n790), .ZN(n12748)
         );
  OAI22_X1 U5370 ( .A1(n8464), .A2(n789), .B1(n14755), .B2(n790), .ZN(n12749)
         );
  OAI22_X1 U5371 ( .A1(n8448), .A2(n789), .B1(n14715), .B2(n790), .ZN(n12750)
         );
  OAI22_X1 U5372 ( .A1(n8432), .A2(n789), .B1(n14675), .B2(n790), .ZN(n12751)
         );
  OAI22_X1 U5373 ( .A1(n8416), .A2(n791), .B1(n14933), .B2(n792), .ZN(n12752)
         );
  OAI22_X1 U5374 ( .A1(n8400), .A2(n791), .B1(n14915), .B2(n792), .ZN(n12753)
         );
  OAI22_X1 U5375 ( .A1(n8384), .A2(n791), .B1(n14875), .B2(n792), .ZN(n12754)
         );
  OAI22_X1 U5376 ( .A1(n8368), .A2(n791), .B1(n14835), .B2(n792), .ZN(n12755)
         );
  OAI22_X1 U5377 ( .A1(n8352), .A2(n791), .B1(n14795), .B2(n792), .ZN(n12756)
         );
  OAI22_X1 U5378 ( .A1(n8336), .A2(n791), .B1(n14755), .B2(n792), .ZN(n12757)
         );
  OAI22_X1 U5379 ( .A1(n8320), .A2(n791), .B1(n14715), .B2(n792), .ZN(n12758)
         );
  OAI22_X1 U5380 ( .A1(n8304), .A2(n791), .B1(n14675), .B2(n792), .ZN(n12759)
         );
  OAI22_X1 U5381 ( .A1(n8288), .A2(n793), .B1(n14933), .B2(n794), .ZN(n12760)
         );
  OAI22_X1 U5382 ( .A1(n8272), .A2(n793), .B1(n14915), .B2(n794), .ZN(n12761)
         );
  OAI22_X1 U5383 ( .A1(n8256), .A2(n793), .B1(n14875), .B2(n794), .ZN(n12762)
         );
  OAI22_X1 U5384 ( .A1(n8240), .A2(n793), .B1(n14835), .B2(n794), .ZN(n12763)
         );
  OAI22_X1 U5385 ( .A1(n8224), .A2(n793), .B1(n14795), .B2(n794), .ZN(n12764)
         );
  OAI22_X1 U5386 ( .A1(n8208), .A2(n793), .B1(n14755), .B2(n794), .ZN(n12765)
         );
  OAI22_X1 U5387 ( .A1(n8192), .A2(n793), .B1(n14715), .B2(n794), .ZN(n12766)
         );
  OAI22_X1 U5388 ( .A1(n8176), .A2(n793), .B1(n14675), .B2(n794), .ZN(n12767)
         );
  OAI22_X1 U5389 ( .A1(n8160), .A2(n795), .B1(n14933), .B2(n796), .ZN(n12768)
         );
  OAI22_X1 U5390 ( .A1(n8144), .A2(n795), .B1(n14915), .B2(n796), .ZN(n12769)
         );
  OAI22_X1 U5391 ( .A1(n8128), .A2(n795), .B1(n14875), .B2(n796), .ZN(n12770)
         );
  OAI22_X1 U5392 ( .A1(n8112), .A2(n795), .B1(n14835), .B2(n796), .ZN(n12771)
         );
  OAI22_X1 U5393 ( .A1(n8096), .A2(n795), .B1(n14795), .B2(n796), .ZN(n12772)
         );
  OAI22_X1 U5394 ( .A1(n8080), .A2(n795), .B1(n14755), .B2(n796), .ZN(n12773)
         );
  OAI22_X1 U5395 ( .A1(n8064), .A2(n795), .B1(n14715), .B2(n796), .ZN(n12774)
         );
  OAI22_X1 U5396 ( .A1(n8048), .A2(n795), .B1(n14675), .B2(n796), .ZN(n12775)
         );
  OAI22_X1 U5397 ( .A1(n8032), .A2(n797), .B1(n14933), .B2(n798), .ZN(n12776)
         );
  OAI22_X1 U5398 ( .A1(n8016), .A2(n797), .B1(n14915), .B2(n798), .ZN(n12777)
         );
  OAI22_X1 U5399 ( .A1(n8000), .A2(n797), .B1(n14875), .B2(n798), .ZN(n12778)
         );
  OAI22_X1 U5400 ( .A1(n7984), .A2(n797), .B1(n14835), .B2(n798), .ZN(n12779)
         );
  OAI22_X1 U5401 ( .A1(n7968), .A2(n797), .B1(n14795), .B2(n798), .ZN(n12780)
         );
  OAI22_X1 U5402 ( .A1(n7952), .A2(n797), .B1(n14755), .B2(n798), .ZN(n12781)
         );
  OAI22_X1 U5403 ( .A1(n7936), .A2(n797), .B1(n14715), .B2(n798), .ZN(n12782)
         );
  OAI22_X1 U5404 ( .A1(n7920), .A2(n797), .B1(n14675), .B2(n798), .ZN(n12783)
         );
  OAI22_X1 U5405 ( .A1(n7904), .A2(n799), .B1(n14933), .B2(n800), .ZN(n12784)
         );
  OAI22_X1 U5406 ( .A1(n7888), .A2(n799), .B1(n14915), .B2(n800), .ZN(n12785)
         );
  OAI22_X1 U5407 ( .A1(n7872), .A2(n799), .B1(n14875), .B2(n800), .ZN(n12786)
         );
  OAI22_X1 U5408 ( .A1(n7856), .A2(n799), .B1(n14835), .B2(n800), .ZN(n12787)
         );
  OAI22_X1 U5409 ( .A1(n7840), .A2(n799), .B1(n14795), .B2(n800), .ZN(n12788)
         );
  OAI22_X1 U5410 ( .A1(n7824), .A2(n799), .B1(n14755), .B2(n800), .ZN(n12789)
         );
  OAI22_X1 U5411 ( .A1(n7808), .A2(n799), .B1(n14715), .B2(n800), .ZN(n12790)
         );
  OAI22_X1 U5412 ( .A1(n7792), .A2(n799), .B1(n14675), .B2(n800), .ZN(n12791)
         );
  OAI22_X1 U5413 ( .A1(n7776), .A2(n801), .B1(n14933), .B2(n802), .ZN(n12792)
         );
  OAI22_X1 U5414 ( .A1(n7760), .A2(n801), .B1(n14916), .B2(n802), .ZN(n12793)
         );
  OAI22_X1 U5415 ( .A1(n7744), .A2(n801), .B1(n14876), .B2(n802), .ZN(n12794)
         );
  OAI22_X1 U5416 ( .A1(n7728), .A2(n801), .B1(n14836), .B2(n802), .ZN(n12795)
         );
  OAI22_X1 U5417 ( .A1(n7712), .A2(n801), .B1(n14796), .B2(n802), .ZN(n12796)
         );
  OAI22_X1 U5418 ( .A1(n7696), .A2(n801), .B1(n14756), .B2(n802), .ZN(n12797)
         );
  OAI22_X1 U5419 ( .A1(n7680), .A2(n801), .B1(n14716), .B2(n802), .ZN(n12798)
         );
  OAI22_X1 U5420 ( .A1(n7664), .A2(n801), .B1(n14676), .B2(n802), .ZN(n12799)
         );
  OAI22_X1 U5421 ( .A1(n7648), .A2(n803), .B1(n14933), .B2(n804), .ZN(n12800)
         );
  OAI22_X1 U5422 ( .A1(n7632), .A2(n803), .B1(n14916), .B2(n804), .ZN(n12801)
         );
  OAI22_X1 U5423 ( .A1(n7616), .A2(n803), .B1(n14876), .B2(n804), .ZN(n12802)
         );
  OAI22_X1 U5424 ( .A1(n7600), .A2(n803), .B1(n14836), .B2(n804), .ZN(n12803)
         );
  OAI22_X1 U5425 ( .A1(n7584), .A2(n803), .B1(n14796), .B2(n804), .ZN(n12804)
         );
  OAI22_X1 U5426 ( .A1(n7568), .A2(n803), .B1(n14756), .B2(n804), .ZN(n12805)
         );
  OAI22_X1 U5427 ( .A1(n7552), .A2(n803), .B1(n14716), .B2(n804), .ZN(n12806)
         );
  OAI22_X1 U5428 ( .A1(n7536), .A2(n803), .B1(n14676), .B2(n804), .ZN(n12807)
         );
  OAI22_X1 U5429 ( .A1(n7520), .A2(n805), .B1(n14933), .B2(n806), .ZN(n12808)
         );
  OAI22_X1 U5430 ( .A1(n7504), .A2(n805), .B1(n14916), .B2(n806), .ZN(n12809)
         );
  OAI22_X1 U5431 ( .A1(n7488), .A2(n805), .B1(n14876), .B2(n806), .ZN(n12810)
         );
  OAI22_X1 U5432 ( .A1(n7472), .A2(n805), .B1(n14836), .B2(n806), .ZN(n12811)
         );
  OAI22_X1 U5433 ( .A1(n7456), .A2(n805), .B1(n14796), .B2(n806), .ZN(n12812)
         );
  OAI22_X1 U5434 ( .A1(n7440), .A2(n805), .B1(n14756), .B2(n806), .ZN(n12813)
         );
  OAI22_X1 U5435 ( .A1(n7424), .A2(n805), .B1(n14716), .B2(n806), .ZN(n12814)
         );
  OAI22_X1 U5436 ( .A1(n7408), .A2(n805), .B1(n14676), .B2(n806), .ZN(n12815)
         );
  OAI22_X1 U5437 ( .A1(n7392), .A2(n807), .B1(n14933), .B2(n808), .ZN(n12816)
         );
  OAI22_X1 U5438 ( .A1(n7376), .A2(n807), .B1(n14916), .B2(n808), .ZN(n12817)
         );
  OAI22_X1 U5439 ( .A1(n7360), .A2(n807), .B1(n14876), .B2(n808), .ZN(n12818)
         );
  OAI22_X1 U5440 ( .A1(n7344), .A2(n807), .B1(n14836), .B2(n808), .ZN(n12819)
         );
  OAI22_X1 U5441 ( .A1(n7328), .A2(n807), .B1(n14796), .B2(n808), .ZN(n12820)
         );
  OAI22_X1 U5442 ( .A1(n7312), .A2(n807), .B1(n14756), .B2(n808), .ZN(n12821)
         );
  OAI22_X1 U5443 ( .A1(n7296), .A2(n807), .B1(n14716), .B2(n808), .ZN(n12822)
         );
  OAI22_X1 U5444 ( .A1(n7280), .A2(n807), .B1(n14676), .B2(n808), .ZN(n12823)
         );
  OAI22_X1 U5445 ( .A1(n7264), .A2(n809), .B1(n14933), .B2(n810), .ZN(n12824)
         );
  OAI22_X1 U5446 ( .A1(n7248), .A2(n809), .B1(n14916), .B2(n810), .ZN(n12825)
         );
  OAI22_X1 U5447 ( .A1(n7232), .A2(n809), .B1(n14876), .B2(n810), .ZN(n12826)
         );
  OAI22_X1 U5448 ( .A1(n7216), .A2(n809), .B1(n14836), .B2(n810), .ZN(n12827)
         );
  OAI22_X1 U5449 ( .A1(n7200), .A2(n809), .B1(n14796), .B2(n810), .ZN(n12828)
         );
  OAI22_X1 U5450 ( .A1(n7184), .A2(n809), .B1(n14756), .B2(n810), .ZN(n12829)
         );
  OAI22_X1 U5451 ( .A1(n7168), .A2(n809), .B1(n14716), .B2(n810), .ZN(n12830)
         );
  OAI22_X1 U5452 ( .A1(n7152), .A2(n809), .B1(n14676), .B2(n810), .ZN(n12831)
         );
  OAI22_X1 U5453 ( .A1(n7136), .A2(n811), .B1(n14933), .B2(n812), .ZN(n12832)
         );
  OAI22_X1 U5454 ( .A1(n7120), .A2(n811), .B1(n14916), .B2(n812), .ZN(n12833)
         );
  OAI22_X1 U5455 ( .A1(n7104), .A2(n811), .B1(n14876), .B2(n812), .ZN(n12834)
         );
  OAI22_X1 U5456 ( .A1(n7088), .A2(n811), .B1(n14836), .B2(n812), .ZN(n12835)
         );
  OAI22_X1 U5457 ( .A1(n7072), .A2(n811), .B1(n14796), .B2(n812), .ZN(n12836)
         );
  OAI22_X1 U5458 ( .A1(n7056), .A2(n811), .B1(n14756), .B2(n812), .ZN(n12837)
         );
  OAI22_X1 U5459 ( .A1(n7040), .A2(n811), .B1(n14716), .B2(n812), .ZN(n12838)
         );
  OAI22_X1 U5460 ( .A1(n7024), .A2(n811), .B1(n14676), .B2(n812), .ZN(n12839)
         );
  OAI22_X1 U5461 ( .A1(n7008), .A2(n813), .B1(n14933), .B2(n814), .ZN(n12840)
         );
  OAI22_X1 U5462 ( .A1(n6992), .A2(n813), .B1(n14916), .B2(n814), .ZN(n12841)
         );
  OAI22_X1 U5463 ( .A1(n6976), .A2(n813), .B1(n14876), .B2(n814), .ZN(n12842)
         );
  OAI22_X1 U5464 ( .A1(n6960), .A2(n813), .B1(n14836), .B2(n814), .ZN(n12843)
         );
  OAI22_X1 U5465 ( .A1(n6944), .A2(n813), .B1(n14796), .B2(n814), .ZN(n12844)
         );
  OAI22_X1 U5466 ( .A1(n6928), .A2(n813), .B1(n14756), .B2(n814), .ZN(n12845)
         );
  OAI22_X1 U5467 ( .A1(n6912), .A2(n813), .B1(n14716), .B2(n814), .ZN(n12846)
         );
  OAI22_X1 U5468 ( .A1(n6896), .A2(n813), .B1(n14676), .B2(n814), .ZN(n12847)
         );
  OAI22_X1 U5469 ( .A1(n6880), .A2(n815), .B1(n14933), .B2(n816), .ZN(n12848)
         );
  OAI22_X1 U5470 ( .A1(n6864), .A2(n815), .B1(n14916), .B2(n816), .ZN(n12849)
         );
  OAI22_X1 U5471 ( .A1(n6848), .A2(n815), .B1(n14876), .B2(n816), .ZN(n12850)
         );
  OAI22_X1 U5472 ( .A1(n6832), .A2(n815), .B1(n14836), .B2(n816), .ZN(n12851)
         );
  OAI22_X1 U5473 ( .A1(n6816), .A2(n815), .B1(n14796), .B2(n816), .ZN(n12852)
         );
  OAI22_X1 U5474 ( .A1(n6800), .A2(n815), .B1(n14756), .B2(n816), .ZN(n12853)
         );
  OAI22_X1 U5475 ( .A1(n6784), .A2(n815), .B1(n14716), .B2(n816), .ZN(n12854)
         );
  OAI22_X1 U5476 ( .A1(n6768), .A2(n815), .B1(n14676), .B2(n816), .ZN(n12855)
         );
  OAI22_X1 U5477 ( .A1(n10084), .A2(n829), .B1(n14932), .B2(n830), .ZN(n12904)
         );
  OAI22_X1 U5478 ( .A1(n10068), .A2(n829), .B1(n14917), .B2(n830), .ZN(n12905)
         );
  OAI22_X1 U5479 ( .A1(n10052), .A2(n829), .B1(n14877), .B2(n830), .ZN(n12906)
         );
  OAI22_X1 U5480 ( .A1(n10036), .A2(n829), .B1(n14837), .B2(n830), .ZN(n12907)
         );
  OAI22_X1 U5481 ( .A1(n10020), .A2(n829), .B1(n14797), .B2(n830), .ZN(n12908)
         );
  OAI22_X1 U5482 ( .A1(n10004), .A2(n829), .B1(n14757), .B2(n830), .ZN(n12909)
         );
  OAI22_X1 U5483 ( .A1(n9988), .A2(n829), .B1(n14717), .B2(n830), .ZN(n12910)
         );
  OAI22_X1 U5484 ( .A1(n9972), .A2(n829), .B1(n14677), .B2(n830), .ZN(n12911)
         );
  OAI22_X1 U5485 ( .A1(n9956), .A2(n832), .B1(n14932), .B2(n833), .ZN(n12912)
         );
  OAI22_X1 U5486 ( .A1(n9940), .A2(n832), .B1(n14917), .B2(n833), .ZN(n12913)
         );
  OAI22_X1 U5487 ( .A1(n9924), .A2(n832), .B1(n14877), .B2(n833), .ZN(n12914)
         );
  OAI22_X1 U5489 ( .A1(n9908), .A2(n832), .B1(n14837), .B2(n833), .ZN(n12915)
         );
  OAI22_X1 U5490 ( .A1(n9892), .A2(n832), .B1(n14797), .B2(n833), .ZN(n12916)
         );
  OAI22_X1 U5491 ( .A1(n9876), .A2(n832), .B1(n14757), .B2(n833), .ZN(n12917)
         );
  OAI22_X1 U5492 ( .A1(n9860), .A2(n832), .B1(n14717), .B2(n833), .ZN(n12918)
         );
  OAI22_X1 U5493 ( .A1(n9844), .A2(n832), .B1(n14677), .B2(n833), .ZN(n12919)
         );
  OAI22_X1 U5494 ( .A1(n9828), .A2(n834), .B1(n14932), .B2(n835), .ZN(n12920)
         );
  OAI22_X1 U5495 ( .A1(n9812), .A2(n834), .B1(n14917), .B2(n835), .ZN(n12921)
         );
  OAI22_X1 U5496 ( .A1(n9796), .A2(n834), .B1(n14877), .B2(n835), .ZN(n12922)
         );
  OAI22_X1 U5497 ( .A1(n9780), .A2(n834), .B1(n14837), .B2(n835), .ZN(n12923)
         );
  OAI22_X1 U5498 ( .A1(n9764), .A2(n834), .B1(n14797), .B2(n835), .ZN(n12924)
         );
  OAI22_X1 U5499 ( .A1(n9748), .A2(n834), .B1(n14757), .B2(n835), .ZN(n12925)
         );
  OAI22_X1 U5500 ( .A1(n9732), .A2(n834), .B1(n14717), .B2(n835), .ZN(n12926)
         );
  OAI22_X1 U5501 ( .A1(n9716), .A2(n834), .B1(n14677), .B2(n835), .ZN(n12927)
         );
  OAI22_X1 U5502 ( .A1(n9700), .A2(n836), .B1(n14932), .B2(n837), .ZN(n12928)
         );
  OAI22_X1 U5503 ( .A1(n9684), .A2(n836), .B1(n14917), .B2(n837), .ZN(n12929)
         );
  OAI22_X1 U5504 ( .A1(n9668), .A2(n836), .B1(n14877), .B2(n837), .ZN(n12930)
         );
  OAI22_X1 U5505 ( .A1(n9652), .A2(n836), .B1(n14837), .B2(n837), .ZN(n12931)
         );
  OAI22_X1 U5506 ( .A1(n9636), .A2(n836), .B1(n14797), .B2(n837), .ZN(n12932)
         );
  OAI22_X1 U5507 ( .A1(n9620), .A2(n836), .B1(n14757), .B2(n837), .ZN(n12933)
         );
  OAI22_X1 U5508 ( .A1(n9604), .A2(n836), .B1(n14717), .B2(n837), .ZN(n12934)
         );
  OAI22_X1 U5509 ( .A1(n9588), .A2(n836), .B1(n14677), .B2(n837), .ZN(n12935)
         );
  OAI22_X1 U5510 ( .A1(n9572), .A2(n838), .B1(n14932), .B2(n839), .ZN(n12936)
         );
  OAI22_X1 U5511 ( .A1(n9556), .A2(n838), .B1(n14917), .B2(n839), .ZN(n12937)
         );
  OAI22_X1 U5512 ( .A1(n9540), .A2(n838), .B1(n14877), .B2(n839), .ZN(n12938)
         );
  OAI22_X1 U5513 ( .A1(n9524), .A2(n838), .B1(n14837), .B2(n839), .ZN(n12939)
         );
  OAI22_X1 U5514 ( .A1(n9508), .A2(n838), .B1(n14797), .B2(n839), .ZN(n12940)
         );
  OAI22_X1 U5515 ( .A1(n9492), .A2(n838), .B1(n14757), .B2(n839), .ZN(n12941)
         );
  OAI22_X1 U5516 ( .A1(n9476), .A2(n838), .B1(n14717), .B2(n839), .ZN(n12942)
         );
  OAI22_X1 U5517 ( .A1(n9460), .A2(n838), .B1(n14677), .B2(n839), .ZN(n12943)
         );
  OAI22_X1 U5518 ( .A1(n9444), .A2(n840), .B1(n14932), .B2(n841), .ZN(n12944)
         );
  OAI22_X1 U5519 ( .A1(n9428), .A2(n840), .B1(n14917), .B2(n841), .ZN(n12945)
         );
  OAI22_X1 U5520 ( .A1(n9412), .A2(n840), .B1(n14877), .B2(n841), .ZN(n12946)
         );
  OAI22_X1 U5521 ( .A1(n9396), .A2(n840), .B1(n14837), .B2(n841), .ZN(n12947)
         );
  OAI22_X1 U5522 ( .A1(n9380), .A2(n840), .B1(n14797), .B2(n841), .ZN(n12948)
         );
  OAI22_X1 U5523 ( .A1(n9364), .A2(n840), .B1(n14757), .B2(n841), .ZN(n12949)
         );
  OAI22_X1 U5524 ( .A1(n9348), .A2(n840), .B1(n14717), .B2(n841), .ZN(n12950)
         );
  OAI22_X1 U5525 ( .A1(n9332), .A2(n840), .B1(n14677), .B2(n841), .ZN(n12951)
         );
  OAI22_X1 U5526 ( .A1(n9316), .A2(n842), .B1(n14932), .B2(n843), .ZN(n12952)
         );
  OAI22_X1 U5527 ( .A1(n9300), .A2(n842), .B1(n14917), .B2(n843), .ZN(n12953)
         );
  OAI22_X1 U5528 ( .A1(n9284), .A2(n842), .B1(n14877), .B2(n843), .ZN(n12954)
         );
  OAI22_X1 U5529 ( .A1(n9268), .A2(n842), .B1(n14837), .B2(n843), .ZN(n12955)
         );
  OAI22_X1 U5530 ( .A1(n9252), .A2(n842), .B1(n14797), .B2(n843), .ZN(n12956)
         );
  OAI22_X1 U5531 ( .A1(n9236), .A2(n842), .B1(n14757), .B2(n843), .ZN(n12957)
         );
  OAI22_X1 U5532 ( .A1(n9220), .A2(n842), .B1(n14717), .B2(n843), .ZN(n12958)
         );
  OAI22_X1 U5533 ( .A1(n9204), .A2(n842), .B1(n14677), .B2(n843), .ZN(n12959)
         );
  OAI22_X1 U5534 ( .A1(n9188), .A2(n844), .B1(n14931), .B2(n845), .ZN(n12960)
         );
  OAI22_X1 U5535 ( .A1(n9172), .A2(n844), .B1(n14917), .B2(n845), .ZN(n12961)
         );
  OAI22_X1 U5536 ( .A1(n9156), .A2(n844), .B1(n14877), .B2(n845), .ZN(n12962)
         );
  OAI22_X1 U5537 ( .A1(n9140), .A2(n844), .B1(n14837), .B2(n845), .ZN(n12963)
         );
  OAI22_X1 U5538 ( .A1(n9124), .A2(n844), .B1(n14797), .B2(n845), .ZN(n12964)
         );
  OAI22_X1 U5539 ( .A1(n9108), .A2(n844), .B1(n14757), .B2(n845), .ZN(n12965)
         );
  OAI22_X1 U5540 ( .A1(n9092), .A2(n844), .B1(n14717), .B2(n845), .ZN(n12966)
         );
  OAI22_X1 U5541 ( .A1(n9076), .A2(n844), .B1(n14677), .B2(n845), .ZN(n12967)
         );
  OAI22_X1 U5542 ( .A1(n9060), .A2(n846), .B1(n14931), .B2(n847), .ZN(n12968)
         );
  OAI22_X1 U5543 ( .A1(n9044), .A2(n846), .B1(n14917), .B2(n847), .ZN(n12969)
         );
  OAI22_X1 U5544 ( .A1(n9028), .A2(n846), .B1(n14877), .B2(n847), .ZN(n12970)
         );
  OAI22_X1 U5545 ( .A1(n9012), .A2(n846), .B1(n14837), .B2(n847), .ZN(n12971)
         );
  OAI22_X1 U5546 ( .A1(n8996), .A2(n846), .B1(n14797), .B2(n847), .ZN(n12972)
         );
  OAI22_X1 U5547 ( .A1(n8980), .A2(n846), .B1(n14757), .B2(n847), .ZN(n12973)
         );
  OAI22_X1 U5548 ( .A1(n8964), .A2(n846), .B1(n14717), .B2(n847), .ZN(n12974)
         );
  OAI22_X1 U5549 ( .A1(n8948), .A2(n846), .B1(n14677), .B2(n847), .ZN(n12975)
         );
  OAI22_X1 U5550 ( .A1(n8932), .A2(n848), .B1(n14931), .B2(n849), .ZN(n12976)
         );
  OAI22_X1 U5551 ( .A1(n8916), .A2(n848), .B1(n14917), .B2(n849), .ZN(n12977)
         );
  OAI22_X1 U5552 ( .A1(n8900), .A2(n848), .B1(n14877), .B2(n849), .ZN(n12978)
         );
  OAI22_X1 U5553 ( .A1(n8884), .A2(n848), .B1(n14837), .B2(n849), .ZN(n12979)
         );
  OAI22_X1 U5554 ( .A1(n8868), .A2(n848), .B1(n14797), .B2(n849), .ZN(n12980)
         );
  OAI22_X1 U5555 ( .A1(n8852), .A2(n848), .B1(n14757), .B2(n849), .ZN(n12981)
         );
  OAI22_X1 U5556 ( .A1(n8836), .A2(n848), .B1(n14717), .B2(n849), .ZN(n12982)
         );
  OAI22_X1 U5557 ( .A1(n8820), .A2(n848), .B1(n14677), .B2(n849), .ZN(n12983)
         );
  OAI22_X1 U5558 ( .A1(n8804), .A2(n850), .B1(n14931), .B2(n851), .ZN(n12984)
         );
  OAI22_X1 U5559 ( .A1(n8788), .A2(n850), .B1(n14917), .B2(n851), .ZN(n12985)
         );
  OAI22_X1 U5560 ( .A1(n8772), .A2(n850), .B1(n14877), .B2(n851), .ZN(n12986)
         );
  OAI22_X1 U5561 ( .A1(n8756), .A2(n850), .B1(n14837), .B2(n851), .ZN(n12987)
         );
  OAI22_X1 U5562 ( .A1(n8740), .A2(n850), .B1(n14797), .B2(n851), .ZN(n12988)
         );
  OAI22_X1 U5563 ( .A1(n8724), .A2(n850), .B1(n14757), .B2(n851), .ZN(n12989)
         );
  OAI22_X1 U5564 ( .A1(n8708), .A2(n850), .B1(n14717), .B2(n851), .ZN(n12990)
         );
  OAI22_X1 U5565 ( .A1(n8692), .A2(n850), .B1(n14677), .B2(n851), .ZN(n12991)
         );
  OAI22_X1 U5566 ( .A1(n8676), .A2(n852), .B1(n14931), .B2(n853), .ZN(n12992)
         );
  OAI22_X1 U5567 ( .A1(n8660), .A2(n852), .B1(n14917), .B2(n853), .ZN(n12993)
         );
  OAI22_X1 U5568 ( .A1(n8644), .A2(n852), .B1(n14877), .B2(n853), .ZN(n12994)
         );
  OAI22_X1 U5569 ( .A1(n8628), .A2(n852), .B1(n14837), .B2(n853), .ZN(n12995)
         );
  OAI22_X1 U5570 ( .A1(n8612), .A2(n852), .B1(n14797), .B2(n853), .ZN(n12996)
         );
  OAI22_X1 U5571 ( .A1(n8596), .A2(n852), .B1(n14757), .B2(n853), .ZN(n12997)
         );
  OAI22_X1 U5572 ( .A1(n8580), .A2(n852), .B1(n14717), .B2(n853), .ZN(n12998)
         );
  OAI22_X1 U5573 ( .A1(n8564), .A2(n852), .B1(n14677), .B2(n853), .ZN(n12999)
         );
  OAI22_X1 U5574 ( .A1(n8548), .A2(n854), .B1(n14931), .B2(n855), .ZN(n13000)
         );
  OAI22_X1 U5575 ( .A1(n8532), .A2(n854), .B1(n14918), .B2(n855), .ZN(n13001)
         );
  OAI22_X1 U5576 ( .A1(n8516), .A2(n854), .B1(n14878), .B2(n855), .ZN(n13002)
         );
  OAI22_X1 U5577 ( .A1(n8500), .A2(n854), .B1(n14838), .B2(n855), .ZN(n13003)
         );
  OAI22_X1 U5578 ( .A1(n8484), .A2(n854), .B1(n14798), .B2(n855), .ZN(n13004)
         );
  OAI22_X1 U5579 ( .A1(n8468), .A2(n854), .B1(n14758), .B2(n855), .ZN(n13005)
         );
  OAI22_X1 U5580 ( .A1(n8452), .A2(n854), .B1(n14718), .B2(n855), .ZN(n13006)
         );
  OAI22_X1 U5581 ( .A1(n8436), .A2(n854), .B1(n14678), .B2(n855), .ZN(n13007)
         );
  OAI22_X1 U5582 ( .A1(n8420), .A2(n856), .B1(n14931), .B2(n857), .ZN(n13008)
         );
  OAI22_X1 U5583 ( .A1(n8404), .A2(n856), .B1(n14918), .B2(n857), .ZN(n13009)
         );
  OAI22_X1 U5584 ( .A1(n8388), .A2(n856), .B1(n14878), .B2(n857), .ZN(n13010)
         );
  OAI22_X1 U5585 ( .A1(n8372), .A2(n856), .B1(n14838), .B2(n857), .ZN(n13011)
         );
  OAI22_X1 U5586 ( .A1(n8356), .A2(n856), .B1(n14798), .B2(n857), .ZN(n13012)
         );
  OAI22_X1 U5587 ( .A1(n8340), .A2(n856), .B1(n14758), .B2(n857), .ZN(n13013)
         );
  OAI22_X1 U5588 ( .A1(n8324), .A2(n856), .B1(n14718), .B2(n857), .ZN(n13014)
         );
  OAI22_X1 U5589 ( .A1(n8308), .A2(n856), .B1(n14678), .B2(n857), .ZN(n13015)
         );
  OAI22_X1 U5590 ( .A1(n8292), .A2(n858), .B1(n14931), .B2(n859), .ZN(n13016)
         );
  OAI22_X1 U5591 ( .A1(n8276), .A2(n858), .B1(n14918), .B2(n859), .ZN(n13017)
         );
  OAI22_X1 U5592 ( .A1(n8260), .A2(n858), .B1(n14878), .B2(n859), .ZN(n13018)
         );
  OAI22_X1 U5593 ( .A1(n8244), .A2(n858), .B1(n14838), .B2(n859), .ZN(n13019)
         );
  OAI22_X1 U5594 ( .A1(n8228), .A2(n858), .B1(n14798), .B2(n859), .ZN(n13020)
         );
  OAI22_X1 U5595 ( .A1(n8212), .A2(n858), .B1(n14758), .B2(n859), .ZN(n13021)
         );
  OAI22_X1 U5596 ( .A1(n8196), .A2(n858), .B1(n14718), .B2(n859), .ZN(n13022)
         );
  OAI22_X1 U5597 ( .A1(n8180), .A2(n858), .B1(n14678), .B2(n859), .ZN(n13023)
         );
  OAI22_X1 U5598 ( .A1(n8164), .A2(n860), .B1(n14931), .B2(n861), .ZN(n13024)
         );
  OAI22_X1 U5599 ( .A1(n8148), .A2(n860), .B1(n14918), .B2(n861), .ZN(n13025)
         );
  OAI22_X1 U5600 ( .A1(n8132), .A2(n860), .B1(n14878), .B2(n861), .ZN(n13026)
         );
  OAI22_X1 U5601 ( .A1(n8116), .A2(n860), .B1(n14838), .B2(n861), .ZN(n13027)
         );
  OAI22_X1 U5602 ( .A1(n8100), .A2(n860), .B1(n14798), .B2(n861), .ZN(n13028)
         );
  OAI22_X1 U5603 ( .A1(n8084), .A2(n860), .B1(n14758), .B2(n861), .ZN(n13029)
         );
  OAI22_X1 U5604 ( .A1(n8068), .A2(n860), .B1(n14718), .B2(n861), .ZN(n13030)
         );
  OAI22_X1 U5605 ( .A1(n8052), .A2(n860), .B1(n14678), .B2(n861), .ZN(n13031)
         );
  OAI22_X1 U5606 ( .A1(n8036), .A2(n862), .B1(n14931), .B2(n863), .ZN(n13032)
         );
  OAI22_X1 U5607 ( .A1(n8020), .A2(n862), .B1(n14918), .B2(n863), .ZN(n13033)
         );
  OAI22_X1 U5608 ( .A1(n8004), .A2(n862), .B1(n14878), .B2(n863), .ZN(n13034)
         );
  OAI22_X1 U5609 ( .A1(n7988), .A2(n862), .B1(n14838), .B2(n863), .ZN(n13035)
         );
  OAI22_X1 U5610 ( .A1(n7972), .A2(n862), .B1(n14798), .B2(n863), .ZN(n13036)
         );
  OAI22_X1 U5611 ( .A1(n7956), .A2(n862), .B1(n14758), .B2(n863), .ZN(n13037)
         );
  OAI22_X1 U5612 ( .A1(n7940), .A2(n862), .B1(n14718), .B2(n863), .ZN(n13038)
         );
  OAI22_X1 U5613 ( .A1(n7924), .A2(n862), .B1(n14678), .B2(n863), .ZN(n13039)
         );
  OAI22_X1 U5614 ( .A1(n7908), .A2(n864), .B1(n14931), .B2(n865), .ZN(n13040)
         );
  OAI22_X1 U5615 ( .A1(n7892), .A2(n864), .B1(n14918), .B2(n865), .ZN(n13041)
         );
  OAI22_X1 U5616 ( .A1(n7876), .A2(n864), .B1(n14878), .B2(n865), .ZN(n13042)
         );
  OAI22_X1 U5617 ( .A1(n7860), .A2(n864), .B1(n14838), .B2(n865), .ZN(n13043)
         );
  OAI22_X1 U5618 ( .A1(n7844), .A2(n864), .B1(n14798), .B2(n865), .ZN(n13044)
         );
  OAI22_X1 U5619 ( .A1(n7828), .A2(n864), .B1(n14758), .B2(n865), .ZN(n13045)
         );
  OAI22_X1 U5620 ( .A1(n7812), .A2(n864), .B1(n14718), .B2(n865), .ZN(n13046)
         );
  OAI22_X1 U5621 ( .A1(n7796), .A2(n864), .B1(n14678), .B2(n865), .ZN(n13047)
         );
  OAI22_X1 U5622 ( .A1(n7780), .A2(n866), .B1(n14931), .B2(n867), .ZN(n13048)
         );
  OAI22_X1 U5623 ( .A1(n7764), .A2(n866), .B1(n14918), .B2(n867), .ZN(n13049)
         );
  OAI22_X1 U5624 ( .A1(n7748), .A2(n866), .B1(n14878), .B2(n867), .ZN(n13050)
         );
  OAI22_X1 U5625 ( .A1(n7732), .A2(n866), .B1(n14838), .B2(n867), .ZN(n13051)
         );
  OAI22_X1 U5626 ( .A1(n7716), .A2(n866), .B1(n14798), .B2(n867), .ZN(n13052)
         );
  OAI22_X1 U5627 ( .A1(n7700), .A2(n866), .B1(n14758), .B2(n867), .ZN(n13053)
         );
  OAI22_X1 U5628 ( .A1(n7684), .A2(n866), .B1(n14718), .B2(n867), .ZN(n13054)
         );
  OAI22_X1 U5629 ( .A1(n7668), .A2(n866), .B1(n14678), .B2(n867), .ZN(n13055)
         );
  OAI22_X1 U5630 ( .A1(n7652), .A2(n868), .B1(n14931), .B2(n869), .ZN(n13056)
         );
  OAI22_X1 U5631 ( .A1(n7636), .A2(n868), .B1(n14918), .B2(n869), .ZN(n13057)
         );
  OAI22_X1 U5632 ( .A1(n7620), .A2(n868), .B1(n14878), .B2(n869), .ZN(n13058)
         );
  OAI22_X1 U5633 ( .A1(n7604), .A2(n868), .B1(n14838), .B2(n869), .ZN(n13059)
         );
  OAI22_X1 U5634 ( .A1(n7588), .A2(n868), .B1(n14798), .B2(n869), .ZN(n13060)
         );
  OAI22_X1 U5635 ( .A1(n7572), .A2(n868), .B1(n14758), .B2(n869), .ZN(n13061)
         );
  OAI22_X1 U5636 ( .A1(n7556), .A2(n868), .B1(n14718), .B2(n869), .ZN(n13062)
         );
  OAI22_X1 U5637 ( .A1(n7540), .A2(n868), .B1(n14678), .B2(n869), .ZN(n13063)
         );
  OAI22_X1 U5638 ( .A1(n7524), .A2(n870), .B1(n14930), .B2(n871), .ZN(n13064)
         );
  OAI22_X1 U5639 ( .A1(n7508), .A2(n870), .B1(n14918), .B2(n871), .ZN(n13065)
         );
  OAI22_X1 U5641 ( .A1(n7492), .A2(n870), .B1(n14878), .B2(n871), .ZN(n13066)
         );
  OAI22_X1 U5642 ( .A1(n7476), .A2(n870), .B1(n14838), .B2(n871), .ZN(n13067)
         );
  OAI22_X1 U5643 ( .A1(n7460), .A2(n870), .B1(n14798), .B2(n871), .ZN(n13068)
         );
  OAI22_X1 U5644 ( .A1(n7444), .A2(n870), .B1(n14758), .B2(n871), .ZN(n13069)
         );
  OAI22_X1 U5645 ( .A1(n7428), .A2(n870), .B1(n14718), .B2(n871), .ZN(n13070)
         );
  OAI22_X1 U5646 ( .A1(n7412), .A2(n870), .B1(n14678), .B2(n871), .ZN(n13071)
         );
  OAI22_X1 U5647 ( .A1(n7396), .A2(n872), .B1(n14930), .B2(n873), .ZN(n13072)
         );
  OAI22_X1 U5648 ( .A1(n7380), .A2(n872), .B1(n14918), .B2(n873), .ZN(n13073)
         );
  OAI22_X1 U5649 ( .A1(n7364), .A2(n872), .B1(n14878), .B2(n873), .ZN(n13074)
         );
  OAI22_X1 U5650 ( .A1(n7348), .A2(n872), .B1(n14838), .B2(n873), .ZN(n13075)
         );
  OAI22_X1 U5651 ( .A1(n7332), .A2(n872), .B1(n14798), .B2(n873), .ZN(n13076)
         );
  OAI22_X1 U5652 ( .A1(n7316), .A2(n872), .B1(n14758), .B2(n873), .ZN(n13077)
         );
  OAI22_X1 U5653 ( .A1(n7300), .A2(n872), .B1(n14718), .B2(n873), .ZN(n13078)
         );
  OAI22_X1 U5654 ( .A1(n7284), .A2(n872), .B1(n14678), .B2(n873), .ZN(n13079)
         );
  OAI22_X1 U5655 ( .A1(n7268), .A2(n874), .B1(n14930), .B2(n875), .ZN(n13080)
         );
  OAI22_X1 U5656 ( .A1(n7252), .A2(n874), .B1(n14918), .B2(n875), .ZN(n13081)
         );
  OAI22_X1 U5657 ( .A1(n7236), .A2(n874), .B1(n14878), .B2(n875), .ZN(n13082)
         );
  OAI22_X1 U5658 ( .A1(n7220), .A2(n874), .B1(n14838), .B2(n875), .ZN(n13083)
         );
  OAI22_X1 U5659 ( .A1(n7204), .A2(n874), .B1(n14798), .B2(n875), .ZN(n13084)
         );
  OAI22_X1 U5660 ( .A1(n7188), .A2(n874), .B1(n14758), .B2(n875), .ZN(n13085)
         );
  OAI22_X1 U5661 ( .A1(n7172), .A2(n874), .B1(n14718), .B2(n875), .ZN(n13086)
         );
  OAI22_X1 U5662 ( .A1(n7156), .A2(n874), .B1(n14678), .B2(n875), .ZN(n13087)
         );
  OAI22_X1 U5663 ( .A1(n7140), .A2(n876), .B1(n14930), .B2(n877), .ZN(n13088)
         );
  OAI22_X1 U5664 ( .A1(n7124), .A2(n876), .B1(n14918), .B2(n877), .ZN(n13089)
         );
  OAI22_X1 U5665 ( .A1(n7108), .A2(n876), .B1(n14878), .B2(n877), .ZN(n13090)
         );
  OAI22_X1 U5666 ( .A1(n7092), .A2(n876), .B1(n14838), .B2(n877), .ZN(n13091)
         );
  OAI22_X1 U5667 ( .A1(n7076), .A2(n876), .B1(n14798), .B2(n877), .ZN(n13092)
         );
  OAI22_X1 U5668 ( .A1(n7060), .A2(n876), .B1(n14758), .B2(n877), .ZN(n13093)
         );
  OAI22_X1 U5669 ( .A1(n7044), .A2(n876), .B1(n14718), .B2(n877), .ZN(n13094)
         );
  OAI22_X1 U5670 ( .A1(n7028), .A2(n876), .B1(n14678), .B2(n877), .ZN(n13095)
         );
  OAI22_X1 U5671 ( .A1(n7012), .A2(n878), .B1(n14930), .B2(n879), .ZN(n13096)
         );
  OAI22_X1 U5672 ( .A1(n6996), .A2(n878), .B1(n14918), .B2(n879), .ZN(n13097)
         );
  OAI22_X1 U5673 ( .A1(n6980), .A2(n878), .B1(n14878), .B2(n879), .ZN(n13098)
         );
  OAI22_X1 U5674 ( .A1(n6964), .A2(n878), .B1(n14838), .B2(n879), .ZN(n13099)
         );
  OAI22_X1 U5675 ( .A1(n6948), .A2(n878), .B1(n14798), .B2(n879), .ZN(n13100)
         );
  OAI22_X1 U5676 ( .A1(n6932), .A2(n878), .B1(n14758), .B2(n879), .ZN(n13101)
         );
  OAI22_X1 U5677 ( .A1(n6916), .A2(n878), .B1(n14718), .B2(n879), .ZN(n13102)
         );
  OAI22_X1 U5678 ( .A1(n6900), .A2(n878), .B1(n14678), .B2(n879), .ZN(n13103)
         );
  OAI22_X1 U5679 ( .A1(n6884), .A2(n880), .B1(n14930), .B2(n881), .ZN(n13104)
         );
  OAI22_X1 U5680 ( .A1(n6868), .A2(n880), .B1(n14919), .B2(n881), .ZN(n13105)
         );
  OAI22_X1 U5681 ( .A1(n6852), .A2(n880), .B1(n14879), .B2(n881), .ZN(n13106)
         );
  OAI22_X1 U5682 ( .A1(n6836), .A2(n880), .B1(n14839), .B2(n881), .ZN(n13107)
         );
  OAI22_X1 U5683 ( .A1(n6820), .A2(n880), .B1(n14799), .B2(n881), .ZN(n13108)
         );
  OAI22_X1 U5684 ( .A1(n6804), .A2(n880), .B1(n14759), .B2(n881), .ZN(n13109)
         );
  OAI22_X1 U5685 ( .A1(n6788), .A2(n880), .B1(n14719), .B2(n881), .ZN(n13110)
         );
  OAI22_X1 U5686 ( .A1(n6772), .A2(n880), .B1(n14679), .B2(n881), .ZN(n13111)
         );
  OAI22_X1 U5687 ( .A1(n9306), .A2(n907), .B1(n14949), .B2(n908), .ZN(n13208)
         );
  OAI22_X1 U5688 ( .A1(n9290), .A2(n907), .B1(n14920), .B2(n908), .ZN(n13209)
         );
  OAI22_X1 U5689 ( .A1(n9274), .A2(n907), .B1(n14880), .B2(n908), .ZN(n13210)
         );
  OAI22_X1 U5690 ( .A1(n9258), .A2(n907), .B1(n14840), .B2(n908), .ZN(n13211)
         );
  OAI22_X1 U5691 ( .A1(n9242), .A2(n907), .B1(n14800), .B2(n908), .ZN(n13212)
         );
  OAI22_X1 U5692 ( .A1(n9226), .A2(n907), .B1(n14760), .B2(n908), .ZN(n13213)
         );
  OAI22_X1 U5693 ( .A1(n9210), .A2(n907), .B1(n14720), .B2(n908), .ZN(n13214)
         );
  OAI22_X1 U5694 ( .A1(n9194), .A2(n907), .B1(n14680), .B2(n908), .ZN(n13215)
         );
  OAI22_X1 U5695 ( .A1(n9178), .A2(n909), .B1(n14949), .B2(n910), .ZN(n13216)
         );
  OAI22_X1 U5696 ( .A1(n9162), .A2(n909), .B1(n14920), .B2(n910), .ZN(n13217)
         );
  OAI22_X1 U5697 ( .A1(n9146), .A2(n909), .B1(n14880), .B2(n910), .ZN(n13218)
         );
  OAI22_X1 U5698 ( .A1(n9130), .A2(n909), .B1(n14840), .B2(n910), .ZN(n13219)
         );
  OAI22_X1 U5699 ( .A1(n9114), .A2(n909), .B1(n14800), .B2(n910), .ZN(n13220)
         );
  OAI22_X1 U5700 ( .A1(n9098), .A2(n909), .B1(n14760), .B2(n910), .ZN(n13221)
         );
  OAI22_X1 U5701 ( .A1(n9082), .A2(n909), .B1(n14720), .B2(n910), .ZN(n13222)
         );
  OAI22_X1 U5702 ( .A1(n9066), .A2(n909), .B1(n14680), .B2(n910), .ZN(n13223)
         );
  OAI22_X1 U5703 ( .A1(n9050), .A2(n911), .B1(n14949), .B2(n912), .ZN(n13224)
         );
  OAI22_X1 U5704 ( .A1(n9034), .A2(n911), .B1(n14920), .B2(n912), .ZN(n13225)
         );
  OAI22_X1 U5705 ( .A1(n9018), .A2(n911), .B1(n14880), .B2(n912), .ZN(n13226)
         );
  OAI22_X1 U5706 ( .A1(n9002), .A2(n911), .B1(n14840), .B2(n912), .ZN(n13227)
         );
  OAI22_X1 U5707 ( .A1(n8986), .A2(n911), .B1(n14800), .B2(n912), .ZN(n13228)
         );
  OAI22_X1 U5708 ( .A1(n8970), .A2(n911), .B1(n14760), .B2(n912), .ZN(n13229)
         );
  OAI22_X1 U5709 ( .A1(n8954), .A2(n911), .B1(n14720), .B2(n912), .ZN(n13230)
         );
  OAI22_X1 U5710 ( .A1(n8938), .A2(n911), .B1(n14680), .B2(n912), .ZN(n13231)
         );
  OAI22_X1 U5711 ( .A1(n8922), .A2(n913), .B1(n14948), .B2(n914), .ZN(n13232)
         );
  OAI22_X1 U5712 ( .A1(n8906), .A2(n913), .B1(n14920), .B2(n914), .ZN(n13233)
         );
  OAI22_X1 U5713 ( .A1(n8890), .A2(n913), .B1(n14880), .B2(n914), .ZN(n13234)
         );
  OAI22_X1 U5714 ( .A1(n8874), .A2(n913), .B1(n14840), .B2(n914), .ZN(n13235)
         );
  OAI22_X1 U5715 ( .A1(n8858), .A2(n913), .B1(n14800), .B2(n914), .ZN(n13236)
         );
  OAI22_X1 U5716 ( .A1(n8842), .A2(n913), .B1(n14760), .B2(n914), .ZN(n13237)
         );
  OAI22_X1 U5717 ( .A1(n8826), .A2(n913), .B1(n14720), .B2(n914), .ZN(n13238)
         );
  OAI22_X1 U5718 ( .A1(n8810), .A2(n913), .B1(n14680), .B2(n914), .ZN(n13239)
         );
  OAI22_X1 U5719 ( .A1(n8794), .A2(n915), .B1(n14948), .B2(n916), .ZN(n13240)
         );
  OAI22_X1 U5720 ( .A1(n8778), .A2(n915), .B1(n14920), .B2(n916), .ZN(n13241)
         );
  OAI22_X1 U5721 ( .A1(n8762), .A2(n915), .B1(n14880), .B2(n916), .ZN(n13242)
         );
  OAI22_X1 U5722 ( .A1(n8746), .A2(n915), .B1(n14840), .B2(n916), .ZN(n13243)
         );
  OAI22_X1 U5723 ( .A1(n8730), .A2(n915), .B1(n14800), .B2(n916), .ZN(n13244)
         );
  OAI22_X1 U5724 ( .A1(n8714), .A2(n915), .B1(n14760), .B2(n916), .ZN(n13245)
         );
  OAI22_X1 U5725 ( .A1(n8698), .A2(n915), .B1(n14720), .B2(n916), .ZN(n13246)
         );
  OAI22_X1 U5726 ( .A1(n8682), .A2(n915), .B1(n14680), .B2(n916), .ZN(n13247)
         );
  OAI22_X1 U5727 ( .A1(n8666), .A2(n917), .B1(n14948), .B2(n918), .ZN(n13248)
         );
  OAI22_X1 U5728 ( .A1(n8650), .A2(n917), .B1(n14920), .B2(n918), .ZN(n13249)
         );
  OAI22_X1 U5729 ( .A1(n8634), .A2(n917), .B1(n14880), .B2(n918), .ZN(n13250)
         );
  OAI22_X1 U5730 ( .A1(n8618), .A2(n917), .B1(n14840), .B2(n918), .ZN(n13251)
         );
  OAI22_X1 U5731 ( .A1(n8602), .A2(n917), .B1(n14800), .B2(n918), .ZN(n13252)
         );
  OAI22_X1 U5732 ( .A1(n8586), .A2(n917), .B1(n14760), .B2(n918), .ZN(n13253)
         );
  OAI22_X1 U5733 ( .A1(n8570), .A2(n917), .B1(n14720), .B2(n918), .ZN(n13254)
         );
  OAI22_X1 U5734 ( .A1(n8554), .A2(n917), .B1(n14680), .B2(n918), .ZN(n13255)
         );
  OAI22_X1 U5735 ( .A1(n8538), .A2(n919), .B1(n14948), .B2(n920), .ZN(n13256)
         );
  OAI22_X1 U5736 ( .A1(n8522), .A2(n919), .B1(n14920), .B2(n920), .ZN(n13257)
         );
  OAI22_X1 U5737 ( .A1(n8506), .A2(n919), .B1(n14880), .B2(n920), .ZN(n13258)
         );
  OAI22_X1 U5738 ( .A1(n8490), .A2(n919), .B1(n14840), .B2(n920), .ZN(n13259)
         );
  OAI22_X1 U5739 ( .A1(n8474), .A2(n919), .B1(n14800), .B2(n920), .ZN(n13260)
         );
  OAI22_X1 U5740 ( .A1(n8458), .A2(n919), .B1(n14760), .B2(n920), .ZN(n13261)
         );
  OAI22_X1 U5741 ( .A1(n8442), .A2(n919), .B1(n14720), .B2(n920), .ZN(n13262)
         );
  OAI22_X1 U5742 ( .A1(n8426), .A2(n919), .B1(n14680), .B2(n920), .ZN(n13263)
         );
  OAI22_X1 U5743 ( .A1(n8410), .A2(n921), .B1(n14948), .B2(n922), .ZN(n13264)
         );
  OAI22_X1 U5744 ( .A1(n8394), .A2(n921), .B1(n14920), .B2(n922), .ZN(n13265)
         );
  OAI22_X1 U5745 ( .A1(n8378), .A2(n921), .B1(n14880), .B2(n922), .ZN(n13266)
         );
  OAI22_X1 U5746 ( .A1(n8362), .A2(n921), .B1(n14840), .B2(n922), .ZN(n13267)
         );
  OAI22_X1 U5747 ( .A1(n8346), .A2(n921), .B1(n14800), .B2(n922), .ZN(n13268)
         );
  OAI22_X1 U5748 ( .A1(n8330), .A2(n921), .B1(n14760), .B2(n922), .ZN(n13269)
         );
  OAI22_X1 U5749 ( .A1(n8314), .A2(n921), .B1(n14720), .B2(n922), .ZN(n13270)
         );
  OAI22_X1 U5750 ( .A1(n8298), .A2(n921), .B1(n14680), .B2(n922), .ZN(n13271)
         );
  OAI22_X1 U5751 ( .A1(n8282), .A2(n923), .B1(n14948), .B2(n924), .ZN(n13272)
         );
  OAI22_X1 U5752 ( .A1(n8266), .A2(n923), .B1(n14920), .B2(n924), .ZN(n13273)
         );
  OAI22_X1 U5753 ( .A1(n8250), .A2(n923), .B1(n14880), .B2(n924), .ZN(n13274)
         );
  OAI22_X1 U5754 ( .A1(n8234), .A2(n923), .B1(n14840), .B2(n924), .ZN(n13275)
         );
  OAI22_X1 U5755 ( .A1(n8218), .A2(n923), .B1(n14800), .B2(n924), .ZN(n13276)
         );
  OAI22_X1 U5756 ( .A1(n8202), .A2(n923), .B1(n14760), .B2(n924), .ZN(n13277)
         );
  OAI22_X1 U5757 ( .A1(n8186), .A2(n923), .B1(n14720), .B2(n924), .ZN(n13278)
         );
  OAI22_X1 U5758 ( .A1(n8170), .A2(n923), .B1(n14680), .B2(n924), .ZN(n13279)
         );
  OAI22_X1 U5759 ( .A1(n8154), .A2(n925), .B1(n14948), .B2(n926), .ZN(n13280)
         );
  OAI22_X1 U5760 ( .A1(n8138), .A2(n925), .B1(n14920), .B2(n926), .ZN(n13281)
         );
  OAI22_X1 U5761 ( .A1(n8122), .A2(n925), .B1(n14880), .B2(n926), .ZN(n13282)
         );
  OAI22_X1 U5762 ( .A1(n8106), .A2(n925), .B1(n14840), .B2(n926), .ZN(n13283)
         );
  OAI22_X1 U5763 ( .A1(n8090), .A2(n925), .B1(n14800), .B2(n926), .ZN(n13284)
         );
  OAI22_X1 U5764 ( .A1(n8074), .A2(n925), .B1(n14760), .B2(n926), .ZN(n13285)
         );
  OAI22_X1 U5765 ( .A1(n8058), .A2(n925), .B1(n14720), .B2(n926), .ZN(n13286)
         );
  OAI22_X1 U5766 ( .A1(n8042), .A2(n925), .B1(n14680), .B2(n926), .ZN(n13287)
         );
  OAI22_X1 U5767 ( .A1(n8026), .A2(n927), .B1(n14948), .B2(n928), .ZN(n13288)
         );
  OAI22_X1 U5768 ( .A1(n8010), .A2(n927), .B1(n14920), .B2(n928), .ZN(n13289)
         );
  OAI22_X1 U5769 ( .A1(n7994), .A2(n927), .B1(n14880), .B2(n928), .ZN(n13290)
         );
  OAI22_X1 U5770 ( .A1(n7978), .A2(n927), .B1(n14840), .B2(n928), .ZN(n13291)
         );
  OAI22_X1 U5771 ( .A1(n7962), .A2(n927), .B1(n14800), .B2(n928), .ZN(n13292)
         );
  OAI22_X1 U5772 ( .A1(n7946), .A2(n927), .B1(n14760), .B2(n928), .ZN(n13293)
         );
  OAI22_X1 U5773 ( .A1(n7930), .A2(n927), .B1(n14720), .B2(n928), .ZN(n13294)
         );
  OAI22_X1 U5774 ( .A1(n7914), .A2(n927), .B1(n14680), .B2(n928), .ZN(n13295)
         );
  OAI22_X1 U5775 ( .A1(n7898), .A2(n929), .B1(n14948), .B2(n930), .ZN(n13296)
         );
  OAI22_X1 U5776 ( .A1(n7882), .A2(n929), .B1(n14920), .B2(n930), .ZN(n13297)
         );
  OAI22_X1 U5777 ( .A1(n7866), .A2(n929), .B1(n14880), .B2(n930), .ZN(n13298)
         );
  OAI22_X1 U5778 ( .A1(n7850), .A2(n929), .B1(n14840), .B2(n930), .ZN(n13299)
         );
  OAI22_X1 U5779 ( .A1(n7834), .A2(n929), .B1(n14800), .B2(n930), .ZN(n13300)
         );
  OAI22_X1 U5780 ( .A1(n7818), .A2(n929), .B1(n14760), .B2(n930), .ZN(n13301)
         );
  OAI22_X1 U5781 ( .A1(n7802), .A2(n929), .B1(n14720), .B2(n930), .ZN(n13302)
         );
  OAI22_X1 U5782 ( .A1(n7786), .A2(n929), .B1(n14680), .B2(n930), .ZN(n13303)
         );
  OAI22_X1 U5783 ( .A1(n7770), .A2(n931), .B1(n14948), .B2(n932), .ZN(n13304)
         );
  OAI22_X1 U5784 ( .A1(n7754), .A2(n931), .B1(n14920), .B2(n932), .ZN(n13305)
         );
  OAI22_X1 U5785 ( .A1(n7738), .A2(n931), .B1(n14880), .B2(n932), .ZN(n13306)
         );
  OAI22_X1 U5786 ( .A1(n7722), .A2(n931), .B1(n14840), .B2(n932), .ZN(n13307)
         );
  OAI22_X1 U5787 ( .A1(n7706), .A2(n931), .B1(n14800), .B2(n932), .ZN(n13308)
         );
  OAI22_X1 U5788 ( .A1(n7690), .A2(n931), .B1(n14760), .B2(n932), .ZN(n13309)
         );
  OAI22_X1 U5789 ( .A1(n7674), .A2(n931), .B1(n14720), .B2(n932), .ZN(n13310)
         );
  OAI22_X1 U5790 ( .A1(n7658), .A2(n931), .B1(n14680), .B2(n932), .ZN(n13311)
         );
  OAI22_X1 U5791 ( .A1(n10078), .A2(n960), .B1(n14947), .B2(n961), .ZN(n13416)
         );
  OAI22_X1 U5793 ( .A1(n10062), .A2(n960), .B1(n14922), .B2(n961), .ZN(n13417)
         );
  OAI22_X1 U5794 ( .A1(n10046), .A2(n960), .B1(n14882), .B2(n961), .ZN(n13418)
         );
  OAI22_X1 U5795 ( .A1(n10030), .A2(n960), .B1(n14842), .B2(n961), .ZN(n13419)
         );
  OAI22_X1 U5796 ( .A1(n10014), .A2(n960), .B1(n14802), .B2(n961), .ZN(n13420)
         );
  OAI22_X1 U5797 ( .A1(n9998), .A2(n960), .B1(n14762), .B2(n961), .ZN(n13421)
         );
  OAI22_X1 U5798 ( .A1(n9982), .A2(n960), .B1(n14722), .B2(n961), .ZN(n13422)
         );
  OAI22_X1 U5799 ( .A1(n9966), .A2(n960), .B1(n14682), .B2(n961), .ZN(n13423)
         );
  OAI22_X1 U5800 ( .A1(n9950), .A2(n963), .B1(n14947), .B2(n964), .ZN(n13424)
         );
  OAI22_X1 U5801 ( .A1(n9934), .A2(n963), .B1(n14922), .B2(n964), .ZN(n13425)
         );
  OAI22_X1 U5802 ( .A1(n9918), .A2(n963), .B1(n14882), .B2(n964), .ZN(n13426)
         );
  OAI22_X1 U5803 ( .A1(n9902), .A2(n963), .B1(n14842), .B2(n964), .ZN(n13427)
         );
  OAI22_X1 U5804 ( .A1(n9886), .A2(n963), .B1(n14802), .B2(n964), .ZN(n13428)
         );
  OAI22_X1 U5805 ( .A1(n9870), .A2(n963), .B1(n14762), .B2(n964), .ZN(n13429)
         );
  OAI22_X1 U5806 ( .A1(n9854), .A2(n963), .B1(n14722), .B2(n964), .ZN(n13430)
         );
  OAI22_X1 U5807 ( .A1(n9838), .A2(n963), .B1(n14682), .B2(n964), .ZN(n13431)
         );
  OAI22_X1 U5808 ( .A1(n9822), .A2(n965), .B1(n14947), .B2(n966), .ZN(n13432)
         );
  OAI22_X1 U5809 ( .A1(n9806), .A2(n965), .B1(n14922), .B2(n966), .ZN(n13433)
         );
  OAI22_X1 U5810 ( .A1(n9790), .A2(n965), .B1(n14882), .B2(n966), .ZN(n13434)
         );
  OAI22_X1 U5811 ( .A1(n9774), .A2(n965), .B1(n14842), .B2(n966), .ZN(n13435)
         );
  OAI22_X1 U5812 ( .A1(n9758), .A2(n965), .B1(n14802), .B2(n966), .ZN(n13436)
         );
  OAI22_X1 U5813 ( .A1(n9742), .A2(n965), .B1(n14762), .B2(n966), .ZN(n13437)
         );
  OAI22_X1 U5814 ( .A1(n9726), .A2(n965), .B1(n14722), .B2(n966), .ZN(n13438)
         );
  OAI22_X1 U5815 ( .A1(n9710), .A2(n965), .B1(n14682), .B2(n966), .ZN(n13439)
         );
  OAI22_X1 U5816 ( .A1(n9694), .A2(n967), .B1(n14946), .B2(n968), .ZN(n13440)
         );
  OAI22_X1 U5817 ( .A1(n9678), .A2(n967), .B1(n14922), .B2(n968), .ZN(n13441)
         );
  OAI22_X1 U5818 ( .A1(n9662), .A2(n967), .B1(n14882), .B2(n968), .ZN(n13442)
         );
  OAI22_X1 U5819 ( .A1(n9646), .A2(n967), .B1(n14842), .B2(n968), .ZN(n13443)
         );
  OAI22_X1 U5820 ( .A1(n9630), .A2(n967), .B1(n14802), .B2(n968), .ZN(n13444)
         );
  OAI22_X1 U5821 ( .A1(n9614), .A2(n967), .B1(n14762), .B2(n968), .ZN(n13445)
         );
  OAI22_X1 U5822 ( .A1(n9598), .A2(n967), .B1(n14722), .B2(n968), .ZN(n13446)
         );
  OAI22_X1 U5823 ( .A1(n9582), .A2(n967), .B1(n14682), .B2(n968), .ZN(n13447)
         );
  OAI22_X1 U5824 ( .A1(n9566), .A2(n969), .B1(n14946), .B2(n970), .ZN(n13448)
         );
  OAI22_X1 U5825 ( .A1(n9550), .A2(n969), .B1(n14922), .B2(n970), .ZN(n13449)
         );
  OAI22_X1 U5826 ( .A1(n9534), .A2(n969), .B1(n14882), .B2(n970), .ZN(n13450)
         );
  OAI22_X1 U5827 ( .A1(n9518), .A2(n969), .B1(n14842), .B2(n970), .ZN(n13451)
         );
  OAI22_X1 U5828 ( .A1(n9502), .A2(n969), .B1(n14802), .B2(n970), .ZN(n13452)
         );
  OAI22_X1 U5829 ( .A1(n9486), .A2(n969), .B1(n14762), .B2(n970), .ZN(n13453)
         );
  OAI22_X1 U5830 ( .A1(n9470), .A2(n969), .B1(n14722), .B2(n970), .ZN(n13454)
         );
  OAI22_X1 U5831 ( .A1(n9454), .A2(n969), .B1(n14682), .B2(n970), .ZN(n13455)
         );
  OAI22_X1 U5832 ( .A1(n9438), .A2(n971), .B1(n14946), .B2(n972), .ZN(n13456)
         );
  OAI22_X1 U5833 ( .A1(n9422), .A2(n971), .B1(n14922), .B2(n972), .ZN(n13457)
         );
  OAI22_X1 U5834 ( .A1(n9406), .A2(n971), .B1(n14882), .B2(n972), .ZN(n13458)
         );
  OAI22_X1 U5835 ( .A1(n9390), .A2(n971), .B1(n14842), .B2(n972), .ZN(n13459)
         );
  OAI22_X1 U5836 ( .A1(n9374), .A2(n971), .B1(n14802), .B2(n972), .ZN(n13460)
         );
  OAI22_X1 U5837 ( .A1(n9358), .A2(n971), .B1(n14762), .B2(n972), .ZN(n13461)
         );
  OAI22_X1 U5838 ( .A1(n9342), .A2(n971), .B1(n14722), .B2(n972), .ZN(n13462)
         );
  OAI22_X1 U5839 ( .A1(n9326), .A2(n971), .B1(n14682), .B2(n972), .ZN(n13463)
         );
  OAI22_X1 U5840 ( .A1(n9310), .A2(n973), .B1(n14946), .B2(n974), .ZN(n13464)
         );
  OAI22_X1 U5841 ( .A1(n9294), .A2(n973), .B1(n14922), .B2(n974), .ZN(n13465)
         );
  OAI22_X1 U5842 ( .A1(n9278), .A2(n973), .B1(n14882), .B2(n974), .ZN(n13466)
         );
  OAI22_X1 U5843 ( .A1(n9262), .A2(n973), .B1(n14842), .B2(n974), .ZN(n13467)
         );
  OAI22_X1 U5844 ( .A1(n9246), .A2(n973), .B1(n14802), .B2(n974), .ZN(n13468)
         );
  OAI22_X1 U5845 ( .A1(n9230), .A2(n973), .B1(n14762), .B2(n974), .ZN(n13469)
         );
  OAI22_X1 U5846 ( .A1(n9214), .A2(n973), .B1(n14722), .B2(n974), .ZN(n13470)
         );
  OAI22_X1 U5847 ( .A1(n9198), .A2(n973), .B1(n14682), .B2(n974), .ZN(n13471)
         );
  OAI22_X1 U5848 ( .A1(n9182), .A2(n975), .B1(n14946), .B2(n976), .ZN(n13472)
         );
  OAI22_X1 U5849 ( .A1(n9166), .A2(n975), .B1(n14922), .B2(n976), .ZN(n13473)
         );
  OAI22_X1 U5850 ( .A1(n9150), .A2(n975), .B1(n14882), .B2(n976), .ZN(n13474)
         );
  OAI22_X1 U5851 ( .A1(n9134), .A2(n975), .B1(n14842), .B2(n976), .ZN(n13475)
         );
  OAI22_X1 U5852 ( .A1(n9118), .A2(n975), .B1(n14802), .B2(n976), .ZN(n13476)
         );
  OAI22_X1 U5853 ( .A1(n9102), .A2(n975), .B1(n14762), .B2(n976), .ZN(n13477)
         );
  OAI22_X1 U5854 ( .A1(n9086), .A2(n975), .B1(n14722), .B2(n976), .ZN(n13478)
         );
  OAI22_X1 U5855 ( .A1(n9070), .A2(n975), .B1(n14682), .B2(n976), .ZN(n13479)
         );
  OAI22_X1 U5856 ( .A1(n9054), .A2(n977), .B1(n14946), .B2(n978), .ZN(n13480)
         );
  OAI22_X1 U5857 ( .A1(n9038), .A2(n977), .B1(n14922), .B2(n978), .ZN(n13481)
         );
  OAI22_X1 U5858 ( .A1(n9022), .A2(n977), .B1(n14882), .B2(n978), .ZN(n13482)
         );
  OAI22_X1 U5859 ( .A1(n9006), .A2(n977), .B1(n14842), .B2(n978), .ZN(n13483)
         );
  OAI22_X1 U5860 ( .A1(n8990), .A2(n977), .B1(n14802), .B2(n978), .ZN(n13484)
         );
  OAI22_X1 U5861 ( .A1(n8974), .A2(n977), .B1(n14762), .B2(n978), .ZN(n13485)
         );
  OAI22_X1 U5862 ( .A1(n8958), .A2(n977), .B1(n14722), .B2(n978), .ZN(n13486)
         );
  OAI22_X1 U5863 ( .A1(n8942), .A2(n977), .B1(n14682), .B2(n978), .ZN(n13487)
         );
  OAI22_X1 U5864 ( .A1(n8926), .A2(n979), .B1(n14946), .B2(n980), .ZN(n13488)
         );
  OAI22_X1 U5865 ( .A1(n8910), .A2(n979), .B1(n14922), .B2(n980), .ZN(n13489)
         );
  OAI22_X1 U5866 ( .A1(n8894), .A2(n979), .B1(n14882), .B2(n980), .ZN(n13490)
         );
  OAI22_X1 U5867 ( .A1(n8878), .A2(n979), .B1(n14842), .B2(n980), .ZN(n13491)
         );
  OAI22_X1 U5868 ( .A1(n8862), .A2(n979), .B1(n14802), .B2(n980), .ZN(n13492)
         );
  OAI22_X1 U5869 ( .A1(n8846), .A2(n979), .B1(n14762), .B2(n980), .ZN(n13493)
         );
  OAI22_X1 U5870 ( .A1(n8830), .A2(n979), .B1(n14722), .B2(n980), .ZN(n13494)
         );
  OAI22_X1 U5871 ( .A1(n8814), .A2(n979), .B1(n14682), .B2(n980), .ZN(n13495)
         );
  OAI22_X1 U5872 ( .A1(n8798), .A2(n981), .B1(n14946), .B2(n982), .ZN(n13496)
         );
  OAI22_X1 U5873 ( .A1(n8782), .A2(n981), .B1(n14922), .B2(n982), .ZN(n13497)
         );
  OAI22_X1 U5874 ( .A1(n8766), .A2(n981), .B1(n14882), .B2(n982), .ZN(n13498)
         );
  OAI22_X1 U5875 ( .A1(n8750), .A2(n981), .B1(n14842), .B2(n982), .ZN(n13499)
         );
  OAI22_X1 U5876 ( .A1(n8734), .A2(n981), .B1(n14802), .B2(n982), .ZN(n13500)
         );
  OAI22_X1 U5877 ( .A1(n8718), .A2(n981), .B1(n14762), .B2(n982), .ZN(n13501)
         );
  OAI22_X1 U5878 ( .A1(n8702), .A2(n981), .B1(n14722), .B2(n982), .ZN(n13502)
         );
  OAI22_X1 U5879 ( .A1(n8686), .A2(n981), .B1(n14682), .B2(n982), .ZN(n13503)
         );
  OAI22_X1 U5880 ( .A1(n8670), .A2(n983), .B1(n14946), .B2(n984), .ZN(n13504)
         );
  OAI22_X1 U5881 ( .A1(n8654), .A2(n983), .B1(n14922), .B2(n984), .ZN(n13505)
         );
  OAI22_X1 U5882 ( .A1(n8638), .A2(n983), .B1(n14882), .B2(n984), .ZN(n13506)
         );
  OAI22_X1 U5883 ( .A1(n8622), .A2(n983), .B1(n14842), .B2(n984), .ZN(n13507)
         );
  OAI22_X1 U5884 ( .A1(n8606), .A2(n983), .B1(n14802), .B2(n984), .ZN(n13508)
         );
  OAI22_X1 U5885 ( .A1(n8590), .A2(n983), .B1(n14762), .B2(n984), .ZN(n13509)
         );
  OAI22_X1 U5886 ( .A1(n8574), .A2(n983), .B1(n14722), .B2(n984), .ZN(n13510)
         );
  OAI22_X1 U5887 ( .A1(n8558), .A2(n983), .B1(n14682), .B2(n984), .ZN(n13511)
         );
  OAI22_X1 U5888 ( .A1(n8542), .A2(n985), .B1(n14946), .B2(n986), .ZN(n13512)
         );
  OAI22_X1 U5889 ( .A1(n8526), .A2(n985), .B1(n14922), .B2(n986), .ZN(n13513)
         );
  OAI22_X1 U5890 ( .A1(n8510), .A2(n985), .B1(n14882), .B2(n986), .ZN(n13514)
         );
  OAI22_X1 U5891 ( .A1(n8494), .A2(n985), .B1(n14842), .B2(n986), .ZN(n13515)
         );
  OAI22_X1 U5892 ( .A1(n8478), .A2(n985), .B1(n14802), .B2(n986), .ZN(n13516)
         );
  OAI22_X1 U5893 ( .A1(n8462), .A2(n985), .B1(n14762), .B2(n986), .ZN(n13517)
         );
  OAI22_X1 U5894 ( .A1(n8446), .A2(n985), .B1(n14722), .B2(n986), .ZN(n13518)
         );
  OAI22_X1 U5895 ( .A1(n8430), .A2(n985), .B1(n14682), .B2(n986), .ZN(n13519)
         );
  OAI22_X1 U5896 ( .A1(n8414), .A2(n987), .B1(n14946), .B2(n988), .ZN(n13520)
         );
  OAI22_X1 U5897 ( .A1(n8398), .A2(n987), .B1(n14923), .B2(n988), .ZN(n13521)
         );
  OAI22_X1 U5898 ( .A1(n8382), .A2(n987), .B1(n14883), .B2(n988), .ZN(n13522)
         );
  OAI22_X1 U5899 ( .A1(n8366), .A2(n987), .B1(n14843), .B2(n988), .ZN(n13523)
         );
  OAI22_X1 U5900 ( .A1(n8350), .A2(n987), .B1(n14803), .B2(n988), .ZN(n13524)
         );
  OAI22_X1 U5901 ( .A1(n8334), .A2(n987), .B1(n14763), .B2(n988), .ZN(n13525)
         );
  OAI22_X1 U5902 ( .A1(n8318), .A2(n987), .B1(n14723), .B2(n988), .ZN(n13526)
         );
  OAI22_X1 U5903 ( .A1(n8302), .A2(n987), .B1(n14683), .B2(n988), .ZN(n13527)
         );
  OAI22_X1 U5904 ( .A1(n8286), .A2(n989), .B1(n14946), .B2(n990), .ZN(n13528)
         );
  OAI22_X1 U5905 ( .A1(n8270), .A2(n989), .B1(n14923), .B2(n990), .ZN(n13529)
         );
  OAI22_X1 U5906 ( .A1(n8254), .A2(n989), .B1(n14883), .B2(n990), .ZN(n13530)
         );
  OAI22_X1 U5907 ( .A1(n8238), .A2(n989), .B1(n14843), .B2(n990), .ZN(n13531)
         );
  OAI22_X1 U5908 ( .A1(n8222), .A2(n989), .B1(n14803), .B2(n990), .ZN(n13532)
         );
  OAI22_X1 U5909 ( .A1(n8206), .A2(n989), .B1(n14763), .B2(n990), .ZN(n13533)
         );
  OAI22_X1 U5910 ( .A1(n8190), .A2(n989), .B1(n14723), .B2(n990), .ZN(n13534)
         );
  OAI22_X1 U5911 ( .A1(n8174), .A2(n989), .B1(n14683), .B2(n990), .ZN(n13535)
         );
  OAI22_X1 U5912 ( .A1(n8158), .A2(n991), .B1(n14946), .B2(n992), .ZN(n13536)
         );
  OAI22_X1 U5913 ( .A1(n8142), .A2(n991), .B1(n14923), .B2(n992), .ZN(n13537)
         );
  OAI22_X1 U5914 ( .A1(n8126), .A2(n991), .B1(n14883), .B2(n992), .ZN(n13538)
         );
  OAI22_X1 U5915 ( .A1(n8110), .A2(n991), .B1(n14843), .B2(n992), .ZN(n13539)
         );
  OAI22_X1 U5916 ( .A1(n8094), .A2(n991), .B1(n14803), .B2(n992), .ZN(n13540)
         );
  OAI22_X1 U5917 ( .A1(n8078), .A2(n991), .B1(n14763), .B2(n992), .ZN(n13541)
         );
  OAI22_X1 U5918 ( .A1(n8062), .A2(n991), .B1(n14723), .B2(n992), .ZN(n13542)
         );
  OAI22_X1 U5919 ( .A1(n8046), .A2(n991), .B1(n14683), .B2(n992), .ZN(n13543)
         );
  OAI22_X1 U5920 ( .A1(n8030), .A2(n993), .B1(n14945), .B2(n994), .ZN(n13544)
         );
  OAI22_X1 U5921 ( .A1(n8014), .A2(n993), .B1(n14923), .B2(n994), .ZN(n13545)
         );
  OAI22_X1 U5922 ( .A1(n7998), .A2(n993), .B1(n14883), .B2(n994), .ZN(n13546)
         );
  OAI22_X1 U5923 ( .A1(n7982), .A2(n993), .B1(n14843), .B2(n994), .ZN(n13547)
         );
  OAI22_X1 U5924 ( .A1(n7966), .A2(n993), .B1(n14803), .B2(n994), .ZN(n13548)
         );
  OAI22_X1 U5925 ( .A1(n7950), .A2(n993), .B1(n14763), .B2(n994), .ZN(n13549)
         );
  OAI22_X1 U5926 ( .A1(n7934), .A2(n993), .B1(n14723), .B2(n994), .ZN(n13550)
         );
  OAI22_X1 U5927 ( .A1(n7918), .A2(n993), .B1(n14683), .B2(n994), .ZN(n13551)
         );
  OAI22_X1 U5928 ( .A1(n7902), .A2(n995), .B1(n14945), .B2(n996), .ZN(n13552)
         );
  OAI22_X1 U5929 ( .A1(n7886), .A2(n995), .B1(n14923), .B2(n996), .ZN(n13553)
         );
  OAI22_X1 U5930 ( .A1(n7870), .A2(n995), .B1(n14883), .B2(n996), .ZN(n13554)
         );
  OAI22_X1 U5931 ( .A1(n7854), .A2(n995), .B1(n14843), .B2(n996), .ZN(n13555)
         );
  OAI22_X1 U5932 ( .A1(n7838), .A2(n995), .B1(n14803), .B2(n996), .ZN(n13556)
         );
  OAI22_X1 U5933 ( .A1(n7822), .A2(n995), .B1(n14763), .B2(n996), .ZN(n13557)
         );
  OAI22_X1 U5934 ( .A1(n7806), .A2(n995), .B1(n14723), .B2(n996), .ZN(n13558)
         );
  OAI22_X1 U5935 ( .A1(n7790), .A2(n995), .B1(n14683), .B2(n996), .ZN(n13559)
         );
  OAI22_X1 U5936 ( .A1(n7774), .A2(n997), .B1(n14945), .B2(n998), .ZN(n13560)
         );
  OAI22_X1 U5937 ( .A1(n7758), .A2(n997), .B1(n14923), .B2(n998), .ZN(n13561)
         );
  OAI22_X1 U5938 ( .A1(n7742), .A2(n997), .B1(n14883), .B2(n998), .ZN(n13562)
         );
  OAI22_X1 U5939 ( .A1(n7726), .A2(n997), .B1(n14843), .B2(n998), .ZN(n13563)
         );
  OAI22_X1 U5940 ( .A1(n7710), .A2(n997), .B1(n14803), .B2(n998), .ZN(n13564)
         );
  OAI22_X1 U5941 ( .A1(n7694), .A2(n997), .B1(n14763), .B2(n998), .ZN(n13565)
         );
  OAI22_X1 U5942 ( .A1(n7678), .A2(n997), .B1(n14723), .B2(n998), .ZN(n13566)
         );
  OAI22_X1 U5943 ( .A1(n7662), .A2(n997), .B1(n14683), .B2(n998), .ZN(n13567)
         );
  OAI22_X1 U5945 ( .A1(n7646), .A2(n999), .B1(n14945), .B2(n1000), .ZN(n13568)
         );
  OAI22_X1 U5946 ( .A1(n7630), .A2(n999), .B1(n14923), .B2(n1000), .ZN(n13569)
         );
  OAI22_X1 U5947 ( .A1(n7614), .A2(n999), .B1(n14883), .B2(n1000), .ZN(n13570)
         );
  OAI22_X1 U5948 ( .A1(n7598), .A2(n999), .B1(n14843), .B2(n1000), .ZN(n13571)
         );
  OAI22_X1 U5949 ( .A1(n7582), .A2(n999), .B1(n14803), .B2(n1000), .ZN(n13572)
         );
  OAI22_X1 U5950 ( .A1(n7566), .A2(n999), .B1(n14763), .B2(n1000), .ZN(n13573)
         );
  OAI22_X1 U5951 ( .A1(n7550), .A2(n999), .B1(n14723), .B2(n1000), .ZN(n13574)
         );
  OAI22_X1 U5952 ( .A1(n7534), .A2(n999), .B1(n14683), .B2(n1000), .ZN(n13575)
         );
  OAI22_X1 U5953 ( .A1(n7518), .A2(n1001), .B1(n14945), .B2(n1002), .ZN(n13576) );
  OAI22_X1 U5954 ( .A1(n7502), .A2(n1001), .B1(n14923), .B2(n1002), .ZN(n13577) );
  OAI22_X1 U5955 ( .A1(n7486), .A2(n1001), .B1(n14883), .B2(n1002), .ZN(n13578) );
  OAI22_X1 U5956 ( .A1(n7470), .A2(n1001), .B1(n14843), .B2(n1002), .ZN(n13579) );
  OAI22_X1 U5957 ( .A1(n7454), .A2(n1001), .B1(n14803), .B2(n1002), .ZN(n13580) );
  OAI22_X1 U5958 ( .A1(n7438), .A2(n1001), .B1(n14763), .B2(n1002), .ZN(n13581) );
  OAI22_X1 U5959 ( .A1(n7422), .A2(n1001), .B1(n14723), .B2(n1002), .ZN(n13582) );
  OAI22_X1 U5960 ( .A1(n7406), .A2(n1001), .B1(n14683), .B2(n1002), .ZN(n13583) );
  OAI22_X1 U5961 ( .A1(n7390), .A2(n1003), .B1(n14945), .B2(n1004), .ZN(n13584) );
  OAI22_X1 U5962 ( .A1(n7374), .A2(n1003), .B1(n14923), .B2(n1004), .ZN(n13585) );
  OAI22_X1 U5963 ( .A1(n7358), .A2(n1003), .B1(n14883), .B2(n1004), .ZN(n13586) );
  OAI22_X1 U5964 ( .A1(n7342), .A2(n1003), .B1(n14843), .B2(n1004), .ZN(n13587) );
  OAI22_X1 U5965 ( .A1(n7326), .A2(n1003), .B1(n14803), .B2(n1004), .ZN(n13588) );
  OAI22_X1 U5966 ( .A1(n7310), .A2(n1003), .B1(n14763), .B2(n1004), .ZN(n13589) );
  OAI22_X1 U5967 ( .A1(n7294), .A2(n1003), .B1(n14723), .B2(n1004), .ZN(n13590) );
  OAI22_X1 U5968 ( .A1(n7278), .A2(n1003), .B1(n14683), .B2(n1004), .ZN(n13591) );
  OAI22_X1 U5969 ( .A1(n7262), .A2(n1005), .B1(n14945), .B2(n1006), .ZN(n13592) );
  OAI22_X1 U5970 ( .A1(n7246), .A2(n1005), .B1(n14923), .B2(n1006), .ZN(n13593) );
  OAI22_X1 U5971 ( .A1(n7230), .A2(n1005), .B1(n14883), .B2(n1006), .ZN(n13594) );
  OAI22_X1 U5972 ( .A1(n7214), .A2(n1005), .B1(n14843), .B2(n1006), .ZN(n13595) );
  OAI22_X1 U5973 ( .A1(n7198), .A2(n1005), .B1(n14803), .B2(n1006), .ZN(n13596) );
  OAI22_X1 U5974 ( .A1(n7182), .A2(n1005), .B1(n14763), .B2(n1006), .ZN(n13597) );
  OAI22_X1 U5975 ( .A1(n7166), .A2(n1005), .B1(n14723), .B2(n1006), .ZN(n13598) );
  OAI22_X1 U5976 ( .A1(n7150), .A2(n1005), .B1(n14683), .B2(n1006), .ZN(n13599) );
  OAI22_X1 U5977 ( .A1(n7134), .A2(n1007), .B1(n14945), .B2(n1008), .ZN(n13600) );
  OAI22_X1 U5978 ( .A1(n7118), .A2(n1007), .B1(n14923), .B2(n1008), .ZN(n13601) );
  OAI22_X1 U5979 ( .A1(n7102), .A2(n1007), .B1(n14883), .B2(n1008), .ZN(n13602) );
  OAI22_X1 U5980 ( .A1(n7086), .A2(n1007), .B1(n14843), .B2(n1008), .ZN(n13603) );
  OAI22_X1 U5981 ( .A1(n7070), .A2(n1007), .B1(n14803), .B2(n1008), .ZN(n13604) );
  OAI22_X1 U5982 ( .A1(n7054), .A2(n1007), .B1(n14763), .B2(n1008), .ZN(n13605) );
  OAI22_X1 U5983 ( .A1(n7038), .A2(n1007), .B1(n14723), .B2(n1008), .ZN(n13606) );
  OAI22_X1 U5984 ( .A1(n7022), .A2(n1007), .B1(n14683), .B2(n1008), .ZN(n13607) );
  OAI22_X1 U5985 ( .A1(n7006), .A2(n1009), .B1(n14945), .B2(n1010), .ZN(n13608) );
  OAI22_X1 U5986 ( .A1(n6990), .A2(n1009), .B1(n14923), .B2(n1010), .ZN(n13609) );
  OAI22_X1 U5987 ( .A1(n6974), .A2(n1009), .B1(n14883), .B2(n1010), .ZN(n13610) );
  OAI22_X1 U5988 ( .A1(n6958), .A2(n1009), .B1(n14843), .B2(n1010), .ZN(n13611) );
  OAI22_X1 U5989 ( .A1(n6942), .A2(n1009), .B1(n14803), .B2(n1010), .ZN(n13612) );
  OAI22_X1 U5990 ( .A1(n6926), .A2(n1009), .B1(n14763), .B2(n1010), .ZN(n13613) );
  OAI22_X1 U5991 ( .A1(n6910), .A2(n1009), .B1(n14723), .B2(n1010), .ZN(n13614) );
  OAI22_X1 U5992 ( .A1(n6894), .A2(n1009), .B1(n14683), .B2(n1010), .ZN(n13615) );
  OAI22_X1 U5993 ( .A1(n6878), .A2(n1011), .B1(n14945), .B2(n1012), .ZN(n13616) );
  OAI22_X1 U5994 ( .A1(n6862), .A2(n1011), .B1(n14923), .B2(n1012), .ZN(n13617) );
  OAI22_X1 U5995 ( .A1(n6846), .A2(n1011), .B1(n14883), .B2(n1012), .ZN(n13618) );
  OAI22_X1 U5996 ( .A1(n6830), .A2(n1011), .B1(n14843), .B2(n1012), .ZN(n13619) );
  OAI22_X1 U5997 ( .A1(n6814), .A2(n1011), .B1(n14803), .B2(n1012), .ZN(n13620) );
  OAI22_X1 U5998 ( .A1(n6798), .A2(n1011), .B1(n14763), .B2(n1012), .ZN(n13621) );
  OAI22_X1 U5999 ( .A1(n6782), .A2(n1011), .B1(n14723), .B2(n1012), .ZN(n13622) );
  OAI22_X1 U6000 ( .A1(n6766), .A2(n1011), .B1(n14683), .B2(n1012), .ZN(n13623) );
  OAI22_X1 U6001 ( .A1(n10086), .A2(n1091), .B1(n14942), .B2(n1092), .ZN(
        n13928) );
  OAI22_X1 U6002 ( .A1(n10070), .A2(n1091), .B1(n14926), .B2(n1092), .ZN(
        n13929) );
  OAI22_X1 U6003 ( .A1(n10054), .A2(n1091), .B1(n14886), .B2(n1092), .ZN(
        n13930) );
  OAI22_X1 U6004 ( .A1(n10038), .A2(n1091), .B1(n14846), .B2(n1092), .ZN(
        n13931) );
  OAI22_X1 U6005 ( .A1(n10022), .A2(n1091), .B1(n14806), .B2(n1092), .ZN(
        n13932) );
  OAI22_X1 U6006 ( .A1(n10006), .A2(n1091), .B1(n14766), .B2(n1092), .ZN(
        n13933) );
  OAI22_X1 U6007 ( .A1(n9990), .A2(n1091), .B1(n14726), .B2(n1092), .ZN(n13934) );
  OAI22_X1 U6008 ( .A1(n9974), .A2(n1091), .B1(n14686), .B2(n1092), .ZN(n13935) );
  OAI22_X1 U6009 ( .A1(n9958), .A2(n1096), .B1(n14942), .B2(n1097), .ZN(n13936) );
  OAI22_X1 U6010 ( .A1(n9942), .A2(n1096), .B1(n14927), .B2(n1097), .ZN(n13937) );
  OAI22_X1 U6011 ( .A1(n9926), .A2(n1096), .B1(n14887), .B2(n1097), .ZN(n13938) );
  OAI22_X1 U6012 ( .A1(n9910), .A2(n1096), .B1(n14847), .B2(n1097), .ZN(n13939) );
  OAI22_X1 U6013 ( .A1(n9894), .A2(n1096), .B1(n14807), .B2(n1097), .ZN(n13940) );
  OAI22_X1 U6014 ( .A1(n9878), .A2(n1096), .B1(n14767), .B2(n1097), .ZN(n13941) );
  OAI22_X1 U6015 ( .A1(n9862), .A2(n1096), .B1(n14727), .B2(n1097), .ZN(n13942) );
  OAI22_X1 U6016 ( .A1(n9846), .A2(n1096), .B1(n14687), .B2(n1097), .ZN(n13943) );
  OAI22_X1 U6017 ( .A1(n9830), .A2(n1099), .B1(n14942), .B2(n1100), .ZN(n13944) );
  OAI22_X1 U6018 ( .A1(n9814), .A2(n1099), .B1(n14927), .B2(n1100), .ZN(n13945) );
  OAI22_X1 U6019 ( .A1(n9798), .A2(n1099), .B1(n14887), .B2(n1100), .ZN(n13946) );
  OAI22_X1 U6020 ( .A1(n9782), .A2(n1099), .B1(n14847), .B2(n1100), .ZN(n13947) );
  OAI22_X1 U6021 ( .A1(n9766), .A2(n1099), .B1(n14807), .B2(n1100), .ZN(n13948) );
  OAI22_X1 U6022 ( .A1(n9750), .A2(n1099), .B1(n14767), .B2(n1100), .ZN(n13949) );
  OAI22_X1 U6023 ( .A1(n9734), .A2(n1099), .B1(n14727), .B2(n1100), .ZN(n13950) );
  OAI22_X1 U6024 ( .A1(n9718), .A2(n1099), .B1(n14687), .B2(n1100), .ZN(n13951) );
  OAI22_X1 U6025 ( .A1(n9702), .A2(n1102), .B1(n14941), .B2(n1103), .ZN(n13952) );
  OAI22_X1 U6026 ( .A1(n9686), .A2(n1102), .B1(n14927), .B2(n1103), .ZN(n13953) );
  OAI22_X1 U6027 ( .A1(n9670), .A2(n1102), .B1(n14887), .B2(n1103), .ZN(n13954) );
  OAI22_X1 U6028 ( .A1(n9654), .A2(n1102), .B1(n14847), .B2(n1103), .ZN(n13955) );
  OAI22_X1 U6029 ( .A1(n9638), .A2(n1102), .B1(n14807), .B2(n1103), .ZN(n13956) );
  OAI22_X1 U6030 ( .A1(n9622), .A2(n1102), .B1(n14767), .B2(n1103), .ZN(n13957) );
  OAI22_X1 U6031 ( .A1(n9606), .A2(n1102), .B1(n14727), .B2(n1103), .ZN(n13958) );
  OAI22_X1 U6032 ( .A1(n9590), .A2(n1102), .B1(n14687), .B2(n1103), .ZN(n13959) );
  OAI22_X1 U6033 ( .A1(n9574), .A2(n1105), .B1(n14941), .B2(n1106), .ZN(n13960) );
  OAI22_X1 U6034 ( .A1(n9558), .A2(n1105), .B1(n14927), .B2(n1106), .ZN(n13961) );
  OAI22_X1 U6035 ( .A1(n9542), .A2(n1105), .B1(n14887), .B2(n1106), .ZN(n13962) );
  OAI22_X1 U6036 ( .A1(n9526), .A2(n1105), .B1(n14847), .B2(n1106), .ZN(n13963) );
  OAI22_X1 U6037 ( .A1(n9510), .A2(n1105), .B1(n14807), .B2(n1106), .ZN(n13964) );
  OAI22_X1 U6038 ( .A1(n9494), .A2(n1105), .B1(n14767), .B2(n1106), .ZN(n13965) );
  OAI22_X1 U6039 ( .A1(n9478), .A2(n1105), .B1(n14727), .B2(n1106), .ZN(n13966) );
  OAI22_X1 U6040 ( .A1(n9462), .A2(n1105), .B1(n14687), .B2(n1106), .ZN(n13967) );
  OAI22_X1 U6041 ( .A1(n9446), .A2(n1108), .B1(n14941), .B2(n1109), .ZN(n13968) );
  OAI22_X1 U6042 ( .A1(n9430), .A2(n1108), .B1(n14927), .B2(n1109), .ZN(n13969) );
  OAI22_X1 U6043 ( .A1(n9414), .A2(n1108), .B1(n14887), .B2(n1109), .ZN(n13970) );
  OAI22_X1 U6044 ( .A1(n9398), .A2(n1108), .B1(n14847), .B2(n1109), .ZN(n13971) );
  OAI22_X1 U6045 ( .A1(n9382), .A2(n1108), .B1(n14807), .B2(n1109), .ZN(n13972) );
  OAI22_X1 U6046 ( .A1(n9366), .A2(n1108), .B1(n14767), .B2(n1109), .ZN(n13973) );
  OAI22_X1 U6047 ( .A1(n9350), .A2(n1108), .B1(n14727), .B2(n1109), .ZN(n13974) );
  OAI22_X1 U6048 ( .A1(n9334), .A2(n1108), .B1(n14687), .B2(n1109), .ZN(n13975) );
  OAI22_X1 U6049 ( .A1(n9318), .A2(n1110), .B1(n14941), .B2(n1111), .ZN(n13976) );
  OAI22_X1 U6050 ( .A1(n9302), .A2(n1110), .B1(n14927), .B2(n1111), .ZN(n13977) );
  OAI22_X1 U6051 ( .A1(n9286), .A2(n1110), .B1(n14887), .B2(n1111), .ZN(n13978) );
  OAI22_X1 U6052 ( .A1(n9270), .A2(n1110), .B1(n14847), .B2(n1111), .ZN(n13979) );
  OAI22_X1 U6053 ( .A1(n9254), .A2(n1110), .B1(n14807), .B2(n1111), .ZN(n13980) );
  OAI22_X1 U6054 ( .A1(n9238), .A2(n1110), .B1(n14767), .B2(n1111), .ZN(n13981) );
  OAI22_X1 U6055 ( .A1(n9222), .A2(n1110), .B1(n14727), .B2(n1111), .ZN(n13982) );
  OAI22_X1 U6056 ( .A1(n9206), .A2(n1110), .B1(n14687), .B2(n1111), .ZN(n13983) );
  OAI22_X1 U6057 ( .A1(n9190), .A2(n1112), .B1(n14941), .B2(n1113), .ZN(n13984) );
  OAI22_X1 U6058 ( .A1(n9174), .A2(n1112), .B1(n14927), .B2(n1113), .ZN(n13985) );
  OAI22_X1 U6059 ( .A1(n9158), .A2(n1112), .B1(n14887), .B2(n1113), .ZN(n13986) );
  OAI22_X1 U6060 ( .A1(n9142), .A2(n1112), .B1(n14847), .B2(n1113), .ZN(n13987) );
  OAI22_X1 U6061 ( .A1(n9126), .A2(n1112), .B1(n14807), .B2(n1113), .ZN(n13988) );
  OAI22_X1 U6062 ( .A1(n9110), .A2(n1112), .B1(n14767), .B2(n1113), .ZN(n13989) );
  OAI22_X1 U6063 ( .A1(n9094), .A2(n1112), .B1(n14727), .B2(n1113), .ZN(n13990) );
  OAI22_X1 U6064 ( .A1(n9078), .A2(n1112), .B1(n14687), .B2(n1113), .ZN(n13991) );
  OAI22_X1 U6065 ( .A1(n9062), .A2(n1114), .B1(n14941), .B2(n1115), .ZN(n13992) );
  OAI22_X1 U6066 ( .A1(n9046), .A2(n1114), .B1(n14927), .B2(n1115), .ZN(n13993) );
  OAI22_X1 U6067 ( .A1(n9030), .A2(n1114), .B1(n14887), .B2(n1115), .ZN(n13994) );
  OAI22_X1 U6068 ( .A1(n9014), .A2(n1114), .B1(n14847), .B2(n1115), .ZN(n13995) );
  OAI22_X1 U6069 ( .A1(n8998), .A2(n1114), .B1(n14807), .B2(n1115), .ZN(n13996) );
  OAI22_X1 U6070 ( .A1(n8982), .A2(n1114), .B1(n14767), .B2(n1115), .ZN(n13997) );
  OAI22_X1 U6071 ( .A1(n8966), .A2(n1114), .B1(n14727), .B2(n1115), .ZN(n13998) );
  OAI22_X1 U6072 ( .A1(n8950), .A2(n1114), .B1(n14687), .B2(n1115), .ZN(n13999) );
  OAI22_X1 U6073 ( .A1(n8934), .A2(n1117), .B1(n14941), .B2(n1118), .ZN(n14000) );
  OAI22_X1 U6074 ( .A1(n8918), .A2(n1117), .B1(n14927), .B2(n1118), .ZN(n14001) );
  OAI22_X1 U6075 ( .A1(n8902), .A2(n1117), .B1(n14887), .B2(n1118), .ZN(n14002) );
  OAI22_X1 U6076 ( .A1(n8886), .A2(n1117), .B1(n14847), .B2(n1118), .ZN(n14003) );
  OAI22_X1 U6077 ( .A1(n8870), .A2(n1117), .B1(n14807), .B2(n1118), .ZN(n14004) );
  OAI22_X1 U6078 ( .A1(n8854), .A2(n1117), .B1(n14767), .B2(n1118), .ZN(n14005) );
  OAI22_X1 U6079 ( .A1(n8838), .A2(n1117), .B1(n14727), .B2(n1118), .ZN(n14006) );
  OAI22_X1 U6080 ( .A1(n8822), .A2(n1117), .B1(n14687), .B2(n1118), .ZN(n14007) );
  OAI22_X1 U6081 ( .A1(n8806), .A2(n1119), .B1(n14941), .B2(n1120), .ZN(n14008) );
  OAI22_X1 U6082 ( .A1(n8790), .A2(n1119), .B1(n14927), .B2(n1120), .ZN(n14009) );
  OAI22_X1 U6083 ( .A1(n8774), .A2(n1119), .B1(n14887), .B2(n1120), .ZN(n14010) );
  OAI22_X1 U6084 ( .A1(n8758), .A2(n1119), .B1(n14847), .B2(n1120), .ZN(n14011) );
  OAI22_X1 U6085 ( .A1(n8742), .A2(n1119), .B1(n14807), .B2(n1120), .ZN(n14012) );
  OAI22_X1 U6086 ( .A1(n8726), .A2(n1119), .B1(n14767), .B2(n1120), .ZN(n14013) );
  OAI22_X1 U6087 ( .A1(n8710), .A2(n1119), .B1(n14727), .B2(n1120), .ZN(n14014) );
  OAI22_X1 U6088 ( .A1(n8694), .A2(n1119), .B1(n14687), .B2(n1120), .ZN(n14015) );
  OAI22_X1 U6089 ( .A1(n8678), .A2(n1121), .B1(n14941), .B2(n1122), .ZN(n14016) );
  OAI22_X1 U6090 ( .A1(n8662), .A2(n1121), .B1(n14927), .B2(n1122), .ZN(n14017) );
  OAI22_X1 U6091 ( .A1(n8646), .A2(n1121), .B1(n14887), .B2(n1122), .ZN(n14018) );
  OAI22_X1 U6092 ( .A1(n8630), .A2(n1121), .B1(n14847), .B2(n1122), .ZN(n14019) );
  OAI22_X1 U6093 ( .A1(n8614), .A2(n1121), .B1(n14807), .B2(n1122), .ZN(n14020) );
  OAI22_X1 U6094 ( .A1(n8598), .A2(n1121), .B1(n14767), .B2(n1122), .ZN(n14021) );
  OAI22_X1 U6095 ( .A1(n8582), .A2(n1121), .B1(n14727), .B2(n1122), .ZN(n14022) );
  OAI22_X1 U6097 ( .A1(n8566), .A2(n1121), .B1(n14687), .B2(n1122), .ZN(n14023) );
  OAI22_X1 U6098 ( .A1(n8550), .A2(n1123), .B1(n14941), .B2(n1124), .ZN(n14024) );
  OAI22_X1 U6099 ( .A1(n8534), .A2(n1123), .B1(n14927), .B2(n1124), .ZN(n14025) );
  OAI22_X1 U6100 ( .A1(n8518), .A2(n1123), .B1(n14887), .B2(n1124), .ZN(n14026) );
  OAI22_X1 U6101 ( .A1(n8502), .A2(n1123), .B1(n14847), .B2(n1124), .ZN(n14027) );
  OAI22_X1 U6102 ( .A1(n8486), .A2(n1123), .B1(n14807), .B2(n1124), .ZN(n14028) );
  OAI22_X1 U6103 ( .A1(n8470), .A2(n1123), .B1(n14767), .B2(n1124), .ZN(n14029) );
  OAI22_X1 U6104 ( .A1(n8454), .A2(n1123), .B1(n14727), .B2(n1124), .ZN(n14030) );
  OAI22_X1 U6105 ( .A1(n8438), .A2(n1123), .B1(n14687), .B2(n1124), .ZN(n14031) );
  OAI22_X1 U6106 ( .A1(n8422), .A2(n1126), .B1(n14941), .B2(n1127), .ZN(n14032) );
  OAI22_X1 U6107 ( .A1(n8406), .A2(n1126), .B1(n14927), .B2(n1127), .ZN(n14033) );
  OAI22_X1 U6108 ( .A1(n8390), .A2(n1126), .B1(n14887), .B2(n1127), .ZN(n14034) );
  OAI22_X1 U6109 ( .A1(n8374), .A2(n1126), .B1(n14847), .B2(n1127), .ZN(n14035) );
  OAI22_X1 U6110 ( .A1(n8358), .A2(n1126), .B1(n14807), .B2(n1127), .ZN(n14036) );
  OAI22_X1 U6111 ( .A1(n8342), .A2(n1126), .B1(n14767), .B2(n1127), .ZN(n14037) );
  OAI22_X1 U6112 ( .A1(n8326), .A2(n1126), .B1(n14727), .B2(n1127), .ZN(n14038) );
  OAI22_X1 U6113 ( .A1(n8310), .A2(n1126), .B1(n14687), .B2(n1127), .ZN(n14039) );
  OAI22_X1 U6114 ( .A1(n8294), .A2(n1128), .B1(n14941), .B2(n1129), .ZN(n14040) );
  OAI22_X1 U6115 ( .A1(n8278), .A2(n1128), .B1(n14928), .B2(n1129), .ZN(n14041) );
  OAI22_X1 U6116 ( .A1(n8262), .A2(n1128), .B1(n14888), .B2(n1129), .ZN(n14042) );
  OAI22_X1 U6117 ( .A1(n8246), .A2(n1128), .B1(n14848), .B2(n1129), .ZN(n14043) );
  OAI22_X1 U6118 ( .A1(n8230), .A2(n1128), .B1(n14808), .B2(n1129), .ZN(n14044) );
  OAI22_X1 U6119 ( .A1(n8214), .A2(n1128), .B1(n14768), .B2(n1129), .ZN(n14045) );
  OAI22_X1 U6120 ( .A1(n8198), .A2(n1128), .B1(n14728), .B2(n1129), .ZN(n14046) );
  OAI22_X1 U6121 ( .A1(n8182), .A2(n1128), .B1(n14688), .B2(n1129), .ZN(n14047) );
  OAI22_X1 U6122 ( .A1(n8166), .A2(n1130), .B1(n14941), .B2(n1131), .ZN(n14048) );
  OAI22_X1 U6123 ( .A1(n8150), .A2(n1130), .B1(n14928), .B2(n1131), .ZN(n14049) );
  OAI22_X1 U6124 ( .A1(n8134), .A2(n1130), .B1(n14888), .B2(n1131), .ZN(n14050) );
  OAI22_X1 U6125 ( .A1(n8118), .A2(n1130), .B1(n14848), .B2(n1131), .ZN(n14051) );
  OAI22_X1 U6126 ( .A1(n8102), .A2(n1130), .B1(n14808), .B2(n1131), .ZN(n14052) );
  OAI22_X1 U6127 ( .A1(n8086), .A2(n1130), .B1(n14768), .B2(n1131), .ZN(n14053) );
  OAI22_X1 U6128 ( .A1(n8070), .A2(n1130), .B1(n14728), .B2(n1131), .ZN(n14054) );
  OAI22_X1 U6129 ( .A1(n8054), .A2(n1130), .B1(n14688), .B2(n1131), .ZN(n14055) );
  OAI22_X1 U6130 ( .A1(n8038), .A2(n1132), .B1(n14940), .B2(n1133), .ZN(n14056) );
  OAI22_X1 U6131 ( .A1(n8022), .A2(n1132), .B1(n14928), .B2(n1133), .ZN(n14057) );
  OAI22_X1 U6132 ( .A1(n8006), .A2(n1132), .B1(n14888), .B2(n1133), .ZN(n14058) );
  OAI22_X1 U6133 ( .A1(n7990), .A2(n1132), .B1(n14848), .B2(n1133), .ZN(n14059) );
  OAI22_X1 U6134 ( .A1(n7974), .A2(n1132), .B1(n14808), .B2(n1133), .ZN(n14060) );
  OAI22_X1 U6135 ( .A1(n7958), .A2(n1132), .B1(n14768), .B2(n1133), .ZN(n14061) );
  OAI22_X1 U6136 ( .A1(n7942), .A2(n1132), .B1(n14728), .B2(n1133), .ZN(n14062) );
  OAI22_X1 U6137 ( .A1(n7926), .A2(n1132), .B1(n14688), .B2(n1133), .ZN(n14063) );
  OAI22_X1 U6138 ( .A1(n7910), .A2(n1135), .B1(n14940), .B2(n1136), .ZN(n14064) );
  OAI22_X1 U6139 ( .A1(n7894), .A2(n1135), .B1(n14928), .B2(n1136), .ZN(n14065) );
  OAI22_X1 U6140 ( .A1(n7878), .A2(n1135), .B1(n14888), .B2(n1136), .ZN(n14066) );
  OAI22_X1 U6141 ( .A1(n7862), .A2(n1135), .B1(n14848), .B2(n1136), .ZN(n14067) );
  OAI22_X1 U6142 ( .A1(n7846), .A2(n1135), .B1(n14808), .B2(n1136), .ZN(n14068) );
  OAI22_X1 U6143 ( .A1(n7830), .A2(n1135), .B1(n14768), .B2(n1136), .ZN(n14069) );
  OAI22_X1 U6144 ( .A1(n7814), .A2(n1135), .B1(n14728), .B2(n1136), .ZN(n14070) );
  OAI22_X1 U6145 ( .A1(n7798), .A2(n1135), .B1(n14688), .B2(n1136), .ZN(n14071) );
  OAI22_X1 U6146 ( .A1(n7782), .A2(n1137), .B1(n14940), .B2(n1138), .ZN(n14072) );
  OAI22_X1 U6147 ( .A1(n7766), .A2(n1137), .B1(n14928), .B2(n1138), .ZN(n14073) );
  OAI22_X1 U6148 ( .A1(n7750), .A2(n1137), .B1(n14888), .B2(n1138), .ZN(n14074) );
  OAI22_X1 U6149 ( .A1(n7734), .A2(n1137), .B1(n14848), .B2(n1138), .ZN(n14075) );
  OAI22_X1 U6150 ( .A1(n7718), .A2(n1137), .B1(n14808), .B2(n1138), .ZN(n14076) );
  OAI22_X1 U6151 ( .A1(n7702), .A2(n1137), .B1(n14768), .B2(n1138), .ZN(n14077) );
  OAI22_X1 U6152 ( .A1(n7686), .A2(n1137), .B1(n14728), .B2(n1138), .ZN(n14078) );
  OAI22_X1 U6153 ( .A1(n7670), .A2(n1137), .B1(n14688), .B2(n1138), .ZN(n14079) );
  OAI22_X1 U6154 ( .A1(n7654), .A2(n1139), .B1(n14940), .B2(n1140), .ZN(n14080) );
  OAI22_X1 U6155 ( .A1(n7638), .A2(n1139), .B1(n14928), .B2(n1140), .ZN(n14081) );
  OAI22_X1 U6156 ( .A1(n7622), .A2(n1139), .B1(n14888), .B2(n1140), .ZN(n14082) );
  OAI22_X1 U6157 ( .A1(n7606), .A2(n1139), .B1(n14848), .B2(n1140), .ZN(n14083) );
  OAI22_X1 U6158 ( .A1(n7590), .A2(n1139), .B1(n14808), .B2(n1140), .ZN(n14084) );
  OAI22_X1 U6159 ( .A1(n7574), .A2(n1139), .B1(n14768), .B2(n1140), .ZN(n14085) );
  OAI22_X1 U6160 ( .A1(n7558), .A2(n1139), .B1(n14728), .B2(n1140), .ZN(n14086) );
  OAI22_X1 U6161 ( .A1(n7542), .A2(n1139), .B1(n14688), .B2(n1140), .ZN(n14087) );
  OAI22_X1 U6162 ( .A1(n7526), .A2(n1141), .B1(n14940), .B2(n1142), .ZN(n14088) );
  OAI22_X1 U6163 ( .A1(n7510), .A2(n1141), .B1(n14928), .B2(n1142), .ZN(n14089) );
  OAI22_X1 U6164 ( .A1(n7494), .A2(n1141), .B1(n14888), .B2(n1142), .ZN(n14090) );
  OAI22_X1 U6165 ( .A1(n7478), .A2(n1141), .B1(n14848), .B2(n1142), .ZN(n14091) );
  OAI22_X1 U6166 ( .A1(n7462), .A2(n1141), .B1(n14808), .B2(n1142), .ZN(n14092) );
  OAI22_X1 U6167 ( .A1(n7446), .A2(n1141), .B1(n14768), .B2(n1142), .ZN(n14093) );
  OAI22_X1 U6168 ( .A1(n7430), .A2(n1141), .B1(n14728), .B2(n1142), .ZN(n14094) );
  OAI22_X1 U6169 ( .A1(n7414), .A2(n1141), .B1(n14688), .B2(n1142), .ZN(n14095) );
  OAI22_X1 U6170 ( .A1(n7398), .A2(n1144), .B1(n14940), .B2(n1145), .ZN(n14096) );
  OAI22_X1 U6171 ( .A1(n7382), .A2(n1144), .B1(n14928), .B2(n1145), .ZN(n14097) );
  OAI22_X1 U6172 ( .A1(n7366), .A2(n1144), .B1(n14888), .B2(n1145), .ZN(n14098) );
  OAI22_X1 U6173 ( .A1(n7350), .A2(n1144), .B1(n14848), .B2(n1145), .ZN(n14099) );
  OAI22_X1 U6174 ( .A1(n7334), .A2(n1144), .B1(n14808), .B2(n1145), .ZN(n14100) );
  OAI22_X1 U6175 ( .A1(n7318), .A2(n1144), .B1(n14768), .B2(n1145), .ZN(n14101) );
  OAI22_X1 U6176 ( .A1(n7302), .A2(n1144), .B1(n14728), .B2(n1145), .ZN(n14102) );
  OAI22_X1 U6177 ( .A1(n7286), .A2(n1144), .B1(n14688), .B2(n1145), .ZN(n14103) );
  OAI22_X1 U6178 ( .A1(n7270), .A2(n1146), .B1(n14940), .B2(n1147), .ZN(n14104) );
  OAI22_X1 U6179 ( .A1(n7254), .A2(n1146), .B1(n14928), .B2(n1147), .ZN(n14105) );
  OAI22_X1 U6180 ( .A1(n7238), .A2(n1146), .B1(n14888), .B2(n1147), .ZN(n14106) );
  OAI22_X1 U6181 ( .A1(n7222), .A2(n1146), .B1(n14848), .B2(n1147), .ZN(n14107) );
  OAI22_X1 U6182 ( .A1(n7206), .A2(n1146), .B1(n14808), .B2(n1147), .ZN(n14108) );
  OAI22_X1 U6183 ( .A1(n7190), .A2(n1146), .B1(n14768), .B2(n1147), .ZN(n14109) );
  OAI22_X1 U6184 ( .A1(n7174), .A2(n1146), .B1(n14728), .B2(n1147), .ZN(n14110) );
  OAI22_X1 U6185 ( .A1(n7158), .A2(n1146), .B1(n14688), .B2(n1147), .ZN(n14111) );
  OAI22_X1 U6186 ( .A1(n7142), .A2(n1148), .B1(n14940), .B2(n1149), .ZN(n14112) );
  OAI22_X1 U6187 ( .A1(n7126), .A2(n1148), .B1(n14928), .B2(n1149), .ZN(n14113) );
  OAI22_X1 U6188 ( .A1(n7110), .A2(n1148), .B1(n14888), .B2(n1149), .ZN(n14114) );
  OAI22_X1 U6189 ( .A1(n7094), .A2(n1148), .B1(n14848), .B2(n1149), .ZN(n14115) );
  OAI22_X1 U6190 ( .A1(n7078), .A2(n1148), .B1(n14808), .B2(n1149), .ZN(n14116) );
  OAI22_X1 U6191 ( .A1(n7062), .A2(n1148), .B1(n14768), .B2(n1149), .ZN(n14117) );
  OAI22_X1 U6192 ( .A1(n7046), .A2(n1148), .B1(n14728), .B2(n1149), .ZN(n14118) );
  OAI22_X1 U6193 ( .A1(n7030), .A2(n1148), .B1(n14688), .B2(n1149), .ZN(n14119) );
  OAI22_X1 U6194 ( .A1(n7014), .A2(n1150), .B1(n14940), .B2(n1151), .ZN(n14120) );
  OAI22_X1 U6195 ( .A1(n6998), .A2(n1150), .B1(n14928), .B2(n1151), .ZN(n14121) );
  OAI22_X1 U6196 ( .A1(n6982), .A2(n1150), .B1(n14888), .B2(n1151), .ZN(n14122) );
  OAI22_X1 U6197 ( .A1(n6966), .A2(n1150), .B1(n14848), .B2(n1151), .ZN(n14123) );
  OAI22_X1 U6198 ( .A1(n6950), .A2(n1150), .B1(n14808), .B2(n1151), .ZN(n14124) );
  OAI22_X1 U6199 ( .A1(n6934), .A2(n1150), .B1(n14768), .B2(n1151), .ZN(n14125) );
  OAI22_X1 U6200 ( .A1(n6918), .A2(n1150), .B1(n14728), .B2(n1151), .ZN(n14126) );
  OAI22_X1 U6201 ( .A1(n6902), .A2(n1150), .B1(n14688), .B2(n1151), .ZN(n14127) );
  OAI22_X1 U6202 ( .A1(n6886), .A2(n1153), .B1(n14940), .B2(n1154), .ZN(n14128) );
  OAI22_X1 U6203 ( .A1(n6870), .A2(n1153), .B1(n14928), .B2(n1154), .ZN(n14129) );
  OAI22_X1 U6204 ( .A1(n6854), .A2(n1153), .B1(n14888), .B2(n1154), .ZN(n14130) );
  OAI22_X1 U6205 ( .A1(n6838), .A2(n1153), .B1(n14848), .B2(n1154), .ZN(n14131) );
  OAI22_X1 U6206 ( .A1(n6822), .A2(n1153), .B1(n14808), .B2(n1154), .ZN(n14132) );
  OAI22_X1 U6207 ( .A1(n6806), .A2(n1153), .B1(n14768), .B2(n1154), .ZN(n14133) );
  OAI22_X1 U6208 ( .A1(n6790), .A2(n1153), .B1(n14728), .B2(n1154), .ZN(n14134) );
  OAI22_X1 U6209 ( .A1(n6774), .A2(n1153), .B1(n14688), .B2(n1154), .ZN(n14135) );
  OAI22_X1 U6210 ( .A1(n14968), .A2(n381), .B1(n9435), .B2(n382), .ZN(n11152)
         );
  OAI22_X1 U6211 ( .A1(n14968), .A2(n383), .B1(n9307), .B2(n384), .ZN(n11160)
         );
  OAI22_X1 U6212 ( .A1(n14968), .A2(n385), .B1(n9179), .B2(n386), .ZN(n11168)
         );
  OAI22_X1 U6213 ( .A1(n14968), .A2(n387), .B1(n9051), .B2(n388), .ZN(n11176)
         );
  OAI22_X1 U6214 ( .A1(n14968), .A2(n389), .B1(n8923), .B2(n390), .ZN(n11184)
         );
  OAI22_X1 U6215 ( .A1(n14968), .A2(n391), .B1(n8795), .B2(n392), .ZN(n11192)
         );
  OAI22_X1 U6216 ( .A1(n14968), .A2(n393), .B1(n8667), .B2(n394), .ZN(n11200)
         );
  OAI22_X1 U6217 ( .A1(n14968), .A2(n395), .B1(n8539), .B2(n396), .ZN(n11208)
         );
  INV_X1 U6218 ( .A(ADDR[0]), .ZN(n14982) );
  AND2_X1 U6219 ( .A1(ADDR[3]), .A2(ADDR[2]), .ZN(n5953) );
  NOR2_X1 U6220 ( .A1(n5960), .A2(n14970), .ZN(n14186) );
  NOR2_X1 U6221 ( .A1(n5961), .A2(n14970), .ZN(n14189) );
  NOR2_X1 U6222 ( .A1(n5962), .A2(n14970), .ZN(n14192) );
  NOR2_X1 U6223 ( .A1(n5963), .A2(n14971), .ZN(n14195) );
  NOR2_X1 U6224 ( .A1(n5964), .A2(n14970), .ZN(n14198) );
  NOR2_X1 U6225 ( .A1(n5965), .A2(n14971), .ZN(n14201) );
  NOR2_X1 U6226 ( .A1(n5966), .A2(n14971), .ZN(n14204) );
  NOR2_X1 U6227 ( .A1(n5967), .A2(n14971), .ZN(n14207) );
  NOR2_X1 U6228 ( .A1(n5968), .A2(n14971), .ZN(n14210) );
  NOR2_X1 U6229 ( .A1(n5969), .A2(n14971), .ZN(n14213) );
  NOR2_X1 U6230 ( .A1(n5970), .A2(n14971), .ZN(n14216) );
  NOR2_X1 U6231 ( .A1(n5971), .A2(n14971), .ZN(n14219) );
  NOR2_X1 U6232 ( .A1(n5972), .A2(n14970), .ZN(n14222) );
  NOR2_X1 U6233 ( .A1(n5973), .A2(n14971), .ZN(n14225) );
  NOR2_X1 U6234 ( .A1(n5974), .A2(n14971), .ZN(n14228) );
  NOR2_X1 U6235 ( .A1(n5975), .A2(n14970), .ZN(n14231) );
  NOR2_X1 U6236 ( .A1(n5976), .A2(n14971), .ZN(n14234) );
  NOR2_X1 U6237 ( .A1(n5977), .A2(n14970), .ZN(n14237) );
  NOR2_X1 U6238 ( .A1(n5978), .A2(n14970), .ZN(n14240) );
  NOR2_X1 U6239 ( .A1(n5979), .A2(n14971), .ZN(n14243) );
  NOR2_X1 U6240 ( .A1(n5980), .A2(n14971), .ZN(n14246) );
  NOR2_X1 U6241 ( .A1(n5981), .A2(n14971), .ZN(n14249) );
  NOR2_X1 U6242 ( .A1(n5982), .A2(n14971), .ZN(n14252) );
  NOR2_X1 U6243 ( .A1(n5983), .A2(n14970), .ZN(n14255) );
  NOR2_X1 U6244 ( .A1(n5984), .A2(n14970), .ZN(n14258) );
  NOR2_X1 U6245 ( .A1(n5985), .A2(n14970), .ZN(n14261) );
  NOR2_X1 U6246 ( .A1(n5986), .A2(n14970), .ZN(n14264) );
  NOR2_X1 U6247 ( .A1(n5987), .A2(n14970), .ZN(n14267) );
  NOR2_X1 U6249 ( .A1(n5988), .A2(n14970), .ZN(n14270) );
  NOR2_X1 U6250 ( .A1(n5989), .A2(n14970), .ZN(n14273) );
  NOR2_X1 U6251 ( .A1(n5990), .A2(n14970), .ZN(n14276) );
  NOR2_X1 U6252 ( .A1(n5991), .A2(n14971), .ZN(n14279) );
  AOI221_X1 U6253 ( .B1(n14351), .B2(n3343), .C1(n5851), .C2(n1), .A(n1192), 
        .ZN(n1188) );
  OAI22_X1 U6254 ( .A1(n9562), .A2(n14361), .B1(n9567), .B2(n14509), .ZN(n1192) );
  AOI221_X1 U6255 ( .B1(n14351), .B2(n3345), .C1(n5851), .C2(n2), .A(n1201), 
        .ZN(n1197) );
  OAI22_X1 U6256 ( .A1(n6490), .A2(n14361), .B1(n6495), .B2(n14509), .ZN(n1201) );
  AOI221_X1 U6257 ( .B1(n14351), .B2(n3346), .C1(n5851), .C2(n3), .A(n1210), 
        .ZN(n1206) );
  OAI22_X1 U6258 ( .A1(n7514), .A2(n14361), .B1(n7519), .B2(n14509), .ZN(n1210) );
  AOI221_X1 U6259 ( .B1(n14350), .B2(n3354), .C1(n5799), .C2(n4), .A(n1355), 
        .ZN(n1352) );
  OAI22_X1 U6260 ( .A1(n9546), .A2(n14362), .B1(n9551), .B2(n14510), .ZN(n1355) );
  AOI221_X1 U6261 ( .B1(n14349), .B2(n3355), .C1(n5799), .C2(n5), .A(n1363), 
        .ZN(n1360) );
  OAI22_X1 U6262 ( .A1(n6474), .A2(n14362), .B1(n6479), .B2(n14510), .ZN(n1363) );
  AOI221_X1 U6263 ( .B1(n14349), .B2(n3357), .C1(n5799), .C2(n6), .A(n1371), 
        .ZN(n1368) );
  OAI22_X1 U6264 ( .A1(n7498), .A2(n14362), .B1(n7503), .B2(n14510), .ZN(n1371) );
  AOI221_X1 U6265 ( .B1(n14348), .B2(n3358), .C1(n5815), .C2(n7), .A(n1504), 
        .ZN(n1501) );
  OAI22_X1 U6266 ( .A1(n9530), .A2(n14363), .B1(n9535), .B2(n14511), .ZN(n1504) );
  AOI221_X1 U6267 ( .B1(n14348), .B2(n3362), .C1(n5815), .C2(n8), .A(n1512), 
        .ZN(n1509) );
  OAI22_X1 U6268 ( .A1(n6458), .A2(n14363), .B1(n6463), .B2(n14511), .ZN(n1512) );
  AOI221_X1 U6269 ( .B1(n14348), .B2(n3363), .C1(n5815), .C2(n9), .A(n1520), 
        .ZN(n1517) );
  OAI22_X1 U6270 ( .A1(n7482), .A2(n14363), .B1(n7487), .B2(n14511), .ZN(n1520) );
  AOI221_X1 U6271 ( .B1(n14347), .B2(n3365), .C1(n5816), .C2(n10), .A(n1653), 
        .ZN(n1650) );
  OAI22_X1 U6272 ( .A1(n9514), .A2(n14364), .B1(n9519), .B2(n14512), .ZN(n1653) );
  AOI221_X1 U6273 ( .B1(n14347), .B2(n3366), .C1(n5816), .C2(n11), .A(n1661), 
        .ZN(n1658) );
  OAI22_X1 U6274 ( .A1(n6442), .A2(n14365), .B1(n6447), .B2(n14513), .ZN(n1661) );
  AOI221_X1 U6275 ( .B1(n14347), .B2(n3370), .C1(n5816), .C2(n12), .A(n1669), 
        .ZN(n1666) );
  OAI22_X1 U6276 ( .A1(n7466), .A2(n14365), .B1(n7471), .B2(n14513), .ZN(n1669) );
  AOI221_X1 U6277 ( .B1(n14346), .B2(n3371), .C1(n5818), .C2(n13), .A(n1802), 
        .ZN(n1799) );
  OAI22_X1 U6278 ( .A1(n9498), .A2(n14366), .B1(n9503), .B2(n14514), .ZN(n1802) );
  AOI221_X1 U6279 ( .B1(n14346), .B2(n3373), .C1(n5818), .C2(n14), .A(n1810), 
        .ZN(n1807) );
  OAI22_X1 U6280 ( .A1(n6426), .A2(n14366), .B1(n6431), .B2(n14514), .ZN(n1810) );
  AOI221_X1 U6281 ( .B1(n14346), .B2(n3374), .C1(n5816), .C2(n15), .A(n1818), 
        .ZN(n1815) );
  OAI22_X1 U6282 ( .A1(n7450), .A2(n14366), .B1(n7455), .B2(n14514), .ZN(n1818) );
  AOI221_X1 U6283 ( .B1(n14345), .B2(n3378), .C1(n5818), .C2(n16), .A(n1951), 
        .ZN(n1948) );
  OAI22_X1 U6284 ( .A1(n9482), .A2(n14367), .B1(n9487), .B2(n14515), .ZN(n1951) );
  AOI221_X1 U6285 ( .B1(n14345), .B2(n3379), .C1(n5818), .C2(n17), .A(n1959), 
        .ZN(n1956) );
  OAI22_X1 U6286 ( .A1(n6410), .A2(n14367), .B1(n6415), .B2(n14515), .ZN(n1959) );
  AOI221_X1 U6287 ( .B1(n14344), .B2(n3381), .C1(n5818), .C2(n18), .A(n1967), 
        .ZN(n1964) );
  OAI22_X1 U6288 ( .A1(n7434), .A2(n14367), .B1(n7439), .B2(n14515), .ZN(n1967) );
  AOI221_X1 U6289 ( .B1(n14343), .B2(n3382), .C1(n5819), .C2(n19), .A(n2100), 
        .ZN(n2097) );
  OAI22_X1 U6290 ( .A1(n9466), .A2(n14368), .B1(n9471), .B2(n14516), .ZN(n2100) );
  AOI221_X1 U6291 ( .B1(n14343), .B2(n3390), .C1(n5824), .C2(n20), .A(n2108), 
        .ZN(n2105) );
  OAI22_X1 U6292 ( .A1(n6394), .A2(n14368), .B1(n6399), .B2(n14516), .ZN(n2108) );
  AOI221_X1 U6293 ( .B1(n14343), .B2(n3391), .C1(n5824), .C2(n21), .A(n2116), 
        .ZN(n2113) );
  OAI22_X1 U6294 ( .A1(n7418), .A2(n14368), .B1(n7423), .B2(n14516), .ZN(n2116) );
  AOI221_X1 U6295 ( .B1(n14342), .B2(n3393), .C1(n5826), .C2(n22), .A(n2249), 
        .ZN(n2246) );
  OAI22_X1 U6296 ( .A1(n9450), .A2(n14369), .B1(n9455), .B2(n14517), .ZN(n2249) );
  AOI221_X1 U6297 ( .B1(n14342), .B2(n3394), .C1(n5826), .C2(n23), .A(n2257), 
        .ZN(n2254) );
  OAI22_X1 U6298 ( .A1(n6378), .A2(n14369), .B1(n6383), .B2(n14517), .ZN(n2257) );
  AOI221_X1 U6299 ( .B1(n14342), .B2(n3398), .C1(n5826), .C2(n24), .A(n2265), 
        .ZN(n2262) );
  OAI22_X1 U6300 ( .A1(n7402), .A2(n14370), .B1(n7407), .B2(n14518), .ZN(n2265) );
  AOI221_X1 U6301 ( .B1(n14341), .B2(n3399), .C1(n5826), .C2(n25), .A(n2398), 
        .ZN(n2395) );
  OAI22_X1 U6302 ( .A1(n9434), .A2(n14371), .B1(n9439), .B2(n14519), .ZN(n2398) );
  AOI221_X1 U6303 ( .B1(n14341), .B2(n3401), .C1(n5827), .C2(n26), .A(n2406), 
        .ZN(n2403) );
  OAI22_X1 U6304 ( .A1(n6362), .A2(n14371), .B1(n6367), .B2(n14519), .ZN(n2406) );
  AOI221_X1 U6305 ( .B1(n14341), .B2(n3402), .C1(n5851), .C2(n27), .A(n2414), 
        .ZN(n2411) );
  OAI22_X1 U6306 ( .A1(n7386), .A2(n14371), .B1(n7391), .B2(n14519), .ZN(n2414) );
  AOI221_X1 U6307 ( .B1(n14340), .B2(n3406), .C1(n5832), .C2(n28), .A(n2547), 
        .ZN(n2544) );
  OAI22_X1 U6308 ( .A1(n9418), .A2(n14372), .B1(n9423), .B2(n14520), .ZN(n2547) );
  AOI221_X1 U6309 ( .B1(n14340), .B2(n3407), .C1(n5827), .C2(n29), .A(n2555), 
        .ZN(n2552) );
  OAI22_X1 U6310 ( .A1(n6346), .A2(n14372), .B1(n6351), .B2(n14520), .ZN(n2555) );
  AOI221_X1 U6311 ( .B1(n14340), .B2(n3409), .C1(n5831), .C2(n30), .A(n2563), 
        .ZN(n2560) );
  OAI22_X1 U6312 ( .A1(n7370), .A2(n14372), .B1(n7375), .B2(n14520), .ZN(n2563) );
  AOI221_X1 U6313 ( .B1(n14338), .B2(n3410), .C1(n5832), .C2(n31), .A(n2696), 
        .ZN(n2693) );
  OAI22_X1 U6314 ( .A1(n9402), .A2(n14373), .B1(n9407), .B2(n14521), .ZN(n2696) );
  AOI221_X1 U6315 ( .B1(n14338), .B2(n3414), .C1(n5832), .C2(n32), .A(n2704), 
        .ZN(n2701) );
  OAI22_X1 U6316 ( .A1(n6330), .A2(n14373), .B1(n6335), .B2(n14521), .ZN(n2704) );
  AOI221_X1 U6317 ( .B1(n14338), .B2(n3415), .C1(n5832), .C2(n33), .A(n2712), 
        .ZN(n2709) );
  OAI22_X1 U6318 ( .A1(n7354), .A2(n14373), .B1(n7359), .B2(n14521), .ZN(n2712) );
  AOI221_X1 U6319 ( .B1(n14337), .B2(n3417), .C1(n5834), .C2(n34), .A(n2845), 
        .ZN(n2842) );
  OAI22_X1 U6320 ( .A1(n9386), .A2(n14374), .B1(n9391), .B2(n14522), .ZN(n2845) );
  AOI221_X1 U6321 ( .B1(n14337), .B2(n3418), .C1(n5834), .C2(n35), .A(n2853), 
        .ZN(n2850) );
  OAI22_X1 U6322 ( .A1(n6314), .A2(n14374), .B1(n6319), .B2(n14522), .ZN(n2853) );
  AOI221_X1 U6323 ( .B1(n14337), .B2(n3431), .C1(n5834), .C2(n36), .A(n2861), 
        .ZN(n2858) );
  OAI22_X1 U6324 ( .A1(n7338), .A2(n14374), .B1(n7343), .B2(n14522), .ZN(n2861) );
  AOI221_X1 U6325 ( .B1(n14336), .B2(n3432), .C1(n5835), .C2(n37), .A(n2994), 
        .ZN(n2991) );
  OAI22_X1 U6326 ( .A1(n9370), .A2(n14376), .B1(n9375), .B2(n14524), .ZN(n2994) );
  AOI221_X1 U6327 ( .B1(n14336), .B2(n3434), .C1(n5835), .C2(n38), .A(n3002), 
        .ZN(n2999) );
  OAI22_X1 U6328 ( .A1(n6298), .A2(n14376), .B1(n6303), .B2(n14524), .ZN(n3002) );
  AOI221_X1 U6329 ( .B1(n14336), .B2(n3435), .C1(n5835), .C2(n39), .A(n3010), 
        .ZN(n3007) );
  OAI22_X1 U6330 ( .A1(n7322), .A2(n14376), .B1(n7327), .B2(n14524), .ZN(n3010) );
  AOI221_X1 U6331 ( .B1(n14335), .B2(n3439), .C1(n5839), .C2(n40), .A(n3143), 
        .ZN(n3140) );
  OAI22_X1 U6332 ( .A1(n9354), .A2(n14377), .B1(n9359), .B2(n14525), .ZN(n3143) );
  AOI221_X1 U6333 ( .B1(n14335), .B2(n3440), .C1(n5842), .C2(n41), .A(n3151), 
        .ZN(n3148) );
  OAI22_X1 U6334 ( .A1(n6282), .A2(n14377), .B1(n6287), .B2(n14525), .ZN(n3151) );
  AOI221_X1 U6335 ( .B1(n14335), .B2(n3442), .C1(n5842), .C2(n42), .A(n3159), 
        .ZN(n3156) );
  OAI22_X1 U6336 ( .A1(n7306), .A2(n14377), .B1(n7311), .B2(n14525), .ZN(n3159) );
  AOI221_X1 U6337 ( .B1(n14334), .B2(n3443), .C1(n5843), .C2(n43), .A(n3292), 
        .ZN(n3289) );
  OAI22_X1 U6338 ( .A1(n9338), .A2(n14378), .B1(n9343), .B2(n14526), .ZN(n3292) );
  AOI221_X1 U6339 ( .B1(n14333), .B2(n3447), .C1(n5842), .C2(n44), .A(n3300), 
        .ZN(n3297) );
  OAI22_X1 U6340 ( .A1(n6266), .A2(n14378), .B1(n6271), .B2(n14526), .ZN(n3300) );
  AOI221_X1 U6341 ( .B1(n14333), .B2(n3448), .C1(n5842), .C2(n45), .A(n3308), 
        .ZN(n3305) );
  OAI22_X1 U6342 ( .A1(n7290), .A2(n14378), .B1(n7295), .B2(n14526), .ZN(n3308) );
  AOI221_X1 U6343 ( .B1(n14332), .B2(n3450), .C1(n5843), .C2(n46), .A(n3441), 
        .ZN(n3438) );
  OAI22_X1 U6344 ( .A1(n9322), .A2(n14379), .B1(n9327), .B2(n14527), .ZN(n3441) );
  AOI221_X1 U6345 ( .B1(n14332), .B2(n3451), .C1(n5843), .C2(n47), .A(n3449), 
        .ZN(n3446) );
  OAI22_X1 U6346 ( .A1(n6250), .A2(n14379), .B1(n6255), .B2(n14527), .ZN(n3449) );
  AOI221_X1 U6347 ( .B1(n14332), .B2(n3455), .C1(n5843), .C2(n48), .A(n3457), 
        .ZN(n3454) );
  OAI22_X1 U6348 ( .A1(n7274), .A2(n14379), .B1(n7279), .B2(n14527), .ZN(n3457) );
  AOI221_X1 U6349 ( .B1(n14331), .B2(n3456), .C1(n5852), .C2(n49), .A(n3590), 
        .ZN(n3587) );
  OAI22_X1 U6350 ( .A1(n9306), .A2(n14380), .B1(n9311), .B2(n14528), .ZN(n3590) );
  AOI221_X1 U6351 ( .B1(n14331), .B2(n3458), .C1(n5852), .C2(n50), .A(n3598), 
        .ZN(n3595) );
  OAI22_X1 U6352 ( .A1(n6234), .A2(n14381), .B1(n6239), .B2(n14529), .ZN(n3598) );
  AOI221_X1 U6353 ( .B1(n14331), .B2(n3459), .C1(n5852), .C2(n51), .A(n3606), 
        .ZN(n3603) );
  OAI22_X1 U6354 ( .A1(n7258), .A2(n14381), .B1(n7263), .B2(n14529), .ZN(n3606) );
  AOI221_X1 U6355 ( .B1(n14330), .B2(n3467), .C1(n5854), .C2(n52), .A(n3739), 
        .ZN(n3736) );
  OAI22_X1 U6356 ( .A1(n9290), .A2(n14382), .B1(n9295), .B2(n14530), .ZN(n3739) );
  AOI221_X1 U6357 ( .B1(n14330), .B2(n3468), .C1(n5854), .C2(n53), .A(n3747), 
        .ZN(n3744) );
  OAI22_X1 U6358 ( .A1(n6218), .A2(n14382), .B1(n6223), .B2(n14530), .ZN(n3747) );
  AOI221_X1 U6359 ( .B1(n14330), .B2(n3470), .C1(n5852), .C2(n54), .A(n3755), 
        .ZN(n3752) );
  OAI22_X1 U6360 ( .A1(n7242), .A2(n14382), .B1(n7247), .B2(n14530), .ZN(n3755) );
  AOI221_X1 U6361 ( .B1(n14329), .B2(n3471), .C1(n5854), .C2(n55), .A(n3888), 
        .ZN(n3885) );
  OAI22_X1 U6362 ( .A1(n9274), .A2(n14383), .B1(n9279), .B2(n14531), .ZN(n3888) );
  AOI221_X1 U6363 ( .B1(n14329), .B2(n3475), .C1(n5854), .C2(n56), .A(n3896), 
        .ZN(n3893) );
  OAI22_X1 U6364 ( .A1(n6202), .A2(n14383), .B1(n6207), .B2(n14531), .ZN(n3896) );
  AOI221_X1 U6365 ( .B1(n14328), .B2(n3476), .C1(n5854), .C2(n57), .A(n3904), 
        .ZN(n3901) );
  OAI22_X1 U6366 ( .A1(n7226), .A2(n14383), .B1(n7231), .B2(n14531), .ZN(n3904) );
  AOI221_X1 U6367 ( .B1(n14327), .B2(n3478), .C1(n5855), .C2(n58), .A(n4037), 
        .ZN(n4034) );
  OAI22_X1 U6368 ( .A1(n9258), .A2(n14384), .B1(n9263), .B2(n14532), .ZN(n4037) );
  AOI221_X1 U6369 ( .B1(n14327), .B2(n3479), .C1(n5860), .C2(n59), .A(n4045), 
        .ZN(n4042) );
  OAI22_X1 U6370 ( .A1(n6186), .A2(n14384), .B1(n6191), .B2(n14532), .ZN(n4045) );
  AOI221_X1 U6371 ( .B1(n14327), .B2(n3483), .C1(n5860), .C2(n60), .A(n4053), 
        .ZN(n4050) );
  OAI22_X1 U6372 ( .A1(n7210), .A2(n14384), .B1(n7215), .B2(n14532), .ZN(n4053) );
  AOI221_X1 U6373 ( .B1(n14326), .B2(n3484), .C1(n5862), .C2(n61), .A(n4186), 
        .ZN(n4183) );
  OAI22_X1 U6374 ( .A1(n9242), .A2(n14385), .B1(n9247), .B2(n14533), .ZN(n4186) );
  AOI221_X1 U6375 ( .B1(n14326), .B2(n3486), .C1(n5862), .C2(n62), .A(n4194), 
        .ZN(n4191) );
  OAI22_X1 U6376 ( .A1(n6170), .A2(n14385), .B1(n6175), .B2(n14533), .ZN(n4194) );
  AOI221_X1 U6377 ( .B1(n14326), .B2(n3487), .C1(n5862), .C2(n63), .A(n4202), 
        .ZN(n4199) );
  OAI22_X1 U6378 ( .A1(n7194), .A2(n14386), .B1(n7199), .B2(n14534), .ZN(n4202) );
  AOI221_X1 U6379 ( .B1(n14325), .B2(n3491), .C1(n5863), .C2(n64), .A(n4335), 
        .ZN(n4332) );
  OAI22_X1 U6380 ( .A1(n9226), .A2(n14387), .B1(n9231), .B2(n14535), .ZN(n4335) );
  AOI221_X1 U6381 ( .B1(n14325), .B2(n3492), .C1(n5863), .C2(n65), .A(n4343), 
        .ZN(n4340) );
  OAI22_X1 U6382 ( .A1(n6154), .A2(n14387), .B1(n6159), .B2(n14535), .ZN(n4343) );
  AOI221_X1 U6383 ( .B1(n14325), .B2(n3494), .C1(n5863), .C2(n76), .A(n4351), 
        .ZN(n4348) );
  OAI22_X1 U6384 ( .A1(n7178), .A2(n14387), .B1(n7183), .B2(n14535), .ZN(n4351) );
  AOI221_X1 U6385 ( .B1(n14324), .B2(n3495), .C1(n5863), .C2(n80), .A(n4484), 
        .ZN(n4481) );
  OAI22_X1 U6386 ( .A1(n9210), .A2(n14388), .B1(n9215), .B2(n14536), .ZN(n4484) );
  AOI221_X1 U6387 ( .B1(n14324), .B2(n3503), .C1(n5863), .C2(n83), .A(n4492), 
        .ZN(n4489) );
  OAI22_X1 U6388 ( .A1(n6138), .A2(n14388), .B1(n6143), .B2(n14536), .ZN(n4492) );
  AOI221_X1 U6389 ( .B1(n14324), .B2(n3504), .C1(n5863), .C2(n86), .A(n4500), 
        .ZN(n4497) );
  OAI22_X1 U6390 ( .A1(n7162), .A2(n14388), .B1(n7167), .B2(n14536), .ZN(n4500) );
  AOI221_X1 U6391 ( .B1(n14322), .B2(n3506), .C1(n5867), .C2(n89), .A(n4633), 
        .ZN(n4630) );
  OAI22_X1 U6392 ( .A1(n9194), .A2(n14389), .B1(n9199), .B2(n14537), .ZN(n4633) );
  AOI221_X1 U6393 ( .B1(n14322), .B2(n3507), .C1(n5799), .C2(n92), .A(n4641), 
        .ZN(n4638) );
  OAI22_X1 U6394 ( .A1(n6122), .A2(n14389), .B1(n6127), .B2(n14537), .ZN(n4641) );
  AOI221_X1 U6395 ( .B1(n14322), .B2(n3511), .C1(n5870), .C2(n95), .A(n4649), 
        .ZN(n4646) );
  OAI22_X1 U6396 ( .A1(n7146), .A2(n14389), .B1(n7151), .B2(n14537), .ZN(n4649) );
  AOI221_X1 U6397 ( .B1(n14321), .B2(n3512), .C1(n5870), .C2(n98), .A(n4782), 
        .ZN(n4779) );
  OAI22_X1 U6398 ( .A1(n9178), .A2(n14390), .B1(n9183), .B2(n14538), .ZN(n4782) );
  AOI221_X1 U6399 ( .B1(n14321), .B2(n3514), .C1(n5870), .C2(n101), .A(n4790), 
        .ZN(n4787) );
  OAI22_X1 U6401 ( .A1(n6106), .A2(n14390), .B1(n6111), .B2(n14538), .ZN(n4790) );
  AOI221_X1 U6402 ( .B1(n14321), .B2(n3515), .C1(n5879), .C2(n104), .A(n4798), 
        .ZN(n4795) );
  OAI22_X1 U6403 ( .A1(n7130), .A2(n14390), .B1(n7135), .B2(n14538), .ZN(n4798) );
  AOI221_X1 U6404 ( .B1(n14320), .B2(n3519), .C1(n5871), .C2(n107), .A(n4931), 
        .ZN(n4928) );
  OAI22_X1 U6405 ( .A1(n9162), .A2(n14392), .B1(n9167), .B2(n14540), .ZN(n4931) );
  AOI221_X1 U6406 ( .B1(n14320), .B2(n3520), .C1(n5871), .C2(n110), .A(n4939), 
        .ZN(n4936) );
  OAI22_X1 U6407 ( .A1(n6090), .A2(n14392), .B1(n6095), .B2(n14540), .ZN(n4939) );
  AOI221_X1 U6408 ( .B1(n14320), .B2(n3522), .C1(n5871), .C2(n113), .A(n4947), 
        .ZN(n4944) );
  OAI22_X1 U6409 ( .A1(n7114), .A2(n14392), .B1(n7119), .B2(n14540), .ZN(n4947) );
  AOI221_X1 U6410 ( .B1(n14319), .B2(n3523), .C1(n5875), .C2(n116), .A(n5080), 
        .ZN(n5077) );
  OAI22_X1 U6411 ( .A1(n9146), .A2(n14393), .B1(n9151), .B2(n14541), .ZN(n5080) );
  AOI221_X1 U6412 ( .B1(n14319), .B2(n3527), .C1(n5878), .C2(n119), .A(n5088), 
        .ZN(n5085) );
  OAI22_X1 U6413 ( .A1(n6074), .A2(n14393), .B1(n6079), .B2(n14541), .ZN(n5088) );
  AOI221_X1 U6414 ( .B1(n14319), .B2(n3528), .C1(n5878), .C2(n122), .A(n5096), 
        .ZN(n5093) );
  OAI22_X1 U6415 ( .A1(n7098), .A2(n14393), .B1(n7103), .B2(n14541), .ZN(n5096) );
  AOI221_X1 U6416 ( .B1(n14318), .B2(n3530), .C1(n5879), .C2(n125), .A(n5229), 
        .ZN(n5226) );
  OAI22_X1 U6417 ( .A1(n9130), .A2(n14394), .B1(n9135), .B2(n14542), .ZN(n5229) );
  AOI221_X1 U6418 ( .B1(n14317), .B2(n3531), .C1(n5878), .C2(n128), .A(n5237), 
        .ZN(n5234) );
  OAI22_X1 U6419 ( .A1(n6058), .A2(n14394), .B1(n6063), .B2(n14542), .ZN(n5237) );
  AOI221_X1 U6420 ( .B1(n14317), .B2(n3539), .C1(n5878), .C2(n131), .A(n5245), 
        .ZN(n5242) );
  OAI22_X1 U6421 ( .A1(n7082), .A2(n14394), .B1(n7087), .B2(n14542), .ZN(n5245) );
  AOI221_X1 U6422 ( .B1(n14316), .B2(n3540), .C1(n5879), .C2(n134), .A(n5378), 
        .ZN(n5375) );
  OAI22_X1 U6423 ( .A1(n9114), .A2(n14395), .B1(n9119), .B2(n14543), .ZN(n5378) );
  AOI221_X1 U6424 ( .B1(n14316), .B2(n3542), .C1(n5879), .C2(n137), .A(n5386), 
        .ZN(n5383) );
  OAI22_X1 U6425 ( .A1(n6042), .A2(n14395), .B1(n6047), .B2(n14543), .ZN(n5386) );
  AOI221_X1 U6426 ( .B1(n14316), .B2(n3543), .C1(n5879), .C2(n140), .A(n5394), 
        .ZN(n5391) );
  OAI22_X1 U6427 ( .A1(n7066), .A2(n14395), .B1(n7071), .B2(n14543), .ZN(n5394) );
  AOI221_X1 U6428 ( .B1(n14315), .B2(n3547), .C1(n5889), .C2(n143), .A(n5527), 
        .ZN(n5524) );
  OAI22_X1 U6429 ( .A1(n9098), .A2(n14396), .B1(n9103), .B2(n14544), .ZN(n5527) );
  AOI221_X1 U6430 ( .B1(n14315), .B2(n3548), .C1(n5889), .C2(n146), .A(n5535), 
        .ZN(n5532) );
  OAI22_X1 U6431 ( .A1(n6026), .A2(n14397), .B1(n6031), .B2(n14545), .ZN(n5535) );
  AOI221_X1 U6432 ( .B1(n14315), .B2(n3550), .C1(n5889), .C2(n149), .A(n5543), 
        .ZN(n5540) );
  OAI22_X1 U6433 ( .A1(n7050), .A2(n14397), .B1(n7055), .B2(n14545), .ZN(n5543) );
  AOI221_X1 U6434 ( .B1(n14314), .B2(n3551), .C1(n5890), .C2(n152), .A(n5676), 
        .ZN(n5673) );
  OAI22_X1 U6435 ( .A1(n9082), .A2(n14398), .B1(n9087), .B2(n14546), .ZN(n5676) );
  AOI221_X1 U6436 ( .B1(n14314), .B2(n3555), .C1(n5893), .C2(n155), .A(n5684), 
        .ZN(n5681) );
  OAI22_X1 U6437 ( .A1(n6010), .A2(n14398), .B1(n6015), .B2(n14546), .ZN(n5684) );
  AOI221_X1 U6438 ( .B1(n14314), .B2(n3556), .C1(n5893), .C2(n158), .A(n5692), 
        .ZN(n5689) );
  OAI22_X1 U6439 ( .A1(n7034), .A2(n14398), .B1(n7039), .B2(n14546), .ZN(n5692) );
  AOI221_X1 U6440 ( .B1(n14313), .B2(n3558), .C1(n5897), .C2(n161), .A(n5817), 
        .ZN(n5814) );
  OAI22_X1 U6441 ( .A1(n8042), .A2(n14399), .B1(n8047), .B2(n14547), .ZN(n5817) );
  AOI221_X1 U6442 ( .B1(n14313), .B2(n3559), .C1(n5897), .C2(n164), .A(n5825), 
        .ZN(n5822) );
  OAI22_X1 U6443 ( .A1(n9066), .A2(n14399), .B1(n9071), .B2(n14547), .ZN(n5825) );
  AOI221_X1 U6444 ( .B1(n14313), .B2(n3563), .C1(n5897), .C2(n167), .A(n5833), 
        .ZN(n5830) );
  OAI22_X1 U6445 ( .A1(n5994), .A2(n14399), .B1(n5999), .B2(n14547), .ZN(n5833) );
  AOI221_X1 U6446 ( .B1(n14450), .B2(n3564), .C1(n14493), .C2(n170), .A(n1195), 
        .ZN(n1187) );
  OAI22_X1 U6447 ( .A1(n9563), .A2(n14553), .B1(n9561), .B2(n14635), .ZN(n1195) );
  AOI221_X1 U6448 ( .B1(n14450), .B2(n3566), .C1(n14493), .C2(n172), .A(n1204), 
        .ZN(n1196) );
  OAI22_X1 U6449 ( .A1(n6491), .A2(n14553), .B1(n6489), .B2(n14635), .ZN(n1204) );
  AOI221_X1 U6450 ( .B1(n14450), .B2(n3567), .C1(n14493), .C2(n238), .A(n1213), 
        .ZN(n1205) );
  OAI22_X1 U6451 ( .A1(n7515), .A2(n14553), .B1(n7513), .B2(n14635), .ZN(n1213) );
  AOI221_X1 U6452 ( .B1(n14449), .B2(n3580), .C1(n14492), .C2(n1181), .A(n1358), .ZN(n1351) );
  OAI22_X1 U6453 ( .A1(n9547), .A2(n14554), .B1(n9545), .B2(n14634), .ZN(n1358) );
  AOI221_X1 U6454 ( .B1(n14448), .B2(n3581), .C1(n14491), .C2(n1182), .A(n1366), .ZN(n1359) );
  OAI22_X1 U6455 ( .A1(n6475), .A2(n14554), .B1(n6473), .B2(n14634), .ZN(n1366) );
  AOI221_X1 U6456 ( .B1(n14448), .B2(n3583), .C1(n14491), .C2(n1184), .A(n1374), .ZN(n1367) );
  OAI22_X1 U6457 ( .A1(n7499), .A2(n14554), .B1(n7497), .B2(n14634), .ZN(n1374) );
  AOI221_X1 U6458 ( .B1(n14447), .B2(n3584), .C1(n14490), .C2(n1185), .A(n1507), .ZN(n1500) );
  OAI22_X1 U6459 ( .A1(n9531), .A2(n14555), .B1(n9529), .B2(n14633), .ZN(n1507) );
  AOI221_X1 U6460 ( .B1(n14447), .B2(n3588), .C1(n14490), .C2(n1190), .A(n1515), .ZN(n1508) );
  OAI22_X1 U6461 ( .A1(n6459), .A2(n14555), .B1(n6457), .B2(n14633), .ZN(n1515) );
  AOI221_X1 U6462 ( .B1(n14447), .B2(n3589), .C1(n14490), .C2(n1191), .A(n1523), .ZN(n1516) );
  OAI22_X1 U6463 ( .A1(n7483), .A2(n14555), .B1(n7481), .B2(n14633), .ZN(n1523) );
  AOI221_X1 U6464 ( .B1(n14446), .B2(n3591), .C1(n14489), .C2(n1193), .A(n1656), .ZN(n1649) );
  OAI22_X1 U6465 ( .A1(n9515), .A2(n14556), .B1(n9513), .B2(n14632), .ZN(n1656) );
  AOI221_X1 U6466 ( .B1(n14446), .B2(n3592), .C1(n14489), .C2(n1194), .A(n1664), .ZN(n1657) );
  OAI22_X1 U6467 ( .A1(n6443), .A2(n14557), .B1(n6441), .B2(n14631), .ZN(n1664) );
  AOI221_X1 U6468 ( .B1(n14446), .B2(n3596), .C1(n14489), .C2(n1199), .A(n1672), .ZN(n1665) );
  OAI22_X1 U6469 ( .A1(n7467), .A2(n14557), .B1(n7465), .B2(n14631), .ZN(n1672) );
  AOI221_X1 U6470 ( .B1(n14445), .B2(n3597), .C1(n14488), .C2(n1200), .A(n1805), .ZN(n1798) );
  OAI22_X1 U6471 ( .A1(n9499), .A2(n14558), .B1(n9497), .B2(n14630), .ZN(n1805) );
  AOI221_X1 U6472 ( .B1(n14445), .B2(n3599), .C1(n14488), .C2(n1202), .A(n1813), .ZN(n1806) );
  OAI22_X1 U6473 ( .A1(n6427), .A2(n14558), .B1(n6425), .B2(n14630), .ZN(n1813) );
  AOI221_X1 U6474 ( .B1(n14445), .B2(n3600), .C1(n14488), .C2(n1203), .A(n1821), .ZN(n1814) );
  OAI22_X1 U6475 ( .A1(n7451), .A2(n14558), .B1(n7449), .B2(n14630), .ZN(n1821) );
  AOI221_X1 U6476 ( .B1(n14444), .B2(n3604), .C1(n14487), .C2(n1208), .A(n1954), .ZN(n1947) );
  OAI22_X1 U6477 ( .A1(n9483), .A2(n14559), .B1(n9481), .B2(n14629), .ZN(n1954) );
  AOI221_X1 U6478 ( .B1(n14444), .B2(n3605), .C1(n14487), .C2(n1209), .A(n1962), .ZN(n1955) );
  OAI22_X1 U6479 ( .A1(n6411), .A2(n14559), .B1(n6409), .B2(n14629), .ZN(n1962) );
  AOI221_X1 U6480 ( .B1(n14443), .B2(n3607), .C1(n14486), .C2(n1211), .A(n1970), .ZN(n1963) );
  OAI22_X1 U6481 ( .A1(n7435), .A2(n14559), .B1(n7433), .B2(n14629), .ZN(n1970) );
  AOI221_X1 U6482 ( .B1(n14442), .B2(n3608), .C1(n14485), .C2(n1212), .A(n2103), .ZN(n2096) );
  OAI22_X1 U6483 ( .A1(n9467), .A2(n14560), .B1(n9465), .B2(n14628), .ZN(n2103) );
  AOI221_X1 U6484 ( .B1(n14442), .B2(n3616), .C1(n14485), .C2(n1221), .A(n2111), .ZN(n2104) );
  OAI22_X1 U6485 ( .A1(n6395), .A2(n14560), .B1(n6393), .B2(n14628), .ZN(n2111) );
  AOI221_X1 U6486 ( .B1(n14442), .B2(n3617), .C1(n14485), .C2(n1222), .A(n2119), .ZN(n2112) );
  OAI22_X1 U6487 ( .A1(n7419), .A2(n14560), .B1(n7417), .B2(n14628), .ZN(n2119) );
  AOI221_X1 U6488 ( .B1(n14441), .B2(n3619), .C1(n14484), .C2(n1224), .A(n2252), .ZN(n2245) );
  OAI22_X1 U6489 ( .A1(n9451), .A2(n14561), .B1(n9449), .B2(n14627), .ZN(n2252) );
  AOI221_X1 U6490 ( .B1(n14441), .B2(n3620), .C1(n14484), .C2(n1225), .A(n2260), .ZN(n2253) );
  OAI22_X1 U6491 ( .A1(n6379), .A2(n14561), .B1(n6377), .B2(n14626), .ZN(n2260) );
  AOI221_X1 U6492 ( .B1(n14441), .B2(n3624), .C1(n14484), .C2(n1230), .A(n2268), .ZN(n2261) );
  OAI22_X1 U6493 ( .A1(n7403), .A2(n14562), .B1(n7401), .B2(n14626), .ZN(n2268) );
  AOI221_X1 U6494 ( .B1(n14440), .B2(n3625), .C1(n14483), .C2(n1231), .A(n2401), .ZN(n2394) );
  OAI22_X1 U6495 ( .A1(n9435), .A2(n14563), .B1(n9433), .B2(n14645), .ZN(n2401) );
  AOI221_X1 U6496 ( .B1(n14440), .B2(n3627), .C1(n14483), .C2(n1233), .A(n2409), .ZN(n2402) );
  OAI22_X1 U6497 ( .A1(n6363), .A2(n14563), .B1(n6361), .B2(n14645), .ZN(n2409) );
  AOI221_X1 U6498 ( .B1(n14440), .B2(n3628), .C1(n14483), .C2(n1234), .A(n2417), .ZN(n2410) );
  OAI22_X1 U6499 ( .A1(n7387), .A2(n14563), .B1(n7385), .B2(n14645), .ZN(n2417) );
  AOI221_X1 U6500 ( .B1(n14439), .B2(n3632), .C1(n14482), .C2(n1239), .A(n2550), .ZN(n2543) );
  OAI22_X1 U6501 ( .A1(n9419), .A2(n14564), .B1(n9417), .B2(n14644), .ZN(n2550) );
  AOI221_X1 U6502 ( .B1(n14439), .B2(n3633), .C1(n14482), .C2(n1240), .A(n2558), .ZN(n2551) );
  OAI22_X1 U6503 ( .A1(n6347), .A2(n14564), .B1(n6345), .B2(n14644), .ZN(n2558) );
  AOI221_X1 U6504 ( .B1(n14439), .B2(n3635), .C1(n14482), .C2(n1242), .A(n2566), .ZN(n2559) );
  OAI22_X1 U6505 ( .A1(n7371), .A2(n14564), .B1(n7369), .B2(n14644), .ZN(n2566) );
  AOI221_X1 U6506 ( .B1(n14437), .B2(n3636), .C1(n14480), .C2(n1243), .A(n2699), .ZN(n2692) );
  OAI22_X1 U6507 ( .A1(n9403), .A2(n14565), .B1(n9401), .B2(n14643), .ZN(n2699) );
  AOI221_X1 U6508 ( .B1(n14437), .B2(n3640), .C1(n14480), .C2(n1248), .A(n2707), .ZN(n2700) );
  OAI22_X1 U6509 ( .A1(n6331), .A2(n14565), .B1(n6329), .B2(n14642), .ZN(n2707) );
  AOI221_X1 U6510 ( .B1(n14437), .B2(n3641), .C1(n14480), .C2(n1249), .A(n2715), .ZN(n2708) );
  OAI22_X1 U6511 ( .A1(n7355), .A2(n14565), .B1(n7353), .B2(n14642), .ZN(n2715) );
  AOI221_X1 U6512 ( .B1(n14436), .B2(n3643), .C1(n14479), .C2(n1251), .A(n2848), .ZN(n2841) );
  OAI22_X1 U6513 ( .A1(n9387), .A2(n14566), .B1(n9385), .B2(n14641), .ZN(n2848) );
  AOI221_X1 U6514 ( .B1(n14436), .B2(n3644), .C1(n14479), .C2(n1252), .A(n2856), .ZN(n2849) );
  OAI22_X1 U6515 ( .A1(n6315), .A2(n14566), .B1(n6313), .B2(n14641), .ZN(n2856) );
  AOI221_X1 U6516 ( .B1(n14436), .B2(n3652), .C1(n14479), .C2(n1261), .A(n2864), .ZN(n2857) );
  OAI22_X1 U6517 ( .A1(n7339), .A2(n14566), .B1(n7337), .B2(n14641), .ZN(n2864) );
  AOI221_X1 U6518 ( .B1(n14435), .B2(n3653), .C1(n14478), .C2(n1262), .A(n2997), .ZN(n2990) );
  OAI22_X1 U6519 ( .A1(n9371), .A2(n14568), .B1(n9369), .B2(n14640), .ZN(n2997) );
  AOI221_X1 U6520 ( .B1(n14435), .B2(n3655), .C1(n14478), .C2(n1264), .A(n3005), .ZN(n2998) );
  OAI22_X1 U6521 ( .A1(n6299), .A2(n14568), .B1(n6297), .B2(n14640), .ZN(n3005) );
  AOI221_X1 U6522 ( .B1(n14435), .B2(n3656), .C1(n14478), .C2(n1265), .A(n3013), .ZN(n3006) );
  OAI22_X1 U6523 ( .A1(n7323), .A2(n14568), .B1(n7321), .B2(n14640), .ZN(n3013) );
  AOI221_X1 U6524 ( .B1(n14434), .B2(n3660), .C1(n14477), .C2(n1270), .A(n3146), .ZN(n3139) );
  OAI22_X1 U6525 ( .A1(n9355), .A2(n14569), .B1(n9353), .B2(n14639), .ZN(n3146) );
  AOI221_X1 U6526 ( .B1(n14434), .B2(n3661), .C1(n14477), .C2(n1271), .A(n3154), .ZN(n3147) );
  OAI22_X1 U6527 ( .A1(n6283), .A2(n14569), .B1(n6281), .B2(n14639), .ZN(n3154) );
  AOI221_X1 U6528 ( .B1(n14434), .B2(n3663), .C1(n14477), .C2(n1273), .A(n3162), .ZN(n3155) );
  OAI22_X1 U6529 ( .A1(n7307), .A2(n14569), .B1(n7305), .B2(n14639), .ZN(n3162) );
  AOI221_X1 U6530 ( .B1(n14433), .B2(n3664), .C1(n14476), .C2(n1274), .A(n3295), .ZN(n3288) );
  OAI22_X1 U6531 ( .A1(n9339), .A2(n14570), .B1(n9337), .B2(n14638), .ZN(n3295) );
  AOI221_X1 U6532 ( .B1(n14432), .B2(n3668), .C1(n14475), .C2(n1279), .A(n3303), .ZN(n3296) );
  OAI22_X1 U6533 ( .A1(n6267), .A2(n14570), .B1(n6265), .B2(n14637), .ZN(n3303) );
  AOI221_X1 U6534 ( .B1(n14432), .B2(n3669), .C1(n14475), .C2(n1280), .A(n3311), .ZN(n3304) );
  OAI22_X1 U6535 ( .A1(n7291), .A2(n14570), .B1(n7289), .B2(n14637), .ZN(n3311) );
  AOI221_X1 U6536 ( .B1(n14431), .B2(n3671), .C1(n14474), .C2(n1282), .A(n3444), .ZN(n3437) );
  OAI22_X1 U6537 ( .A1(n9323), .A2(n14571), .B1(n9321), .B2(n14636), .ZN(n3444) );
  AOI221_X1 U6538 ( .B1(n14431), .B2(n3672), .C1(n14474), .C2(n1283), .A(n3452), .ZN(n3445) );
  OAI22_X1 U6539 ( .A1(n6251), .A2(n14571), .B1(n6249), .B2(n14636), .ZN(n3452) );
  AOI221_X1 U6540 ( .B1(n14431), .B2(n3676), .C1(n14474), .C2(n1288), .A(n3460), .ZN(n3453) );
  OAI22_X1 U6541 ( .A1(n7275), .A2(n14571), .B1(n7273), .B2(n14636), .ZN(n3460) );
  AOI221_X1 U6542 ( .B1(n14430), .B2(n3677), .C1(n14473), .C2(n1289), .A(n3593), .ZN(n3586) );
  OAI22_X1 U6543 ( .A1(n9307), .A2(n14572), .B1(n9305), .B2(n14615), .ZN(n3593) );
  AOI221_X1 U6544 ( .B1(n14430), .B2(n3679), .C1(n14473), .C2(n1291), .A(n3601), .ZN(n3594) );
  OAI22_X1 U6545 ( .A1(n6235), .A2(n14573), .B1(n6233), .B2(n14615), .ZN(n3601) );
  AOI221_X1 U6546 ( .B1(n14430), .B2(n3680), .C1(n14473), .C2(n1292), .A(n3609), .ZN(n3602) );
  OAI22_X1 U6547 ( .A1(n7259), .A2(n14573), .B1(n7257), .B2(n14615), .ZN(n3609) );
  AOI221_X1 U6548 ( .B1(n14429), .B2(n3688), .C1(n14472), .C2(n1301), .A(n3742), .ZN(n3735) );
  OAI22_X1 U6549 ( .A1(n9291), .A2(n14574), .B1(n9289), .B2(n14614), .ZN(n3742) );
  AOI221_X1 U6550 ( .B1(n14429), .B2(n3689), .C1(n14472), .C2(n1302), .A(n3750), .ZN(n3743) );
  OAI22_X1 U6551 ( .A1(n6219), .A2(n14574), .B1(n6217), .B2(n14614), .ZN(n3750) );
  AOI221_X1 U6553 ( .B1(n14429), .B2(n3691), .C1(n14472), .C2(n1304), .A(n3758), .ZN(n3751) );
  OAI22_X1 U6554 ( .A1(n7243), .A2(n14574), .B1(n7241), .B2(n14614), .ZN(n3758) );
  AOI221_X1 U6555 ( .B1(n14428), .B2(n3692), .C1(n14471), .C2(n1305), .A(n3891), .ZN(n3884) );
  OAI22_X1 U6556 ( .A1(n9275), .A2(n14575), .B1(n9273), .B2(n14613), .ZN(n3891) );
  AOI221_X1 U6557 ( .B1(n14428), .B2(n3696), .C1(n14471), .C2(n1310), .A(n3899), .ZN(n3892) );
  OAI22_X1 U6558 ( .A1(n6203), .A2(n14575), .B1(n6201), .B2(n14613), .ZN(n3899) );
  AOI221_X1 U6559 ( .B1(n14427), .B2(n3697), .C1(n14470), .C2(n1311), .A(n3907), .ZN(n3900) );
  OAI22_X1 U6560 ( .A1(n7227), .A2(n14575), .B1(n7225), .B2(n14613), .ZN(n3907) );
  AOI221_X1 U6561 ( .B1(n14426), .B2(n3699), .C1(n14469), .C2(n1313), .A(n4040), .ZN(n4033) );
  OAI22_X1 U6562 ( .A1(n9259), .A2(n14576), .B1(n9257), .B2(n14612), .ZN(n4040) );
  AOI221_X1 U6563 ( .B1(n14426), .B2(n3700), .C1(n14469), .C2(n1314), .A(n4048), .ZN(n4041) );
  OAI22_X1 U6564 ( .A1(n6187), .A2(n14576), .B1(n6185), .B2(n14612), .ZN(n4048) );
  AOI221_X1 U6565 ( .B1(n14426), .B2(n3704), .C1(n14469), .C2(n1319), .A(n4056), .ZN(n4049) );
  OAI22_X1 U6566 ( .A1(n7211), .A2(n14576), .B1(n7209), .B2(n14612), .ZN(n4056) );
  AOI221_X1 U6567 ( .B1(n14425), .B2(n3705), .C1(n14468), .C2(n1320), .A(n4189), .ZN(n4182) );
  OAI22_X1 U6568 ( .A1(n9243), .A2(n14577), .B1(n9241), .B2(n14610), .ZN(n4189) );
  AOI221_X1 U6569 ( .B1(n14425), .B2(n3707), .C1(n14468), .C2(n1322), .A(n4197), .ZN(n4190) );
  OAI22_X1 U6570 ( .A1(n6171), .A2(n14577), .B1(n6169), .B2(n14610), .ZN(n4197) );
  AOI221_X1 U6571 ( .B1(n14425), .B2(n3708), .C1(n14468), .C2(n1323), .A(n4205), .ZN(n4198) );
  OAI22_X1 U6572 ( .A1(n7195), .A2(n14578), .B1(n7193), .B2(n14610), .ZN(n4205) );
  AOI221_X1 U6573 ( .B1(n14424), .B2(n3712), .C1(n14467), .C2(n1328), .A(n4338), .ZN(n4331) );
  OAI22_X1 U6574 ( .A1(n9227), .A2(n14579), .B1(n9225), .B2(n14609), .ZN(n4338) );
  AOI221_X1 U6575 ( .B1(n14424), .B2(n3713), .C1(n14467), .C2(n1329), .A(n4346), .ZN(n4339) );
  OAI22_X1 U6576 ( .A1(n6155), .A2(n14579), .B1(n6153), .B2(n14609), .ZN(n4346) );
  AOI221_X1 U6577 ( .B1(n14424), .B2(n3715), .C1(n14467), .C2(n1331), .A(n4354), .ZN(n4347) );
  OAI22_X1 U6578 ( .A1(n7179), .A2(n14579), .B1(n7177), .B2(n14609), .ZN(n4354) );
  AOI221_X1 U6579 ( .B1(n14423), .B2(n3716), .C1(n14466), .C2(n1332), .A(n4487), .ZN(n4480) );
  OAI22_X1 U6580 ( .A1(n9211), .A2(n14580), .B1(n9209), .B2(n14608), .ZN(n4487) );
  AOI221_X1 U6581 ( .B1(n14423), .B2(n3729), .C1(n14466), .C2(n1345), .A(n4495), .ZN(n4488) );
  OAI22_X1 U6582 ( .A1(n6139), .A2(n14580), .B1(n6137), .B2(n14608), .ZN(n4495) );
  AOI221_X1 U6583 ( .B1(n14423), .B2(n3730), .C1(n14466), .C2(n1346), .A(n4503), .ZN(n4496) );
  OAI22_X1 U6584 ( .A1(n7163), .A2(n14580), .B1(n7161), .B2(n14608), .ZN(n4503) );
  AOI221_X1 U6585 ( .B1(n14421), .B2(n3732), .C1(n14464), .C2(n1348), .A(n4636), .ZN(n4629) );
  OAI22_X1 U6586 ( .A1(n9195), .A2(n14581), .B1(n9193), .B2(n14607), .ZN(n4636) );
  AOI221_X1 U6587 ( .B1(n14421), .B2(n3733), .C1(n14464), .C2(n1349), .A(n4644), .ZN(n4637) );
  OAI22_X1 U6588 ( .A1(n6123), .A2(n14581), .B1(n6121), .B2(n14607), .ZN(n4644) );
  AOI221_X1 U6589 ( .B1(n14421), .B2(n3737), .C1(n14464), .C2(n1353), .A(n4652), .ZN(n4645) );
  OAI22_X1 U6590 ( .A1(n7147), .A2(n14581), .B1(n7145), .B2(n14607), .ZN(n4652) );
  AOI221_X1 U6591 ( .B1(n14420), .B2(n3738), .C1(n14463), .C2(n1354), .A(n4785), .ZN(n4778) );
  OAI22_X1 U6592 ( .A1(n9179), .A2(n14582), .B1(n9177), .B2(n14625), .ZN(n4785) );
  AOI221_X1 U6593 ( .B1(n14420), .B2(n3740), .C1(n14463), .C2(n1356), .A(n4793), .ZN(n4786) );
  OAI22_X1 U6594 ( .A1(n6107), .A2(n14582), .B1(n6105), .B2(n14625), .ZN(n4793) );
  AOI221_X1 U6595 ( .B1(n14420), .B2(n3741), .C1(n14463), .C2(n1357), .A(n4801), .ZN(n4794) );
  OAI22_X1 U6596 ( .A1(n7131), .A2(n14582), .B1(n7129), .B2(n14625), .ZN(n4801) );
  AOI221_X1 U6597 ( .B1(n14419), .B2(n3745), .C1(n14462), .C2(n1361), .A(n4934), .ZN(n4927) );
  OAI22_X1 U6598 ( .A1(n9163), .A2(n14584), .B1(n9161), .B2(n14624), .ZN(n4934) );
  AOI221_X1 U6599 ( .B1(n14419), .B2(n3746), .C1(n14462), .C2(n1362), .A(n4942), .ZN(n4935) );
  OAI22_X1 U6600 ( .A1(n6091), .A2(n14584), .B1(n6089), .B2(n14624), .ZN(n4942) );
  AOI221_X1 U6601 ( .B1(n14419), .B2(n3748), .C1(n14462), .C2(n1364), .A(n4950), .ZN(n4943) );
  OAI22_X1 U6602 ( .A1(n7115), .A2(n14584), .B1(n7113), .B2(n14624), .ZN(n4950) );
  AOI221_X1 U6603 ( .B1(n14418), .B2(n3749), .C1(n14461), .C2(n1365), .A(n5083), .ZN(n5076) );
  OAI22_X1 U6604 ( .A1(n9147), .A2(n14585), .B1(n9145), .B2(n14623), .ZN(n5083) );
  AOI221_X1 U6605 ( .B1(n14418), .B2(n3753), .C1(n14461), .C2(n1369), .A(n5091), .ZN(n5084) );
  OAI22_X1 U6606 ( .A1(n6075), .A2(n14585), .B1(n6073), .B2(n14623), .ZN(n5091) );
  AOI221_X1 U6607 ( .B1(n14418), .B2(n3754), .C1(n14461), .C2(n1370), .A(n5099), .ZN(n5092) );
  OAI22_X1 U6608 ( .A1(n7099), .A2(n14585), .B1(n7097), .B2(n14623), .ZN(n5099) );
  AOI221_X1 U6609 ( .B1(n14417), .B2(n3756), .C1(n14460), .C2(n1372), .A(n5232), .ZN(n5225) );
  OAI22_X1 U6610 ( .A1(n9131), .A2(n14586), .B1(n9129), .B2(n14622), .ZN(n5232) );
  AOI221_X1 U6611 ( .B1(n14416), .B2(n3757), .C1(n14459), .C2(n1373), .A(n5240), .ZN(n5233) );
  OAI22_X1 U6612 ( .A1(n6059), .A2(n14586), .B1(n6057), .B2(n14621), .ZN(n5240) );
  AOI221_X1 U6613 ( .B1(n14416), .B2(n3765), .C1(n14459), .C2(n1381), .A(n5248), .ZN(n5241) );
  OAI22_X1 U6614 ( .A1(n7083), .A2(n14586), .B1(n7081), .B2(n14621), .ZN(n5248) );
  AOI221_X1 U6615 ( .B1(n14415), .B2(n3766), .C1(n14458), .C2(n1382), .A(n5381), .ZN(n5374) );
  OAI22_X1 U6616 ( .A1(n9115), .A2(n14587), .B1(n9113), .B2(n14620), .ZN(n5381) );
  AOI221_X1 U6617 ( .B1(n14415), .B2(n3768), .C1(n14458), .C2(n1384), .A(n5389), .ZN(n5382) );
  OAI22_X1 U6618 ( .A1(n6043), .A2(n14587), .B1(n6041), .B2(n14620), .ZN(n5389) );
  AOI221_X1 U6619 ( .B1(n14415), .B2(n3769), .C1(n14458), .C2(n1385), .A(n5397), .ZN(n5390) );
  OAI22_X1 U6620 ( .A1(n7067), .A2(n14587), .B1(n7065), .B2(n14620), .ZN(n5397) );
  AOI221_X1 U6621 ( .B1(n14414), .B2(n3773), .C1(n14457), .C2(n1389), .A(n5530), .ZN(n5523) );
  OAI22_X1 U6622 ( .A1(n9099), .A2(n14588), .B1(n9097), .B2(n14619), .ZN(n5530) );
  AOI221_X1 U6623 ( .B1(n14414), .B2(n3774), .C1(n14457), .C2(n1390), .A(n5538), .ZN(n5531) );
  OAI22_X1 U6624 ( .A1(n6027), .A2(n14589), .B1(n6025), .B2(n14619), .ZN(n5538) );
  AOI221_X1 U6625 ( .B1(n14414), .B2(n3776), .C1(n14457), .C2(n1392), .A(n5546), .ZN(n5539) );
  OAI22_X1 U6626 ( .A1(n7051), .A2(n14589), .B1(n7049), .B2(n14619), .ZN(n5546) );
  AOI221_X1 U6627 ( .B1(n14413), .B2(n3777), .C1(n14456), .C2(n1393), .A(n5679), .ZN(n5672) );
  OAI22_X1 U6628 ( .A1(n9083), .A2(n14590), .B1(n9081), .B2(n14618), .ZN(n5679) );
  AOI221_X1 U6629 ( .B1(n14413), .B2(n3781), .C1(n14456), .C2(n1397), .A(n5687), .ZN(n5680) );
  OAI22_X1 U6630 ( .A1(n6011), .A2(n14590), .B1(n6009), .B2(n14618), .ZN(n5687) );
  AOI221_X1 U6631 ( .B1(n14413), .B2(n3782), .C1(n14456), .C2(n1398), .A(n5695), .ZN(n5688) );
  OAI22_X1 U6632 ( .A1(n7035), .A2(n14590), .B1(n7033), .B2(n14618), .ZN(n5695) );
  AOI221_X1 U6633 ( .B1(n14412), .B2(n3784), .C1(n14455), .C2(n1400), .A(n5820), .ZN(n5813) );
  OAI22_X1 U6634 ( .A1(n8043), .A2(n14591), .B1(n8041), .B2(n14617), .ZN(n5820) );
  AOI221_X1 U6635 ( .B1(n14412), .B2(n3785), .C1(n14455), .C2(n1401), .A(n5828), .ZN(n5821) );
  OAI22_X1 U6636 ( .A1(n9067), .A2(n14591), .B1(n9065), .B2(n14617), .ZN(n5828) );
  AOI221_X1 U6637 ( .B1(n14412), .B2(n3789), .C1(n14455), .C2(n1405), .A(n5836), .ZN(n5829) );
  OAI22_X1 U6638 ( .A1(n5995), .A2(n14591), .B1(n5993), .B2(n14616), .ZN(n5836) );
  OAI22_X1 U6639 ( .A1(n8923), .A2(n14563), .B1(n8921), .B2(n14645), .ZN(n2429) );
  OAI22_X1 U6640 ( .A1(n9947), .A2(n14563), .B1(n9945), .B2(n14645), .ZN(n2437) );
  OAI22_X1 U6641 ( .A1(n6875), .A2(n14563), .B1(n6873), .B2(n14645), .ZN(n2445) );
  OAI22_X1 U6642 ( .A1(n7899), .A2(n14563), .B1(n7897), .B2(n14645), .ZN(n2453) );
  OAI22_X1 U6643 ( .A1(n9074), .A2(n14400), .B1(n9079), .B2(n14548), .ZN(n5899) );
  OAI22_X1 U6644 ( .A1(n6002), .A2(n14400), .B1(n6007), .B2(n14548), .ZN(n5907) );
  OAI22_X1 U6645 ( .A1(n7026), .A2(n14400), .B1(n7031), .B2(n14548), .ZN(n5915) );
  OAI22_X1 U6646 ( .A1(n8562), .A2(n14400), .B1(n8567), .B2(n14548), .ZN(n5927) );
  OAI22_X1 U6647 ( .A1(n9586), .A2(n14400), .B1(n9591), .B2(n14548), .ZN(n5935) );
  OAI22_X1 U6648 ( .A1(n6514), .A2(n14400), .B1(n6519), .B2(n14548), .ZN(n5943) );
  OAI22_X1 U6649 ( .A1(n7538), .A2(n14400), .B1(n7543), .B2(n14548), .ZN(n5951) );
  OAI22_X1 U6650 ( .A1(n8538), .A2(n14361), .B1(n8543), .B2(n14509), .ZN(n1183) );
  OAI22_X1 U6651 ( .A1(n8539), .A2(n14553), .B1(n8537), .B2(n14606), .ZN(n1186) );
  OAI22_X1 U6652 ( .A1(n9050), .A2(n14361), .B1(n9055), .B2(n14509), .ZN(n1223) );
  OAI22_X1 U6653 ( .A1(n9051), .A2(n14553), .B1(n9049), .B2(n14635), .ZN(n1226) );
  OAI22_X1 U6654 ( .A1(n10074), .A2(n14361), .B1(n10079), .B2(n14509), .ZN(
        n1232) );
  OAI22_X1 U6655 ( .A1(n10075), .A2(n14553), .B1(n10073), .B2(n14635), .ZN(
        n1235) );
  OAI22_X1 U6656 ( .A1(n7002), .A2(n14361), .B1(n7007), .B2(n14509), .ZN(n1241) );
  OAI22_X1 U6657 ( .A1(n7003), .A2(n14553), .B1(n7001), .B2(n14635), .ZN(n1244) );
  OAI22_X1 U6658 ( .A1(n8026), .A2(n14361), .B1(n8031), .B2(n14509), .ZN(n1250) );
  OAI22_X1 U6659 ( .A1(n8027), .A2(n14553), .B1(n8025), .B2(n14635), .ZN(n1253) );
  OAI22_X1 U6660 ( .A1(n8546), .A2(n14361), .B1(n8551), .B2(n14509), .ZN(n1263) );
  OAI22_X1 U6661 ( .A1(n8547), .A2(n14553), .B1(n8545), .B2(n14635), .ZN(n1266) );
  OAI22_X1 U6662 ( .A1(n9570), .A2(n14361), .B1(n9575), .B2(n14509), .ZN(n1272) );
  OAI22_X1 U6663 ( .A1(n9571), .A2(n14553), .B1(n9569), .B2(n14635), .ZN(n1275) );
  OAI22_X1 U6664 ( .A1(n6498), .A2(n14361), .B1(n6503), .B2(n14509), .ZN(n1281) );
  OAI22_X1 U6665 ( .A1(n6499), .A2(n14553), .B1(n6497), .B2(n14635), .ZN(n1284) );
  OAI22_X1 U6666 ( .A1(n7522), .A2(n14362), .B1(n7527), .B2(n14510), .ZN(n1290) );
  OAI22_X1 U6667 ( .A1(n7523), .A2(n14554), .B1(n7521), .B2(n14634), .ZN(n1293) );
  OAI22_X1 U6668 ( .A1(n9058), .A2(n14362), .B1(n9063), .B2(n14510), .ZN(n1303) );
  OAI22_X1 U6669 ( .A1(n9059), .A2(n14554), .B1(n9057), .B2(n14634), .ZN(n1306) );
  OAI22_X1 U6670 ( .A1(n10082), .A2(n14362), .B1(n10087), .B2(n14510), .ZN(
        n1312) );
  OAI22_X1 U6671 ( .A1(n10083), .A2(n14554), .B1(n10081), .B2(n14634), .ZN(
        n1315) );
  OAI22_X1 U6672 ( .A1(n7010), .A2(n14362), .B1(n7015), .B2(n14510), .ZN(n1321) );
  OAI22_X1 U6673 ( .A1(n7011), .A2(n14554), .B1(n7009), .B2(n14634), .ZN(n1324) );
  OAI22_X1 U6674 ( .A1(n8034), .A2(n14362), .B1(n8039), .B2(n14510), .ZN(n1330) );
  OAI22_X1 U6675 ( .A1(n8035), .A2(n14554), .B1(n8033), .B2(n14634), .ZN(n1333) );
  OAI22_X1 U6676 ( .A1(n8522), .A2(n14362), .B1(n8527), .B2(n14510), .ZN(n1347) );
  OAI22_X1 U6677 ( .A1(n8523), .A2(n14554), .B1(n8521), .B2(n14634), .ZN(n1350) );
  OAI22_X1 U6678 ( .A1(n9034), .A2(n14362), .B1(n9039), .B2(n14510), .ZN(n1383) );
  OAI22_X1 U6679 ( .A1(n9035), .A2(n14554), .B1(n9033), .B2(n14634), .ZN(n1386) );
  OAI22_X1 U6680 ( .A1(n10058), .A2(n14362), .B1(n10063), .B2(n14510), .ZN(
        n1391) );
  OAI22_X1 U6681 ( .A1(n10059), .A2(n14554), .B1(n10057), .B2(n14634), .ZN(
        n1394) );
  OAI22_X1 U6682 ( .A1(n6986), .A2(n14362), .B1(n6991), .B2(n14510), .ZN(n1399) );
  OAI22_X1 U6683 ( .A1(n6987), .A2(n14554), .B1(n6985), .B2(n14634), .ZN(n1402) );
  OAI22_X1 U6684 ( .A1(n8010), .A2(n14362), .B1(n8015), .B2(n14510), .ZN(n1407) );
  OAI22_X1 U6685 ( .A1(n8011), .A2(n14554), .B1(n8009), .B2(n14634), .ZN(n1410) );
  OAI22_X1 U6686 ( .A1(n8530), .A2(n14363), .B1(n8535), .B2(n14511), .ZN(n1419) );
  OAI22_X1 U6687 ( .A1(n8531), .A2(n14555), .B1(n8529), .B2(n14633), .ZN(n1422) );
  OAI22_X1 U6688 ( .A1(n9554), .A2(n14363), .B1(n9559), .B2(n14511), .ZN(n1427) );
  OAI22_X1 U6689 ( .A1(n9555), .A2(n14555), .B1(n9553), .B2(n14633), .ZN(n1430) );
  OAI22_X1 U6690 ( .A1(n6482), .A2(n14363), .B1(n6487), .B2(n14511), .ZN(n1435) );
  OAI22_X1 U6691 ( .A1(n6483), .A2(n14555), .B1(n6481), .B2(n14633), .ZN(n1438) );
  OAI22_X1 U6692 ( .A1(n7506), .A2(n14363), .B1(n7511), .B2(n14511), .ZN(n1443) );
  OAI22_X1 U6693 ( .A1(n7507), .A2(n14555), .B1(n7505), .B2(n14633), .ZN(n1446) );
  OAI22_X1 U6694 ( .A1(n9042), .A2(n14363), .B1(n9047), .B2(n14511), .ZN(n1455) );
  OAI22_X1 U6695 ( .A1(n9043), .A2(n14555), .B1(n9041), .B2(n14633), .ZN(n1458) );
  OAI22_X1 U6696 ( .A1(n10066), .A2(n14363), .B1(n10071), .B2(n14511), .ZN(
        n1463) );
  OAI22_X1 U6697 ( .A1(n10067), .A2(n14555), .B1(n10065), .B2(n14633), .ZN(
        n1466) );
  OAI22_X1 U6698 ( .A1(n6994), .A2(n14363), .B1(n6999), .B2(n14511), .ZN(n1471) );
  OAI22_X1 U6699 ( .A1(n6995), .A2(n14555), .B1(n6993), .B2(n14633), .ZN(n1474) );
  OAI22_X1 U6700 ( .A1(n8018), .A2(n14363), .B1(n8023), .B2(n14511), .ZN(n1479) );
  OAI22_X1 U6701 ( .A1(n8019), .A2(n14555), .B1(n8017), .B2(n14633), .ZN(n1482) );
  OAI22_X1 U6702 ( .A1(n8506), .A2(n14363), .B1(n8511), .B2(n14511), .ZN(n1496) );
  OAI22_X1 U6703 ( .A1(n8507), .A2(n14555), .B1(n8505), .B2(n14633), .ZN(n1499) );
  OAI22_X1 U6705 ( .A1(n9018), .A2(n14363), .B1(n9023), .B2(n14511), .ZN(n1532) );
  OAI22_X1 U6706 ( .A1(n9019), .A2(n14555), .B1(n9017), .B2(n14633), .ZN(n1535) );
  OAI22_X1 U6707 ( .A1(n10042), .A2(n14364), .B1(n10047), .B2(n14512), .ZN(
        n1540) );
  OAI22_X1 U6708 ( .A1(n10043), .A2(n14556), .B1(n10041), .B2(n14632), .ZN(
        n1543) );
  OAI22_X1 U6709 ( .A1(n6970), .A2(n14364), .B1(n6975), .B2(n14512), .ZN(n1548) );
  OAI22_X1 U6710 ( .A1(n6971), .A2(n14556), .B1(n6969), .B2(n14632), .ZN(n1551) );
  OAI22_X1 U6711 ( .A1(n7994), .A2(n14364), .B1(n7999), .B2(n14512), .ZN(n1556) );
  OAI22_X1 U6712 ( .A1(n7995), .A2(n14556), .B1(n7993), .B2(n14632), .ZN(n1559) );
  OAI22_X1 U6713 ( .A1(n8514), .A2(n14364), .B1(n8519), .B2(n14512), .ZN(n1568) );
  OAI22_X1 U6714 ( .A1(n8515), .A2(n14556), .B1(n8513), .B2(n14632), .ZN(n1571) );
  OAI22_X1 U6715 ( .A1(n9538), .A2(n14364), .B1(n9543), .B2(n14512), .ZN(n1576) );
  OAI22_X1 U6716 ( .A1(n9539), .A2(n14556), .B1(n9537), .B2(n14632), .ZN(n1579) );
  OAI22_X1 U6717 ( .A1(n6466), .A2(n14364), .B1(n6471), .B2(n14512), .ZN(n1584) );
  OAI22_X1 U6718 ( .A1(n6467), .A2(n14556), .B1(n6465), .B2(n14632), .ZN(n1587) );
  OAI22_X1 U6719 ( .A1(n7490), .A2(n14364), .B1(n7495), .B2(n14512), .ZN(n1592) );
  OAI22_X1 U6720 ( .A1(n7491), .A2(n14556), .B1(n7489), .B2(n14632), .ZN(n1595) );
  OAI22_X1 U6721 ( .A1(n9026), .A2(n14364), .B1(n9031), .B2(n14512), .ZN(n1604) );
  OAI22_X1 U6722 ( .A1(n9027), .A2(n14556), .B1(n9025), .B2(n14632), .ZN(n1607) );
  OAI22_X1 U6723 ( .A1(n10050), .A2(n14364), .B1(n10055), .B2(n14512), .ZN(
        n1612) );
  OAI22_X1 U6724 ( .A1(n10051), .A2(n14556), .B1(n10049), .B2(n14632), .ZN(
        n1615) );
  OAI22_X1 U6725 ( .A1(n6978), .A2(n14364), .B1(n6983), .B2(n14512), .ZN(n1620) );
  OAI22_X1 U6726 ( .A1(n6979), .A2(n14556), .B1(n6977), .B2(n14632), .ZN(n1623) );
  OAI22_X1 U6727 ( .A1(n8002), .A2(n14364), .B1(n8007), .B2(n14512), .ZN(n1628) );
  OAI22_X1 U6728 ( .A1(n8003), .A2(n14556), .B1(n8001), .B2(n14632), .ZN(n1631) );
  OAI22_X1 U6729 ( .A1(n8490), .A2(n14364), .B1(n8495), .B2(n14512), .ZN(n1645) );
  OAI22_X1 U6730 ( .A1(n8491), .A2(n14556), .B1(n8489), .B2(n14632), .ZN(n1648) );
  OAI22_X1 U6731 ( .A1(n9002), .A2(n14365), .B1(n9007), .B2(n14513), .ZN(n1681) );
  OAI22_X1 U6732 ( .A1(n9003), .A2(n14557), .B1(n9001), .B2(n14631), .ZN(n1684) );
  OAI22_X1 U6733 ( .A1(n10026), .A2(n14365), .B1(n10031), .B2(n14513), .ZN(
        n1689) );
  OAI22_X1 U6734 ( .A1(n10027), .A2(n14557), .B1(n10025), .B2(n14631), .ZN(
        n1692) );
  OAI22_X1 U6735 ( .A1(n6954), .A2(n14365), .B1(n6959), .B2(n14513), .ZN(n1697) );
  OAI22_X1 U6736 ( .A1(n6955), .A2(n14557), .B1(n6953), .B2(n14631), .ZN(n1700) );
  OAI22_X1 U6737 ( .A1(n7978), .A2(n14365), .B1(n7983), .B2(n14513), .ZN(n1705) );
  OAI22_X1 U6738 ( .A1(n7979), .A2(n14557), .B1(n7977), .B2(n14631), .ZN(n1708) );
  OAI22_X1 U6739 ( .A1(n8498), .A2(n14365), .B1(n8503), .B2(n14513), .ZN(n1717) );
  OAI22_X1 U6740 ( .A1(n8499), .A2(n14557), .B1(n8497), .B2(n14631), .ZN(n1720) );
  OAI22_X1 U6741 ( .A1(n9522), .A2(n14365), .B1(n9527), .B2(n14513), .ZN(n1725) );
  OAI22_X1 U6742 ( .A1(n9523), .A2(n14557), .B1(n9521), .B2(n14631), .ZN(n1728) );
  OAI22_X1 U6743 ( .A1(n6450), .A2(n14365), .B1(n6455), .B2(n14513), .ZN(n1733) );
  OAI22_X1 U6744 ( .A1(n6451), .A2(n14557), .B1(n6449), .B2(n14631), .ZN(n1736) );
  OAI22_X1 U6745 ( .A1(n7474), .A2(n14365), .B1(n7479), .B2(n14513), .ZN(n1741) );
  OAI22_X1 U6746 ( .A1(n7475), .A2(n14557), .B1(n7473), .B2(n14631), .ZN(n1744) );
  OAI22_X1 U6747 ( .A1(n9010), .A2(n14365), .B1(n9015), .B2(n14513), .ZN(n1753) );
  OAI22_X1 U6748 ( .A1(n9011), .A2(n14557), .B1(n9009), .B2(n14631), .ZN(n1756) );
  OAI22_X1 U6749 ( .A1(n10034), .A2(n14365), .B1(n10039), .B2(n14513), .ZN(
        n1761) );
  OAI22_X1 U6750 ( .A1(n10035), .A2(n14557), .B1(n10033), .B2(n14631), .ZN(
        n1764) );
  OAI22_X1 U6751 ( .A1(n6962), .A2(n14365), .B1(n6967), .B2(n14513), .ZN(n1769) );
  OAI22_X1 U6752 ( .A1(n6963), .A2(n14557), .B1(n6961), .B2(n14631), .ZN(n1772) );
  OAI22_X1 U6753 ( .A1(n7986), .A2(n14366), .B1(n7991), .B2(n14514), .ZN(n1777) );
  OAI22_X1 U6754 ( .A1(n7987), .A2(n14558), .B1(n7985), .B2(n14630), .ZN(n1780) );
  OAI22_X1 U6755 ( .A1(n8474), .A2(n14366), .B1(n8479), .B2(n14514), .ZN(n1794) );
  OAI22_X1 U6756 ( .A1(n8475), .A2(n14558), .B1(n8473), .B2(n14630), .ZN(n1797) );
  OAI22_X1 U6757 ( .A1(n8986), .A2(n14366), .B1(n8991), .B2(n14514), .ZN(n1830) );
  OAI22_X1 U6758 ( .A1(n8987), .A2(n14558), .B1(n8985), .B2(n14630), .ZN(n1833) );
  OAI22_X1 U6759 ( .A1(n10010), .A2(n14366), .B1(n10015), .B2(n14514), .ZN(
        n1838) );
  OAI22_X1 U6760 ( .A1(n10011), .A2(n14558), .B1(n10009), .B2(n14630), .ZN(
        n1841) );
  OAI22_X1 U6761 ( .A1(n6938), .A2(n14366), .B1(n6943), .B2(n14514), .ZN(n1846) );
  OAI22_X1 U6762 ( .A1(n6939), .A2(n14558), .B1(n6937), .B2(n14630), .ZN(n1849) );
  OAI22_X1 U6763 ( .A1(n7962), .A2(n14366), .B1(n7967), .B2(n14514), .ZN(n1854) );
  OAI22_X1 U6764 ( .A1(n7963), .A2(n14558), .B1(n7961), .B2(n14630), .ZN(n1857) );
  OAI22_X1 U6765 ( .A1(n8482), .A2(n14366), .B1(n8487), .B2(n14514), .ZN(n1866) );
  OAI22_X1 U6766 ( .A1(n8483), .A2(n14558), .B1(n8481), .B2(n14630), .ZN(n1869) );
  OAI22_X1 U6767 ( .A1(n9506), .A2(n14366), .B1(n9511), .B2(n14514), .ZN(n1874) );
  OAI22_X1 U6768 ( .A1(n9507), .A2(n14558), .B1(n9505), .B2(n14630), .ZN(n1877) );
  OAI22_X1 U6769 ( .A1(n6434), .A2(n14366), .B1(n6439), .B2(n14514), .ZN(n1882) );
  OAI22_X1 U6770 ( .A1(n6435), .A2(n14558), .B1(n6433), .B2(n14630), .ZN(n1885) );
  OAI22_X1 U6771 ( .A1(n7458), .A2(n14366), .B1(n7463), .B2(n14514), .ZN(n1890) );
  OAI22_X1 U6772 ( .A1(n7459), .A2(n14558), .B1(n7457), .B2(n14629), .ZN(n1893) );
  OAI22_X1 U6773 ( .A1(n8994), .A2(n14367), .B1(n8999), .B2(n14515), .ZN(n1902) );
  OAI22_X1 U6774 ( .A1(n8995), .A2(n14559), .B1(n8993), .B2(n14629), .ZN(n1905) );
  OAI22_X1 U6775 ( .A1(n10018), .A2(n14367), .B1(n10023), .B2(n14515), .ZN(
        n1910) );
  OAI22_X1 U6776 ( .A1(n10019), .A2(n14559), .B1(n10017), .B2(n14629), .ZN(
        n1913) );
  OAI22_X1 U6777 ( .A1(n6946), .A2(n14367), .B1(n6951), .B2(n14515), .ZN(n1918) );
  OAI22_X1 U6778 ( .A1(n6947), .A2(n14559), .B1(n6945), .B2(n14629), .ZN(n1921) );
  OAI22_X1 U6779 ( .A1(n7970), .A2(n14367), .B1(n7975), .B2(n14515), .ZN(n1926) );
  OAI22_X1 U6780 ( .A1(n7971), .A2(n14559), .B1(n7969), .B2(n14629), .ZN(n1929) );
  OAI22_X1 U6781 ( .A1(n8458), .A2(n14367), .B1(n8463), .B2(n14515), .ZN(n1943) );
  OAI22_X1 U6782 ( .A1(n8459), .A2(n14559), .B1(n8457), .B2(n14629), .ZN(n1946) );
  OAI22_X1 U6783 ( .A1(n8970), .A2(n14367), .B1(n8975), .B2(n14515), .ZN(n1979) );
  OAI22_X1 U6784 ( .A1(n8971), .A2(n14559), .B1(n8969), .B2(n14629), .ZN(n1982) );
  OAI22_X1 U6785 ( .A1(n9994), .A2(n14367), .B1(n9999), .B2(n14515), .ZN(n1987) );
  OAI22_X1 U6786 ( .A1(n9995), .A2(n14559), .B1(n9993), .B2(n14629), .ZN(n1990) );
  OAI22_X1 U6787 ( .A1(n6922), .A2(n14367), .B1(n6927), .B2(n14515), .ZN(n1995) );
  OAI22_X1 U6788 ( .A1(n6923), .A2(n14559), .B1(n6921), .B2(n14629), .ZN(n1998) );
  OAI22_X1 U6789 ( .A1(n7946), .A2(n14367), .B1(n7951), .B2(n14515), .ZN(n2003) );
  OAI22_X1 U6790 ( .A1(n7947), .A2(n14559), .B1(n7945), .B2(n14629), .ZN(n2006) );
  OAI22_X1 U6791 ( .A1(n8466), .A2(n14367), .B1(n8471), .B2(n14515), .ZN(n2015) );
  OAI22_X1 U6792 ( .A1(n8467), .A2(n14559), .B1(n8465), .B2(n14628), .ZN(n2018) );
  OAI22_X1 U6793 ( .A1(n9490), .A2(n14368), .B1(n9495), .B2(n14516), .ZN(n2023) );
  OAI22_X1 U6794 ( .A1(n9491), .A2(n14560), .B1(n9489), .B2(n14628), .ZN(n2026) );
  OAI22_X1 U6795 ( .A1(n6418), .A2(n14368), .B1(n6423), .B2(n14516), .ZN(n2031) );
  OAI22_X1 U6796 ( .A1(n6419), .A2(n14560), .B1(n6417), .B2(n14628), .ZN(n2034) );
  OAI22_X1 U6797 ( .A1(n7442), .A2(n14368), .B1(n7447), .B2(n14516), .ZN(n2039) );
  OAI22_X1 U6798 ( .A1(n7443), .A2(n14560), .B1(n7441), .B2(n14628), .ZN(n2042) );
  OAI22_X1 U6799 ( .A1(n8978), .A2(n14368), .B1(n8983), .B2(n14516), .ZN(n2051) );
  OAI22_X1 U6800 ( .A1(n8979), .A2(n14560), .B1(n8977), .B2(n14628), .ZN(n2054) );
  OAI22_X1 U6801 ( .A1(n10002), .A2(n14368), .B1(n10007), .B2(n14516), .ZN(
        n2059) );
  OAI22_X1 U6802 ( .A1(n10003), .A2(n14560), .B1(n10001), .B2(n14628), .ZN(
        n2062) );
  OAI22_X1 U6803 ( .A1(n6930), .A2(n14368), .B1(n6935), .B2(n14516), .ZN(n2067) );
  OAI22_X1 U6804 ( .A1(n6931), .A2(n14560), .B1(n6929), .B2(n14628), .ZN(n2070) );
  OAI22_X1 U6805 ( .A1(n7954), .A2(n14368), .B1(n7959), .B2(n14516), .ZN(n2075) );
  OAI22_X1 U6806 ( .A1(n7955), .A2(n14560), .B1(n7953), .B2(n14628), .ZN(n2078) );
  OAI22_X1 U6807 ( .A1(n8442), .A2(n14368), .B1(n8447), .B2(n14516), .ZN(n2092) );
  OAI22_X1 U6808 ( .A1(n8443), .A2(n14560), .B1(n8441), .B2(n14628), .ZN(n2095) );
  OAI22_X1 U6809 ( .A1(n8954), .A2(n14368), .B1(n8959), .B2(n14516), .ZN(n2128) );
  OAI22_X1 U6810 ( .A1(n8955), .A2(n14560), .B1(n8953), .B2(n14628), .ZN(n2131) );
  OAI22_X1 U6811 ( .A1(n9978), .A2(n14368), .B1(n9983), .B2(n14516), .ZN(n2136) );
  OAI22_X1 U6812 ( .A1(n9979), .A2(n14560), .B1(n9977), .B2(n14627), .ZN(n2139) );
  OAI22_X1 U6813 ( .A1(n6906), .A2(n14369), .B1(n6911), .B2(n14517), .ZN(n2144) );
  OAI22_X1 U6814 ( .A1(n6907), .A2(n14561), .B1(n6905), .B2(n14627), .ZN(n2147) );
  OAI22_X1 U6815 ( .A1(n7930), .A2(n14369), .B1(n7935), .B2(n14517), .ZN(n2152) );
  OAI22_X1 U6816 ( .A1(n7931), .A2(n14561), .B1(n7929), .B2(n14627), .ZN(n2155) );
  OAI22_X1 U6817 ( .A1(n8450), .A2(n14369), .B1(n8455), .B2(n14517), .ZN(n2164) );
  OAI22_X1 U6818 ( .A1(n8451), .A2(n14561), .B1(n8449), .B2(n14627), .ZN(n2167) );
  OAI22_X1 U6819 ( .A1(n9474), .A2(n14369), .B1(n9479), .B2(n14517), .ZN(n2172) );
  OAI22_X1 U6820 ( .A1(n9475), .A2(n14561), .B1(n9473), .B2(n14627), .ZN(n2175) );
  OAI22_X1 U6821 ( .A1(n6402), .A2(n14369), .B1(n6407), .B2(n14517), .ZN(n2180) );
  OAI22_X1 U6822 ( .A1(n6403), .A2(n14561), .B1(n6401), .B2(n14627), .ZN(n2183) );
  OAI22_X1 U6823 ( .A1(n7426), .A2(n14369), .B1(n7431), .B2(n14517), .ZN(n2188) );
  OAI22_X1 U6824 ( .A1(n7427), .A2(n14561), .B1(n7425), .B2(n14627), .ZN(n2191) );
  OAI22_X1 U6825 ( .A1(n8962), .A2(n14369), .B1(n8967), .B2(n14517), .ZN(n2200) );
  OAI22_X1 U6826 ( .A1(n8963), .A2(n14561), .B1(n8961), .B2(n14627), .ZN(n2203) );
  OAI22_X1 U6827 ( .A1(n9986), .A2(n14369), .B1(n9991), .B2(n14517), .ZN(n2208) );
  OAI22_X1 U6828 ( .A1(n9987), .A2(n14561), .B1(n9985), .B2(n14627), .ZN(n2211) );
  OAI22_X1 U6829 ( .A1(n6914), .A2(n14369), .B1(n6919), .B2(n14517), .ZN(n2216) );
  OAI22_X1 U6830 ( .A1(n6915), .A2(n14561), .B1(n6913), .B2(n14627), .ZN(n2219) );
  OAI22_X1 U6831 ( .A1(n7938), .A2(n14369), .B1(n7943), .B2(n14517), .ZN(n2224) );
  OAI22_X1 U6832 ( .A1(n7939), .A2(n14561), .B1(n7937), .B2(n14627), .ZN(n2227) );
  OAI22_X1 U6833 ( .A1(n8426), .A2(n14369), .B1(n8431), .B2(n14517), .ZN(n2241) );
  OAI22_X1 U6834 ( .A1(n8427), .A2(n14561), .B1(n8425), .B2(n14627), .ZN(n2244) );
  OAI22_X1 U6835 ( .A1(n8938), .A2(n14370), .B1(n8943), .B2(n14518), .ZN(n2277) );
  OAI22_X1 U6836 ( .A1(n8939), .A2(n14562), .B1(n8937), .B2(n14626), .ZN(n2280) );
  OAI22_X1 U6837 ( .A1(n9962), .A2(n14370), .B1(n9967), .B2(n14518), .ZN(n2285) );
  OAI22_X1 U6838 ( .A1(n9963), .A2(n14562), .B1(n9961), .B2(n14626), .ZN(n2288) );
  OAI22_X1 U6839 ( .A1(n6890), .A2(n14370), .B1(n6895), .B2(n14518), .ZN(n2293) );
  OAI22_X1 U6840 ( .A1(n6891), .A2(n14562), .B1(n6889), .B2(n14626), .ZN(n2296) );
  OAI22_X1 U6841 ( .A1(n7914), .A2(n14370), .B1(n7919), .B2(n14518), .ZN(n2301) );
  OAI22_X1 U6842 ( .A1(n7915), .A2(n14562), .B1(n7913), .B2(n14626), .ZN(n2304) );
  OAI22_X1 U6843 ( .A1(n8434), .A2(n14370), .B1(n8439), .B2(n14518), .ZN(n2313) );
  OAI22_X1 U6844 ( .A1(n8435), .A2(n14562), .B1(n8433), .B2(n14626), .ZN(n2316) );
  OAI22_X1 U6845 ( .A1(n9458), .A2(n14370), .B1(n9463), .B2(n14518), .ZN(n2321) );
  OAI22_X1 U6846 ( .A1(n9459), .A2(n14562), .B1(n9457), .B2(n14626), .ZN(n2324) );
  OAI22_X1 U6847 ( .A1(n6386), .A2(n14370), .B1(n6391), .B2(n14518), .ZN(n2329) );
  OAI22_X1 U6848 ( .A1(n6387), .A2(n14562), .B1(n6385), .B2(n14626), .ZN(n2332) );
  OAI22_X1 U6849 ( .A1(n7410), .A2(n14370), .B1(n7415), .B2(n14518), .ZN(n2337) );
  OAI22_X1 U6850 ( .A1(n7411), .A2(n14562), .B1(n7409), .B2(n14626), .ZN(n2340) );
  OAI22_X1 U6851 ( .A1(n8946), .A2(n14370), .B1(n8951), .B2(n14518), .ZN(n2349) );
  OAI22_X1 U6852 ( .A1(n8947), .A2(n14562), .B1(n8945), .B2(n14626), .ZN(n2352) );
  OAI22_X1 U6853 ( .A1(n9970), .A2(n14370), .B1(n9975), .B2(n14518), .ZN(n2357) );
  OAI22_X1 U6854 ( .A1(n9971), .A2(n14562), .B1(n9969), .B2(n14626), .ZN(n2360) );
  OAI22_X1 U6855 ( .A1(n6898), .A2(n14370), .B1(n6903), .B2(n14518), .ZN(n2365) );
  OAI22_X1 U6857 ( .A1(n6899), .A2(n14562), .B1(n6897), .B2(n14626), .ZN(n2368) );
  OAI22_X1 U6858 ( .A1(n7922), .A2(n14370), .B1(n7927), .B2(n14518), .ZN(n2373) );
  OAI22_X1 U6859 ( .A1(n7923), .A2(n14562), .B1(n7921), .B2(n14625), .ZN(n2376) );
  OAI22_X1 U6860 ( .A1(n8410), .A2(n14371), .B1(n8415), .B2(n14519), .ZN(n2390) );
  OAI22_X1 U6861 ( .A1(n8411), .A2(n14563), .B1(n8409), .B2(n14630), .ZN(n2393) );
  OAI22_X1 U6862 ( .A1(n8922), .A2(n14371), .B1(n8927), .B2(n14519), .ZN(n2426) );
  OAI22_X1 U6863 ( .A1(n9946), .A2(n14371), .B1(n9951), .B2(n14519), .ZN(n2434) );
  OAI22_X1 U6864 ( .A1(n6874), .A2(n14371), .B1(n6879), .B2(n14519), .ZN(n2442) );
  OAI22_X1 U6865 ( .A1(n7898), .A2(n14371), .B1(n7903), .B2(n14519), .ZN(n2450) );
  OAI22_X1 U6866 ( .A1(n8418), .A2(n14371), .B1(n8423), .B2(n14519), .ZN(n2462) );
  OAI22_X1 U6867 ( .A1(n8419), .A2(n14563), .B1(n8417), .B2(n14644), .ZN(n2465) );
  OAI22_X1 U6868 ( .A1(n9442), .A2(n14371), .B1(n9447), .B2(n14519), .ZN(n2470) );
  OAI22_X1 U6869 ( .A1(n9443), .A2(n14563), .B1(n9441), .B2(n14644), .ZN(n2473) );
  OAI22_X1 U6870 ( .A1(n6370), .A2(n14371), .B1(n6375), .B2(n14519), .ZN(n2478) );
  OAI22_X1 U6871 ( .A1(n6371), .A2(n14563), .B1(n6369), .B2(n14644), .ZN(n2481) );
  OAI22_X1 U6872 ( .A1(n7394), .A2(n14371), .B1(n7399), .B2(n14519), .ZN(n2486) );
  OAI22_X1 U6873 ( .A1(n7395), .A2(n14563), .B1(n7393), .B2(n14644), .ZN(n2489) );
  OAI22_X1 U6874 ( .A1(n8930), .A2(n14371), .B1(n8935), .B2(n14519), .ZN(n2498) );
  OAI22_X1 U6875 ( .A1(n8931), .A2(n14563), .B1(n8929), .B2(n14644), .ZN(n2501) );
  OAI22_X1 U6876 ( .A1(n9954), .A2(n14372), .B1(n9959), .B2(n14520), .ZN(n2506) );
  OAI22_X1 U6877 ( .A1(n9955), .A2(n14564), .B1(n9953), .B2(n14644), .ZN(n2509) );
  OAI22_X1 U6878 ( .A1(n6882), .A2(n14372), .B1(n6887), .B2(n14520), .ZN(n2514) );
  OAI22_X1 U6879 ( .A1(n6883), .A2(n14564), .B1(n6881), .B2(n14644), .ZN(n2517) );
  OAI22_X1 U6880 ( .A1(n7906), .A2(n14372), .B1(n7911), .B2(n14520), .ZN(n2522) );
  OAI22_X1 U6881 ( .A1(n7907), .A2(n14564), .B1(n7905), .B2(n14644), .ZN(n2525) );
  OAI22_X1 U6882 ( .A1(n8394), .A2(n14372), .B1(n8399), .B2(n14520), .ZN(n2539) );
  OAI22_X1 U6883 ( .A1(n8395), .A2(n14564), .B1(n8393), .B2(n14644), .ZN(n2542) );
  OAI22_X1 U6884 ( .A1(n8906), .A2(n14372), .B1(n8911), .B2(n14520), .ZN(n2575) );
  OAI22_X1 U6885 ( .A1(n8907), .A2(n14564), .B1(n8905), .B2(n14644), .ZN(n2578) );
  OAI22_X1 U6886 ( .A1(n9930), .A2(n14372), .B1(n9935), .B2(n14520), .ZN(n2583) );
  OAI22_X1 U6887 ( .A1(n9931), .A2(n14564), .B1(n9929), .B2(n14643), .ZN(n2586) );
  OAI22_X1 U6888 ( .A1(n6858), .A2(n14372), .B1(n6863), .B2(n14520), .ZN(n2591) );
  OAI22_X1 U6889 ( .A1(n6859), .A2(n14564), .B1(n6857), .B2(n14643), .ZN(n2594) );
  OAI22_X1 U6890 ( .A1(n7882), .A2(n14372), .B1(n7887), .B2(n14520), .ZN(n2599) );
  OAI22_X1 U6891 ( .A1(n7883), .A2(n14564), .B1(n7881), .B2(n14643), .ZN(n2602) );
  OAI22_X1 U6892 ( .A1(n8402), .A2(n14372), .B1(n8407), .B2(n14520), .ZN(n2611) );
  OAI22_X1 U6893 ( .A1(n8403), .A2(n14564), .B1(n8401), .B2(n14643), .ZN(n2614) );
  OAI22_X1 U6894 ( .A1(n9426), .A2(n14372), .B1(n9431), .B2(n14520), .ZN(n2619) );
  OAI22_X1 U6895 ( .A1(n9427), .A2(n14564), .B1(n9425), .B2(n14643), .ZN(n2622) );
  OAI22_X1 U6896 ( .A1(n6354), .A2(n14373), .B1(n6359), .B2(n14521), .ZN(n2627) );
  OAI22_X1 U6897 ( .A1(n6355), .A2(n14565), .B1(n6353), .B2(n14643), .ZN(n2630) );
  OAI22_X1 U6898 ( .A1(n7378), .A2(n14373), .B1(n7383), .B2(n14521), .ZN(n2635) );
  OAI22_X1 U6899 ( .A1(n7379), .A2(n14565), .B1(n7377), .B2(n14643), .ZN(n2638) );
  OAI22_X1 U6900 ( .A1(n8914), .A2(n14373), .B1(n8919), .B2(n14521), .ZN(n2647) );
  OAI22_X1 U6901 ( .A1(n8915), .A2(n14565), .B1(n8913), .B2(n14643), .ZN(n2650) );
  OAI22_X1 U6902 ( .A1(n9938), .A2(n14373), .B1(n9943), .B2(n14521), .ZN(n2655) );
  OAI22_X1 U6903 ( .A1(n9939), .A2(n14565), .B1(n9937), .B2(n14643), .ZN(n2658) );
  OAI22_X1 U6904 ( .A1(n6866), .A2(n14373), .B1(n6871), .B2(n14521), .ZN(n2663) );
  OAI22_X1 U6905 ( .A1(n6867), .A2(n14565), .B1(n6865), .B2(n14643), .ZN(n2666) );
  OAI22_X1 U6906 ( .A1(n7890), .A2(n14373), .B1(n7895), .B2(n14521), .ZN(n2671) );
  OAI22_X1 U6907 ( .A1(n7891), .A2(n14565), .B1(n7889), .B2(n14643), .ZN(n2674) );
  OAI22_X1 U6908 ( .A1(n8378), .A2(n14373), .B1(n8383), .B2(n14521), .ZN(n2688) );
  OAI22_X1 U6909 ( .A1(n8379), .A2(n14565), .B1(n8377), .B2(n14643), .ZN(n2691) );
  OAI22_X1 U6910 ( .A1(n8890), .A2(n14373), .B1(n8895), .B2(n14521), .ZN(n2724) );
  OAI22_X1 U6911 ( .A1(n8891), .A2(n14565), .B1(n8889), .B2(n14642), .ZN(n2727) );
  OAI22_X1 U6912 ( .A1(n9914), .A2(n14373), .B1(n9919), .B2(n14521), .ZN(n2732) );
  OAI22_X1 U6913 ( .A1(n9915), .A2(n14565), .B1(n9913), .B2(n14642), .ZN(n2735) );
  OAI22_X1 U6914 ( .A1(n6842), .A2(n14373), .B1(n6847), .B2(n14521), .ZN(n2740) );
  OAI22_X1 U6915 ( .A1(n6843), .A2(n14565), .B1(n6841), .B2(n14642), .ZN(n2743) );
  OAI22_X1 U6916 ( .A1(n7866), .A2(n14374), .B1(n7871), .B2(n14522), .ZN(n2748) );
  OAI22_X1 U6917 ( .A1(n7867), .A2(n14566), .B1(n7865), .B2(n14642), .ZN(n2751) );
  OAI22_X1 U6918 ( .A1(n8386), .A2(n14374), .B1(n8391), .B2(n14522), .ZN(n2760) );
  OAI22_X1 U6919 ( .A1(n8387), .A2(n14566), .B1(n8385), .B2(n14642), .ZN(n2763) );
  OAI22_X1 U6920 ( .A1(n9410), .A2(n14374), .B1(n9415), .B2(n14522), .ZN(n2768) );
  OAI22_X1 U6921 ( .A1(n9411), .A2(n14566), .B1(n9409), .B2(n14642), .ZN(n2771) );
  OAI22_X1 U6922 ( .A1(n6338), .A2(n14374), .B1(n6343), .B2(n14522), .ZN(n2776) );
  OAI22_X1 U6923 ( .A1(n6339), .A2(n14566), .B1(n6337), .B2(n14642), .ZN(n2779) );
  OAI22_X1 U6924 ( .A1(n7362), .A2(n14374), .B1(n7367), .B2(n14522), .ZN(n2784) );
  OAI22_X1 U6925 ( .A1(n7363), .A2(n14566), .B1(n7361), .B2(n14642), .ZN(n2787) );
  OAI22_X1 U6926 ( .A1(n8898), .A2(n14374), .B1(n8903), .B2(n14522), .ZN(n2796) );
  OAI22_X1 U6927 ( .A1(n8899), .A2(n14566), .B1(n8897), .B2(n14642), .ZN(n2799) );
  OAI22_X1 U6928 ( .A1(n9922), .A2(n14374), .B1(n9927), .B2(n14522), .ZN(n2804) );
  OAI22_X1 U6929 ( .A1(n9923), .A2(n14566), .B1(n9921), .B2(n14642), .ZN(n2807) );
  OAI22_X1 U6930 ( .A1(n6850), .A2(n14374), .B1(n6855), .B2(n14522), .ZN(n2812) );
  OAI22_X1 U6931 ( .A1(n6851), .A2(n14566), .B1(n6849), .B2(n14642), .ZN(n2815) );
  OAI22_X1 U6932 ( .A1(n7874), .A2(n14374), .B1(n7879), .B2(n14522), .ZN(n2820) );
  OAI22_X1 U6933 ( .A1(n7875), .A2(n14566), .B1(n7873), .B2(n14641), .ZN(n2823) );
  OAI22_X1 U6934 ( .A1(n8362), .A2(n14374), .B1(n8367), .B2(n14522), .ZN(n2837) );
  OAI22_X1 U6935 ( .A1(n8363), .A2(n14566), .B1(n8361), .B2(n14641), .ZN(n2840) );
  OAI22_X1 U6936 ( .A1(n8874), .A2(n14375), .B1(n8879), .B2(n14523), .ZN(n2873) );
  OAI22_X1 U6937 ( .A1(n8875), .A2(n14567), .B1(n8873), .B2(n14641), .ZN(n2876) );
  OAI22_X1 U6938 ( .A1(n9898), .A2(n14375), .B1(n9903), .B2(n14523), .ZN(n2881) );
  OAI22_X1 U6939 ( .A1(n9899), .A2(n14567), .B1(n9897), .B2(n14641), .ZN(n2884) );
  OAI22_X1 U6940 ( .A1(n6826), .A2(n14375), .B1(n6831), .B2(n14523), .ZN(n2889) );
  OAI22_X1 U6941 ( .A1(n6827), .A2(n14567), .B1(n6825), .B2(n14641), .ZN(n2892) );
  OAI22_X1 U6942 ( .A1(n7850), .A2(n14375), .B1(n7855), .B2(n14523), .ZN(n2897) );
  OAI22_X1 U6943 ( .A1(n7851), .A2(n14567), .B1(n7849), .B2(n14641), .ZN(n2900) );
  OAI22_X1 U6944 ( .A1(n8370), .A2(n14375), .B1(n8375), .B2(n14523), .ZN(n2909) );
  OAI22_X1 U6945 ( .A1(n8371), .A2(n14567), .B1(n8369), .B2(n14641), .ZN(n2912) );
  OAI22_X1 U6946 ( .A1(n9394), .A2(n14375), .B1(n9399), .B2(n14523), .ZN(n2917) );
  OAI22_X1 U6947 ( .A1(n9395), .A2(n14567), .B1(n9393), .B2(n14641), .ZN(n2920) );
  OAI22_X1 U6948 ( .A1(n6322), .A2(n14375), .B1(n6327), .B2(n14523), .ZN(n2925) );
  OAI22_X1 U6949 ( .A1(n6323), .A2(n14567), .B1(n6321), .B2(n14641), .ZN(n2928) );
  OAI22_X1 U6950 ( .A1(n7346), .A2(n14375), .B1(n7351), .B2(n14523), .ZN(n2933) );
  OAI22_X1 U6951 ( .A1(n7347), .A2(n14567), .B1(n7345), .B2(n14641), .ZN(n2936) );
  OAI22_X1 U6952 ( .A1(n8882), .A2(n14375), .B1(n8887), .B2(n14523), .ZN(n2945) );
  OAI22_X1 U6953 ( .A1(n8883), .A2(n14567), .B1(n8881), .B2(n14640), .ZN(n2948) );
  OAI22_X1 U6954 ( .A1(n9906), .A2(n14375), .B1(n9911), .B2(n14523), .ZN(n2953) );
  OAI22_X1 U6955 ( .A1(n9907), .A2(n14567), .B1(n9905), .B2(n14640), .ZN(n2956) );
  OAI22_X1 U6956 ( .A1(n6834), .A2(n14375), .B1(n6839), .B2(n14523), .ZN(n2961) );
  OAI22_X1 U6957 ( .A1(n6835), .A2(n14567), .B1(n6833), .B2(n14640), .ZN(n2964) );
  OAI22_X1 U6958 ( .A1(n7858), .A2(n14375), .B1(n7863), .B2(n14523), .ZN(n2969) );
  OAI22_X1 U6959 ( .A1(n7859), .A2(n14567), .B1(n7857), .B2(n14640), .ZN(n2972) );
  OAI22_X1 U6960 ( .A1(n8346), .A2(n14375), .B1(n8351), .B2(n14523), .ZN(n2986) );
  OAI22_X1 U6961 ( .A1(n8347), .A2(n14567), .B1(n8345), .B2(n14640), .ZN(n2989) );
  OAI22_X1 U6962 ( .A1(n8858), .A2(n14376), .B1(n8863), .B2(n14524), .ZN(n3022) );
  OAI22_X1 U6963 ( .A1(n8859), .A2(n14568), .B1(n8857), .B2(n14640), .ZN(n3025) );
  OAI22_X1 U6964 ( .A1(n9882), .A2(n14376), .B1(n9887), .B2(n14524), .ZN(n3030) );
  OAI22_X1 U6965 ( .A1(n9883), .A2(n14568), .B1(n9881), .B2(n14640), .ZN(n3033) );
  OAI22_X1 U6966 ( .A1(n6810), .A2(n14376), .B1(n6815), .B2(n14524), .ZN(n3038) );
  OAI22_X1 U6967 ( .A1(n6811), .A2(n14568), .B1(n6809), .B2(n14640), .ZN(n3041) );
  OAI22_X1 U6968 ( .A1(n7834), .A2(n14376), .B1(n7839), .B2(n14524), .ZN(n3046) );
  OAI22_X1 U6969 ( .A1(n7835), .A2(n14568), .B1(n7833), .B2(n14640), .ZN(n3049) );
  OAI22_X1 U6970 ( .A1(n8354), .A2(n14376), .B1(n8359), .B2(n14524), .ZN(n3058) );
  OAI22_X1 U6971 ( .A1(n8355), .A2(n14568), .B1(n8353), .B2(n14639), .ZN(n3061) );
  OAI22_X1 U6972 ( .A1(n9378), .A2(n14376), .B1(n9383), .B2(n14524), .ZN(n3066) );
  OAI22_X1 U6973 ( .A1(n9379), .A2(n14568), .B1(n9377), .B2(n14639), .ZN(n3069) );
  OAI22_X1 U6974 ( .A1(n6306), .A2(n14376), .B1(n6311), .B2(n14524), .ZN(n3074) );
  OAI22_X1 U6975 ( .A1(n6307), .A2(n14568), .B1(n6305), .B2(n14639), .ZN(n3077) );
  OAI22_X1 U6976 ( .A1(n7330), .A2(n14376), .B1(n7335), .B2(n14524), .ZN(n3082) );
  OAI22_X1 U6977 ( .A1(n7331), .A2(n14568), .B1(n7329), .B2(n14639), .ZN(n3085) );
  OAI22_X1 U6978 ( .A1(n8866), .A2(n14376), .B1(n8871), .B2(n14524), .ZN(n3094) );
  OAI22_X1 U6979 ( .A1(n8867), .A2(n14568), .B1(n8865), .B2(n14639), .ZN(n3097) );
  OAI22_X1 U6980 ( .A1(n9890), .A2(n14376), .B1(n9895), .B2(n14524), .ZN(n3102) );
  OAI22_X1 U6981 ( .A1(n9891), .A2(n14568), .B1(n9889), .B2(n14639), .ZN(n3105) );
  OAI22_X1 U6982 ( .A1(n6818), .A2(n14377), .B1(n6823), .B2(n14525), .ZN(n3110) );
  OAI22_X1 U6983 ( .A1(n6819), .A2(n14569), .B1(n6817), .B2(n14639), .ZN(n3113) );
  OAI22_X1 U6984 ( .A1(n7842), .A2(n14377), .B1(n7847), .B2(n14525), .ZN(n3118) );
  OAI22_X1 U6985 ( .A1(n7843), .A2(n14569), .B1(n7841), .B2(n14639), .ZN(n3121) );
  OAI22_X1 U6986 ( .A1(n8330), .A2(n14377), .B1(n8335), .B2(n14525), .ZN(n3135) );
  OAI22_X1 U6987 ( .A1(n8331), .A2(n14569), .B1(n8329), .B2(n14639), .ZN(n3138) );
  OAI22_X1 U6988 ( .A1(n8842), .A2(n14377), .B1(n8847), .B2(n14525), .ZN(n3171) );
  OAI22_X1 U6989 ( .A1(n8843), .A2(n14569), .B1(n8841), .B2(n14639), .ZN(n3174) );
  OAI22_X1 U6990 ( .A1(n9866), .A2(n14377), .B1(n9871), .B2(n14525), .ZN(n3179) );
  OAI22_X1 U6991 ( .A1(n9867), .A2(n14569), .B1(n9865), .B2(n14638), .ZN(n3182) );
  OAI22_X1 U6992 ( .A1(n6794), .A2(n14377), .B1(n6799), .B2(n14525), .ZN(n3187) );
  OAI22_X1 U6993 ( .A1(n6795), .A2(n14569), .B1(n6793), .B2(n14638), .ZN(n3190) );
  OAI22_X1 U6994 ( .A1(n7818), .A2(n14377), .B1(n7823), .B2(n14525), .ZN(n3195) );
  OAI22_X1 U6995 ( .A1(n7819), .A2(n14569), .B1(n7817), .B2(n14638), .ZN(n3198) );
  OAI22_X1 U6996 ( .A1(n8338), .A2(n14377), .B1(n8343), .B2(n14525), .ZN(n3207) );
  OAI22_X1 U6997 ( .A1(n8339), .A2(n14569), .B1(n8337), .B2(n14638), .ZN(n3210) );
  OAI22_X1 U6998 ( .A1(n9362), .A2(n14377), .B1(n9367), .B2(n14525), .ZN(n3215) );
  OAI22_X1 U6999 ( .A1(n9363), .A2(n14569), .B1(n9361), .B2(n14638), .ZN(n3218) );
  OAI22_X1 U7000 ( .A1(n6290), .A2(n14377), .B1(n6295), .B2(n14525), .ZN(n3223) );
  OAI22_X1 U7001 ( .A1(n6291), .A2(n14569), .B1(n6289), .B2(n14638), .ZN(n3226) );
  OAI22_X1 U7002 ( .A1(n7314), .A2(n14378), .B1(n7319), .B2(n14526), .ZN(n3231) );
  OAI22_X1 U7003 ( .A1(n7315), .A2(n14570), .B1(n7313), .B2(n14638), .ZN(n3234) );
  OAI22_X1 U7004 ( .A1(n8850), .A2(n14378), .B1(n8855), .B2(n14526), .ZN(n3243) );
  OAI22_X1 U7005 ( .A1(n8851), .A2(n14570), .B1(n8849), .B2(n14638), .ZN(n3246) );
  OAI22_X1 U7006 ( .A1(n9874), .A2(n14378), .B1(n9879), .B2(n14526), .ZN(n3251) );
  OAI22_X1 U7007 ( .A1(n9875), .A2(n14570), .B1(n9873), .B2(n14638), .ZN(n3254) );
  OAI22_X1 U7009 ( .A1(n6802), .A2(n14378), .B1(n6807), .B2(n14526), .ZN(n3259) );
  OAI22_X1 U7010 ( .A1(n6803), .A2(n14570), .B1(n6801), .B2(n14638), .ZN(n3262) );
  OAI22_X1 U7011 ( .A1(n7826), .A2(n14378), .B1(n7831), .B2(n14526), .ZN(n3267) );
  OAI22_X1 U7012 ( .A1(n7827), .A2(n14570), .B1(n7825), .B2(n14638), .ZN(n3270) );
  OAI22_X1 U7013 ( .A1(n8314), .A2(n14378), .B1(n8319), .B2(n14526), .ZN(n3284) );
  OAI22_X1 U7014 ( .A1(n8315), .A2(n14570), .B1(n8313), .B2(n14638), .ZN(n3287) );
  OAI22_X1 U7015 ( .A1(n8826), .A2(n14378), .B1(n8831), .B2(n14526), .ZN(n3320) );
  OAI22_X1 U7016 ( .A1(n8827), .A2(n14570), .B1(n8825), .B2(n14637), .ZN(n3323) );
  OAI22_X1 U7017 ( .A1(n9850), .A2(n14378), .B1(n9855), .B2(n14526), .ZN(n3328) );
  OAI22_X1 U7018 ( .A1(n9851), .A2(n14570), .B1(n9849), .B2(n14637), .ZN(n3331) );
  OAI22_X1 U7019 ( .A1(n6778), .A2(n14378), .B1(n6783), .B2(n14526), .ZN(n3336) );
  OAI22_X1 U7020 ( .A1(n6779), .A2(n14570), .B1(n6777), .B2(n14637), .ZN(n3339) );
  OAI22_X1 U7021 ( .A1(n7802), .A2(n14378), .B1(n7807), .B2(n14526), .ZN(n3344) );
  OAI22_X1 U7022 ( .A1(n7803), .A2(n14570), .B1(n7801), .B2(n14637), .ZN(n3347) );
  OAI22_X1 U7023 ( .A1(n8322), .A2(n14379), .B1(n8327), .B2(n14527), .ZN(n3356) );
  OAI22_X1 U7024 ( .A1(n8323), .A2(n14571), .B1(n8321), .B2(n14637), .ZN(n3359) );
  OAI22_X1 U7025 ( .A1(n9346), .A2(n14379), .B1(n9351), .B2(n14527), .ZN(n3364) );
  OAI22_X1 U7026 ( .A1(n9347), .A2(n14571), .B1(n9345), .B2(n14637), .ZN(n3367) );
  OAI22_X1 U7027 ( .A1(n6274), .A2(n14379), .B1(n6279), .B2(n14527), .ZN(n3372) );
  OAI22_X1 U7028 ( .A1(n6275), .A2(n14571), .B1(n6273), .B2(n14637), .ZN(n3375) );
  OAI22_X1 U7029 ( .A1(n7298), .A2(n14379), .B1(n7303), .B2(n14527), .ZN(n3380) );
  OAI22_X1 U7030 ( .A1(n7299), .A2(n14571), .B1(n7297), .B2(n14637), .ZN(n3383) );
  OAI22_X1 U7031 ( .A1(n8834), .A2(n14379), .B1(n8839), .B2(n14527), .ZN(n3392) );
  OAI22_X1 U7032 ( .A1(n8835), .A2(n14571), .B1(n8833), .B2(n14637), .ZN(n3395) );
  OAI22_X1 U7033 ( .A1(n9858), .A2(n14379), .B1(n9863), .B2(n14527), .ZN(n3400) );
  OAI22_X1 U7034 ( .A1(n9859), .A2(n14571), .B1(n9857), .B2(n14637), .ZN(n3403) );
  OAI22_X1 U7035 ( .A1(n6786), .A2(n14379), .B1(n6791), .B2(n14527), .ZN(n3408) );
  OAI22_X1 U7036 ( .A1(n6787), .A2(n14571), .B1(n6785), .B2(n14637), .ZN(n3411) );
  OAI22_X1 U7037 ( .A1(n7810), .A2(n14379), .B1(n7815), .B2(n14527), .ZN(n3416) );
  OAI22_X1 U7038 ( .A1(n7811), .A2(n14571), .B1(n7809), .B2(n14636), .ZN(n3419) );
  OAI22_X1 U7039 ( .A1(n8298), .A2(n14379), .B1(n8303), .B2(n14527), .ZN(n3433) );
  OAI22_X1 U7040 ( .A1(n8299), .A2(n14571), .B1(n8297), .B2(n14636), .ZN(n3436) );
  OAI22_X1 U7041 ( .A1(n8810), .A2(n14379), .B1(n8815), .B2(n14527), .ZN(n3469) );
  OAI22_X1 U7042 ( .A1(n8811), .A2(n14571), .B1(n8809), .B2(n14636), .ZN(n3472) );
  OAI22_X1 U7043 ( .A1(n9834), .A2(n14380), .B1(n9839), .B2(n14528), .ZN(n3477) );
  OAI22_X1 U7044 ( .A1(n9835), .A2(n14572), .B1(n9833), .B2(n14636), .ZN(n3480) );
  OAI22_X1 U7045 ( .A1(n6762), .A2(n14380), .B1(n6767), .B2(n14528), .ZN(n3485) );
  OAI22_X1 U7046 ( .A1(n6763), .A2(n14572), .B1(n6761), .B2(n14636), .ZN(n3488) );
  OAI22_X1 U7047 ( .A1(n7786), .A2(n14380), .B1(n7791), .B2(n14528), .ZN(n3493) );
  OAI22_X1 U7048 ( .A1(n7787), .A2(n14572), .B1(n7785), .B2(n14636), .ZN(n3496) );
  OAI22_X1 U7049 ( .A1(n8306), .A2(n14380), .B1(n8311), .B2(n14528), .ZN(n3505) );
  OAI22_X1 U7050 ( .A1(n8307), .A2(n14572), .B1(n8305), .B2(n14636), .ZN(n3508) );
  OAI22_X1 U7051 ( .A1(n9330), .A2(n14380), .B1(n9335), .B2(n14528), .ZN(n3513) );
  OAI22_X1 U7052 ( .A1(n9331), .A2(n14572), .B1(n9329), .B2(n14636), .ZN(n3516) );
  OAI22_X1 U7053 ( .A1(n6258), .A2(n14380), .B1(n6263), .B2(n14528), .ZN(n3521) );
  OAI22_X1 U7054 ( .A1(n6259), .A2(n14572), .B1(n6257), .B2(n14636), .ZN(n3524) );
  OAI22_X1 U7055 ( .A1(n7282), .A2(n14380), .B1(n7287), .B2(n14528), .ZN(n3529) );
  OAI22_X1 U7056 ( .A1(n7283), .A2(n14572), .B1(n7281), .B2(n14636), .ZN(n3532) );
  OAI22_X1 U7057 ( .A1(n8818), .A2(n14380), .B1(n8823), .B2(n14528), .ZN(n3541) );
  OAI22_X1 U7058 ( .A1(n8819), .A2(n14572), .B1(n8817), .B2(n14635), .ZN(n3544) );
  OAI22_X1 U7059 ( .A1(n9842), .A2(n14380), .B1(n9847), .B2(n14528), .ZN(n3549) );
  OAI22_X1 U7060 ( .A1(n9843), .A2(n14572), .B1(n9841), .B2(n14635), .ZN(n3552) );
  OAI22_X1 U7061 ( .A1(n6770), .A2(n14380), .B1(n6775), .B2(n14528), .ZN(n3557) );
  OAI22_X1 U7062 ( .A1(n6771), .A2(n14572), .B1(n6769), .B2(n14635), .ZN(n3560) );
  OAI22_X1 U7063 ( .A1(n7794), .A2(n14380), .B1(n7799), .B2(n14528), .ZN(n3565) );
  OAI22_X1 U7064 ( .A1(n7795), .A2(n14572), .B1(n7793), .B2(n14640), .ZN(n3568) );
  OAI22_X1 U7065 ( .A1(n8282), .A2(n14380), .B1(n8287), .B2(n14528), .ZN(n3582) );
  OAI22_X1 U7066 ( .A1(n8283), .A2(n14572), .B1(n8281), .B2(n14616), .ZN(n3585) );
  OAI22_X1 U7067 ( .A1(n8794), .A2(n14381), .B1(n8799), .B2(n14529), .ZN(n3618) );
  OAI22_X1 U7068 ( .A1(n8795), .A2(n14573), .B1(n8793), .B2(n14615), .ZN(n3621) );
  OAI22_X1 U7069 ( .A1(n9818), .A2(n14381), .B1(n9823), .B2(n14529), .ZN(n3626) );
  OAI22_X1 U7070 ( .A1(n9819), .A2(n14573), .B1(n9817), .B2(n14615), .ZN(n3629) );
  OAI22_X1 U7071 ( .A1(n6746), .A2(n14381), .B1(n6751), .B2(n14529), .ZN(n3634) );
  OAI22_X1 U7072 ( .A1(n6747), .A2(n14573), .B1(n6745), .B2(n14615), .ZN(n3637) );
  OAI22_X1 U7073 ( .A1(n7770), .A2(n14381), .B1(n7775), .B2(n14529), .ZN(n3642) );
  OAI22_X1 U7074 ( .A1(n7771), .A2(n14573), .B1(n7769), .B2(n14615), .ZN(n3645) );
  OAI22_X1 U7075 ( .A1(n8290), .A2(n14381), .B1(n8295), .B2(n14529), .ZN(n3654) );
  OAI22_X1 U7076 ( .A1(n8291), .A2(n14573), .B1(n8289), .B2(n14615), .ZN(n3657) );
  OAI22_X1 U7077 ( .A1(n9314), .A2(n14381), .B1(n9319), .B2(n14529), .ZN(n3662) );
  OAI22_X1 U7078 ( .A1(n9315), .A2(n14573), .B1(n9313), .B2(n14615), .ZN(n3665) );
  OAI22_X1 U7079 ( .A1(n7266), .A2(n14381), .B1(n7271), .B2(n14529), .ZN(n3678) );
  OAI22_X1 U7080 ( .A1(n7267), .A2(n14573), .B1(n7265), .B2(n14615), .ZN(n3681) );
  OAI22_X1 U7081 ( .A1(n6242), .A2(n14381), .B1(n6247), .B2(n14529), .ZN(n3670) );
  OAI22_X1 U7082 ( .A1(n6243), .A2(n14573), .B1(n6241), .B2(n14615), .ZN(n3673) );
  OAI22_X1 U7083 ( .A1(n8802), .A2(n14381), .B1(n8807), .B2(n14529), .ZN(n3690) );
  OAI22_X1 U7084 ( .A1(n8803), .A2(n14573), .B1(n8801), .B2(n14615), .ZN(n3693) );
  OAI22_X1 U7085 ( .A1(n9826), .A2(n14381), .B1(n9831), .B2(n14529), .ZN(n3698) );
  OAI22_X1 U7086 ( .A1(n9827), .A2(n14573), .B1(n9825), .B2(n14615), .ZN(n3701) );
  OAI22_X1 U7087 ( .A1(n6754), .A2(n14381), .B1(n6759), .B2(n14529), .ZN(n3706) );
  OAI22_X1 U7088 ( .A1(n6755), .A2(n14573), .B1(n6753), .B2(n14614), .ZN(n3709) );
  OAI22_X1 U7089 ( .A1(n7778), .A2(n14382), .B1(n7783), .B2(n14530), .ZN(n3714) );
  OAI22_X1 U7090 ( .A1(n7779), .A2(n14574), .B1(n7777), .B2(n14614), .ZN(n3717) );
  OAI22_X1 U7091 ( .A1(n8266), .A2(n14382), .B1(n8271), .B2(n14530), .ZN(n3731) );
  OAI22_X1 U7092 ( .A1(n8267), .A2(n14574), .B1(n8265), .B2(n14614), .ZN(n3734) );
  OAI22_X1 U7093 ( .A1(n8778), .A2(n14382), .B1(n8783), .B2(n14530), .ZN(n3767) );
  OAI22_X1 U7094 ( .A1(n8779), .A2(n14574), .B1(n8777), .B2(n14614), .ZN(n3770) );
  OAI22_X1 U7095 ( .A1(n9802), .A2(n14382), .B1(n9807), .B2(n14530), .ZN(n3775) );
  OAI22_X1 U7096 ( .A1(n9803), .A2(n14574), .B1(n9801), .B2(n14614), .ZN(n3778) );
  OAI22_X1 U7097 ( .A1(n6730), .A2(n14382), .B1(n6735), .B2(n14530), .ZN(n3783) );
  OAI22_X1 U7098 ( .A1(n6731), .A2(n14574), .B1(n6729), .B2(n14614), .ZN(n3786) );
  OAI22_X1 U7099 ( .A1(n7754), .A2(n14382), .B1(n7759), .B2(n14530), .ZN(n3791) );
  OAI22_X1 U7100 ( .A1(n7755), .A2(n14574), .B1(n7753), .B2(n14614), .ZN(n3794) );
  OAI22_X1 U7101 ( .A1(n8274), .A2(n14382), .B1(n8279), .B2(n14530), .ZN(n3803) );
  OAI22_X1 U7102 ( .A1(n8275), .A2(n14574), .B1(n8273), .B2(n14614), .ZN(n3806) );
  OAI22_X1 U7103 ( .A1(n9298), .A2(n14382), .B1(n9303), .B2(n14530), .ZN(n3811) );
  OAI22_X1 U7104 ( .A1(n9299), .A2(n14574), .B1(n9297), .B2(n14614), .ZN(n3814) );
  OAI22_X1 U7105 ( .A1(n6226), .A2(n14382), .B1(n6231), .B2(n14530), .ZN(n3819) );
  OAI22_X1 U7106 ( .A1(n6227), .A2(n14574), .B1(n6225), .B2(n14614), .ZN(n3822) );
  OAI22_X1 U7107 ( .A1(n7250), .A2(n14382), .B1(n7255), .B2(n14530), .ZN(n3827) );
  OAI22_X1 U7108 ( .A1(n7251), .A2(n14574), .B1(n7249), .B2(n14613), .ZN(n3830) );
  OAI22_X1 U7109 ( .A1(n8786), .A2(n14383), .B1(n8791), .B2(n14531), .ZN(n3839) );
  OAI22_X1 U7110 ( .A1(n8787), .A2(n14575), .B1(n8785), .B2(n14613), .ZN(n3842) );
  OAI22_X1 U7111 ( .A1(n9810), .A2(n14383), .B1(n9815), .B2(n14531), .ZN(n3847) );
  OAI22_X1 U7112 ( .A1(n9811), .A2(n14575), .B1(n9809), .B2(n14613), .ZN(n3850) );
  OAI22_X1 U7113 ( .A1(n6738), .A2(n14383), .B1(n6743), .B2(n14531), .ZN(n3855) );
  OAI22_X1 U7114 ( .A1(n6739), .A2(n14575), .B1(n6737), .B2(n14613), .ZN(n3858) );
  OAI22_X1 U7115 ( .A1(n7762), .A2(n14383), .B1(n7767), .B2(n14531), .ZN(n3863) );
  OAI22_X1 U7116 ( .A1(n7763), .A2(n14575), .B1(n7761), .B2(n14613), .ZN(n3866) );
  OAI22_X1 U7117 ( .A1(n8250), .A2(n14383), .B1(n8255), .B2(n14531), .ZN(n3880) );
  OAI22_X1 U7118 ( .A1(n8251), .A2(n14575), .B1(n8249), .B2(n14613), .ZN(n3883) );
  OAI22_X1 U7119 ( .A1(n8762), .A2(n14383), .B1(n8767), .B2(n14531), .ZN(n3916) );
  OAI22_X1 U7120 ( .A1(n8763), .A2(n14575), .B1(n8761), .B2(n14613), .ZN(n3919) );
  OAI22_X1 U7121 ( .A1(n9786), .A2(n14383), .B1(n9791), .B2(n14531), .ZN(n3924) );
  OAI22_X1 U7122 ( .A1(n9787), .A2(n14575), .B1(n9785), .B2(n14613), .ZN(n3927) );
  OAI22_X1 U7123 ( .A1(n6714), .A2(n14383), .B1(n6719), .B2(n14531), .ZN(n3932) );
  OAI22_X1 U7124 ( .A1(n6715), .A2(n14575), .B1(n6713), .B2(n14613), .ZN(n3935) );
  OAI22_X1 U7125 ( .A1(n7738), .A2(n14383), .B1(n7743), .B2(n14531), .ZN(n3940) );
  OAI22_X1 U7126 ( .A1(n7739), .A2(n14575), .B1(n7737), .B2(n14613), .ZN(n3943) );
  OAI22_X1 U7127 ( .A1(n8258), .A2(n14383), .B1(n8263), .B2(n14531), .ZN(n3952) );
  OAI22_X1 U7128 ( .A1(n8259), .A2(n14575), .B1(n8257), .B2(n14612), .ZN(n3955) );
  OAI22_X1 U7129 ( .A1(n9282), .A2(n14384), .B1(n9287), .B2(n14532), .ZN(n3960) );
  OAI22_X1 U7130 ( .A1(n9283), .A2(n14576), .B1(n9281), .B2(n14612), .ZN(n3963) );
  OAI22_X1 U7131 ( .A1(n6210), .A2(n14384), .B1(n6215), .B2(n14532), .ZN(n3968) );
  OAI22_X1 U7132 ( .A1(n6211), .A2(n14576), .B1(n6209), .B2(n14612), .ZN(n3971) );
  OAI22_X1 U7133 ( .A1(n7234), .A2(n14384), .B1(n7239), .B2(n14532), .ZN(n3976) );
  OAI22_X1 U7134 ( .A1(n7235), .A2(n14576), .B1(n7233), .B2(n14612), .ZN(n3979) );
  OAI22_X1 U7135 ( .A1(n8770), .A2(n14384), .B1(n8775), .B2(n14532), .ZN(n3988) );
  OAI22_X1 U7136 ( .A1(n8771), .A2(n14576), .B1(n8769), .B2(n14612), .ZN(n3991) );
  OAI22_X1 U7137 ( .A1(n9794), .A2(n14384), .B1(n9799), .B2(n14532), .ZN(n3996) );
  OAI22_X1 U7138 ( .A1(n9795), .A2(n14576), .B1(n9793), .B2(n14612), .ZN(n3999) );
  OAI22_X1 U7139 ( .A1(n6722), .A2(n14384), .B1(n6727), .B2(n14532), .ZN(n4004) );
  OAI22_X1 U7140 ( .A1(n6723), .A2(n14576), .B1(n6721), .B2(n14612), .ZN(n4007) );
  OAI22_X1 U7141 ( .A1(n7746), .A2(n14384), .B1(n7751), .B2(n14532), .ZN(n4012) );
  OAI22_X1 U7142 ( .A1(n7747), .A2(n14576), .B1(n7745), .B2(n14612), .ZN(n4015) );
  OAI22_X1 U7143 ( .A1(n8234), .A2(n14384), .B1(n8239), .B2(n14532), .ZN(n4029) );
  OAI22_X1 U7144 ( .A1(n8235), .A2(n14576), .B1(n8233), .B2(n14612), .ZN(n4032) );
  OAI22_X1 U7145 ( .A1(n8746), .A2(n14384), .B1(n8751), .B2(n14532), .ZN(n4065) );
  OAI22_X1 U7146 ( .A1(n8747), .A2(n14576), .B1(n8745), .B2(n14612), .ZN(n4068) );
  OAI22_X1 U7147 ( .A1(n9770), .A2(n14384), .B1(n9775), .B2(n14532), .ZN(n4073) );
  OAI22_X1 U7148 ( .A1(n9771), .A2(n14576), .B1(n9769), .B2(n14611), .ZN(n4076) );
  OAI22_X1 U7149 ( .A1(n6698), .A2(n14385), .B1(n6703), .B2(n14533), .ZN(n4081) );
  OAI22_X1 U7150 ( .A1(n6699), .A2(n14577), .B1(n6697), .B2(n14611), .ZN(n4084) );
  OAI22_X1 U7151 ( .A1(n7722), .A2(n14385), .B1(n7727), .B2(n14533), .ZN(n4089) );
  OAI22_X1 U7152 ( .A1(n7723), .A2(n14577), .B1(n7721), .B2(n14611), .ZN(n4092) );
  OAI22_X1 U7153 ( .A1(n8242), .A2(n14385), .B1(n8247), .B2(n14533), .ZN(n4101) );
  OAI22_X1 U7154 ( .A1(n8243), .A2(n14577), .B1(n8241), .B2(n14611), .ZN(n4104) );
  OAI22_X1 U7155 ( .A1(n9266), .A2(n14385), .B1(n9271), .B2(n14533), .ZN(n4109) );
  OAI22_X1 U7156 ( .A1(n9267), .A2(n14577), .B1(n9265), .B2(n14611), .ZN(n4112) );
  OAI22_X1 U7157 ( .A1(n6194), .A2(n14385), .B1(n6199), .B2(n14533), .ZN(n4117) );
  OAI22_X1 U7158 ( .A1(n6195), .A2(n14577), .B1(n6193), .B2(n14611), .ZN(n4120) );
  OAI22_X1 U7159 ( .A1(n7218), .A2(n14385), .B1(n7223), .B2(n14533), .ZN(n4125) );
  OAI22_X1 U7161 ( .A1(n7219), .A2(n14577), .B1(n7217), .B2(n14611), .ZN(n4128) );
  OAI22_X1 U7162 ( .A1(n8754), .A2(n14385), .B1(n8759), .B2(n14533), .ZN(n4137) );
  OAI22_X1 U7163 ( .A1(n8755), .A2(n14577), .B1(n8753), .B2(n14611), .ZN(n4140) );
  OAI22_X1 U7164 ( .A1(n9778), .A2(n14385), .B1(n9783), .B2(n14533), .ZN(n4145) );
  OAI22_X1 U7165 ( .A1(n9779), .A2(n14577), .B1(n9777), .B2(n14611), .ZN(n4148) );
  OAI22_X1 U7166 ( .A1(n6706), .A2(n14385), .B1(n6711), .B2(n14533), .ZN(n4153) );
  OAI22_X1 U7167 ( .A1(n6707), .A2(n14577), .B1(n6705), .B2(n14611), .ZN(n4156) );
  OAI22_X1 U7168 ( .A1(n7730), .A2(n14385), .B1(n7735), .B2(n14533), .ZN(n4161) );
  OAI22_X1 U7169 ( .A1(n7731), .A2(n14577), .B1(n7729), .B2(n14611), .ZN(n4164) );
  OAI22_X1 U7170 ( .A1(n8218), .A2(n14385), .B1(n8223), .B2(n14533), .ZN(n4178) );
  OAI22_X1 U7171 ( .A1(n8219), .A2(n14577), .B1(n8217), .B2(n14611), .ZN(n4181) );
  OAI22_X1 U7172 ( .A1(n8730), .A2(n14386), .B1(n8735), .B2(n14534), .ZN(n4214) );
  OAI22_X1 U7173 ( .A1(n8731), .A2(n14578), .B1(n8729), .B2(n14610), .ZN(n4217) );
  OAI22_X1 U7174 ( .A1(n9754), .A2(n14386), .B1(n9759), .B2(n14534), .ZN(n4222) );
  OAI22_X1 U7175 ( .A1(n9755), .A2(n14578), .B1(n9753), .B2(n14610), .ZN(n4225) );
  OAI22_X1 U7176 ( .A1(n6682), .A2(n14386), .B1(n6687), .B2(n14534), .ZN(n4230) );
  OAI22_X1 U7177 ( .A1(n6683), .A2(n14578), .B1(n6681), .B2(n14610), .ZN(n4233) );
  OAI22_X1 U7178 ( .A1(n7706), .A2(n14386), .B1(n7711), .B2(n14534), .ZN(n4238) );
  OAI22_X1 U7179 ( .A1(n7707), .A2(n14578), .B1(n7705), .B2(n14610), .ZN(n4241) );
  OAI22_X1 U7180 ( .A1(n8226), .A2(n14386), .B1(n8231), .B2(n14534), .ZN(n4250) );
  OAI22_X1 U7181 ( .A1(n8227), .A2(n14578), .B1(n8225), .B2(n14610), .ZN(n4253) );
  OAI22_X1 U7182 ( .A1(n9250), .A2(n14386), .B1(n9255), .B2(n14534), .ZN(n4258) );
  OAI22_X1 U7183 ( .A1(n9251), .A2(n14578), .B1(n9249), .B2(n14610), .ZN(n4261) );
  OAI22_X1 U7184 ( .A1(n6178), .A2(n14386), .B1(n6183), .B2(n14534), .ZN(n4266) );
  OAI22_X1 U7185 ( .A1(n6179), .A2(n14578), .B1(n6177), .B2(n14610), .ZN(n4269) );
  OAI22_X1 U7186 ( .A1(n7202), .A2(n14386), .B1(n7207), .B2(n14534), .ZN(n4274) );
  OAI22_X1 U7187 ( .A1(n7203), .A2(n14578), .B1(n7201), .B2(n14610), .ZN(n4277) );
  OAI22_X1 U7188 ( .A1(n8738), .A2(n14386), .B1(n8743), .B2(n14534), .ZN(n4286) );
  OAI22_X1 U7189 ( .A1(n8739), .A2(n14578), .B1(n8737), .B2(n14610), .ZN(n4289) );
  OAI22_X1 U7190 ( .A1(n9762), .A2(n14386), .B1(n9767), .B2(n14534), .ZN(n4294) );
  OAI22_X1 U7191 ( .A1(n9763), .A2(n14578), .B1(n9761), .B2(n14610), .ZN(n4297) );
  OAI22_X1 U7192 ( .A1(n6690), .A2(n14386), .B1(n6695), .B2(n14534), .ZN(n4302) );
  OAI22_X1 U7193 ( .A1(n6691), .A2(n14578), .B1(n6689), .B2(n14609), .ZN(n4305) );
  OAI22_X1 U7194 ( .A1(n7714), .A2(n14386), .B1(n7719), .B2(n14534), .ZN(n4310) );
  OAI22_X1 U7195 ( .A1(n7715), .A2(n14578), .B1(n7713), .B2(n14609), .ZN(n4313) );
  OAI22_X1 U7196 ( .A1(n8202), .A2(n14387), .B1(n8207), .B2(n14535), .ZN(n4327) );
  OAI22_X1 U7197 ( .A1(n8203), .A2(n14579), .B1(n8201), .B2(n14609), .ZN(n4330) );
  OAI22_X1 U7198 ( .A1(n8714), .A2(n14387), .B1(n8719), .B2(n14535), .ZN(n4363) );
  OAI22_X1 U7199 ( .A1(n8715), .A2(n14579), .B1(n8713), .B2(n14609), .ZN(n4366) );
  OAI22_X1 U7200 ( .A1(n9738), .A2(n14387), .B1(n9743), .B2(n14535), .ZN(n4371) );
  OAI22_X1 U7201 ( .A1(n9739), .A2(n14579), .B1(n9737), .B2(n14609), .ZN(n4374) );
  OAI22_X1 U7202 ( .A1(n6666), .A2(n14387), .B1(n6671), .B2(n14535), .ZN(n4379) );
  OAI22_X1 U7203 ( .A1(n6667), .A2(n14579), .B1(n6665), .B2(n14609), .ZN(n4382) );
  OAI22_X1 U7204 ( .A1(n7690), .A2(n14387), .B1(n7695), .B2(n14535), .ZN(n4387) );
  OAI22_X1 U7205 ( .A1(n7691), .A2(n14579), .B1(n7689), .B2(n14609), .ZN(n4390) );
  OAI22_X1 U7206 ( .A1(n8210), .A2(n14387), .B1(n8215), .B2(n14535), .ZN(n4399) );
  OAI22_X1 U7207 ( .A1(n8211), .A2(n14579), .B1(n8209), .B2(n14609), .ZN(n4402) );
  OAI22_X1 U7208 ( .A1(n9234), .A2(n14387), .B1(n9239), .B2(n14535), .ZN(n4407) );
  OAI22_X1 U7209 ( .A1(n9235), .A2(n14579), .B1(n9233), .B2(n14609), .ZN(n4410) );
  OAI22_X1 U7210 ( .A1(n6162), .A2(n14387), .B1(n6167), .B2(n14535), .ZN(n4415) );
  OAI22_X1 U7211 ( .A1(n6163), .A2(n14579), .B1(n6161), .B2(n14609), .ZN(n4418) );
  OAI22_X1 U7212 ( .A1(n7186), .A2(n14387), .B1(n7191), .B2(n14535), .ZN(n4423) );
  OAI22_X1 U7213 ( .A1(n7187), .A2(n14579), .B1(n7185), .B2(n14608), .ZN(n4426) );
  OAI22_X1 U7214 ( .A1(n8722), .A2(n14387), .B1(n8727), .B2(n14535), .ZN(n4435) );
  OAI22_X1 U7215 ( .A1(n8723), .A2(n14579), .B1(n8721), .B2(n14608), .ZN(n4438) );
  OAI22_X1 U7216 ( .A1(n9746), .A2(n14388), .B1(n9751), .B2(n14536), .ZN(n4443) );
  OAI22_X1 U7217 ( .A1(n9747), .A2(n14580), .B1(n9745), .B2(n14608), .ZN(n4446) );
  OAI22_X1 U7218 ( .A1(n6674), .A2(n14388), .B1(n6679), .B2(n14536), .ZN(n4451) );
  OAI22_X1 U7219 ( .A1(n6675), .A2(n14580), .B1(n6673), .B2(n14608), .ZN(n4454) );
  OAI22_X1 U7220 ( .A1(n7698), .A2(n14388), .B1(n7703), .B2(n14536), .ZN(n4459) );
  OAI22_X1 U7221 ( .A1(n7699), .A2(n14580), .B1(n7697), .B2(n14608), .ZN(n4462) );
  OAI22_X1 U7222 ( .A1(n8186), .A2(n14388), .B1(n8191), .B2(n14536), .ZN(n4476) );
  OAI22_X1 U7223 ( .A1(n8187), .A2(n14580), .B1(n8185), .B2(n14608), .ZN(n4479) );
  OAI22_X1 U7224 ( .A1(n8698), .A2(n14388), .B1(n8703), .B2(n14536), .ZN(n4512) );
  OAI22_X1 U7225 ( .A1(n8699), .A2(n14580), .B1(n8697), .B2(n14608), .ZN(n4515) );
  OAI22_X1 U7226 ( .A1(n9722), .A2(n14388), .B1(n9727), .B2(n14536), .ZN(n4520) );
  OAI22_X1 U7227 ( .A1(n9723), .A2(n14580), .B1(n9721), .B2(n14608), .ZN(n4523) );
  OAI22_X1 U7228 ( .A1(n6650), .A2(n14388), .B1(n6655), .B2(n14536), .ZN(n4528) );
  OAI22_X1 U7229 ( .A1(n6651), .A2(n14580), .B1(n6649), .B2(n14608), .ZN(n4531) );
  OAI22_X1 U7230 ( .A1(n7674), .A2(n14388), .B1(n7679), .B2(n14536), .ZN(n4536) );
  OAI22_X1 U7231 ( .A1(n7675), .A2(n14580), .B1(n7673), .B2(n14608), .ZN(n4539) );
  OAI22_X1 U7232 ( .A1(n8194), .A2(n14388), .B1(n8199), .B2(n14536), .ZN(n4548) );
  OAI22_X1 U7233 ( .A1(n8195), .A2(n14580), .B1(n8193), .B2(n14607), .ZN(n4551) );
  OAI22_X1 U7234 ( .A1(n9218), .A2(n14388), .B1(n9223), .B2(n14536), .ZN(n4556) );
  OAI22_X1 U7235 ( .A1(n9219), .A2(n14580), .B1(n9217), .B2(n14607), .ZN(n4559) );
  OAI22_X1 U7236 ( .A1(n6146), .A2(n14389), .B1(n6151), .B2(n14537), .ZN(n4564) );
  OAI22_X1 U7237 ( .A1(n6147), .A2(n14581), .B1(n6145), .B2(n14607), .ZN(n4567) );
  OAI22_X1 U7238 ( .A1(n7170), .A2(n14389), .B1(n7175), .B2(n14537), .ZN(n4572) );
  OAI22_X1 U7239 ( .A1(n7171), .A2(n14581), .B1(n7169), .B2(n14607), .ZN(n4575) );
  OAI22_X1 U7240 ( .A1(n8706), .A2(n14389), .B1(n8711), .B2(n14537), .ZN(n4584) );
  OAI22_X1 U7241 ( .A1(n8707), .A2(n14581), .B1(n8705), .B2(n14607), .ZN(n4587) );
  OAI22_X1 U7242 ( .A1(n9730), .A2(n14389), .B1(n9735), .B2(n14537), .ZN(n4592) );
  OAI22_X1 U7243 ( .A1(n9731), .A2(n14581), .B1(n9729), .B2(n14607), .ZN(n4595) );
  OAI22_X1 U7244 ( .A1(n6658), .A2(n14389), .B1(n6663), .B2(n14537), .ZN(n4600) );
  OAI22_X1 U7245 ( .A1(n6659), .A2(n14581), .B1(n6657), .B2(n14607), .ZN(n4603) );
  OAI22_X1 U7246 ( .A1(n7682), .A2(n14389), .B1(n7687), .B2(n14537), .ZN(n4608) );
  OAI22_X1 U7247 ( .A1(n7683), .A2(n14581), .B1(n7681), .B2(n14607), .ZN(n4611) );
  OAI22_X1 U7248 ( .A1(n8170), .A2(n14389), .B1(n8175), .B2(n14537), .ZN(n4625) );
  OAI22_X1 U7249 ( .A1(n8171), .A2(n14581), .B1(n8169), .B2(n14607), .ZN(n4628) );
  OAI22_X1 U7250 ( .A1(n8682), .A2(n14389), .B1(n8687), .B2(n14537), .ZN(n4661) );
  OAI22_X1 U7251 ( .A1(n8683), .A2(n14581), .B1(n8681), .B2(n14607), .ZN(n4664) );
  OAI22_X1 U7252 ( .A1(n9706), .A2(n14389), .B1(n9711), .B2(n14537), .ZN(n4669) );
  OAI22_X1 U7253 ( .A1(n9707), .A2(n14581), .B1(n9705), .B2(n14606), .ZN(n4672) );
  OAI22_X1 U7254 ( .A1(n6634), .A2(n14389), .B1(n6639), .B2(n14537), .ZN(n4677) );
  OAI22_X1 U7255 ( .A1(n6635), .A2(n14581), .B1(n6633), .B2(n14606), .ZN(n4680) );
  OAI22_X1 U7256 ( .A1(n7658), .A2(n14390), .B1(n7663), .B2(n14538), .ZN(n4685) );
  OAI22_X1 U7257 ( .A1(n7659), .A2(n14582), .B1(n7657), .B2(n14606), .ZN(n4688) );
  OAI22_X1 U7258 ( .A1(n8178), .A2(n14390), .B1(n8183), .B2(n14538), .ZN(n4697) );
  OAI22_X1 U7259 ( .A1(n8179), .A2(n14582), .B1(n8177), .B2(n14606), .ZN(n4700) );
  OAI22_X1 U7260 ( .A1(n9202), .A2(n14390), .B1(n9207), .B2(n14538), .ZN(n4705) );
  OAI22_X1 U7261 ( .A1(n9203), .A2(n14582), .B1(n9201), .B2(n14606), .ZN(n4708) );
  OAI22_X1 U7262 ( .A1(n6130), .A2(n14390), .B1(n6135), .B2(n14538), .ZN(n4713) );
  OAI22_X1 U7263 ( .A1(n6131), .A2(n14582), .B1(n6129), .B2(n14606), .ZN(n4716) );
  OAI22_X1 U7264 ( .A1(n7154), .A2(n14390), .B1(n7159), .B2(n14538), .ZN(n4721) );
  OAI22_X1 U7265 ( .A1(n7155), .A2(n14582), .B1(n7153), .B2(n14606), .ZN(n4724) );
  OAI22_X1 U7266 ( .A1(n8690), .A2(n14390), .B1(n8695), .B2(n14538), .ZN(n4733) );
  OAI22_X1 U7267 ( .A1(n8691), .A2(n14582), .B1(n8689), .B2(n14606), .ZN(n4736) );
  OAI22_X1 U7268 ( .A1(n9714), .A2(n14390), .B1(n9719), .B2(n14538), .ZN(n4741) );
  OAI22_X1 U7269 ( .A1(n9715), .A2(n14582), .B1(n9713), .B2(n14606), .ZN(n4744) );
  OAI22_X1 U7270 ( .A1(n6642), .A2(n14390), .B1(n6647), .B2(n14538), .ZN(n4749) );
  OAI22_X1 U7271 ( .A1(n6643), .A2(n14582), .B1(n6641), .B2(n14606), .ZN(n4752) );
  OAI22_X1 U7272 ( .A1(n7666), .A2(n14390), .B1(n7671), .B2(n14538), .ZN(n4757) );
  OAI22_X1 U7273 ( .A1(n7667), .A2(n14582), .B1(n7665), .B2(n14611), .ZN(n4760) );
  OAI22_X1 U7274 ( .A1(n8154), .A2(n14390), .B1(n8159), .B2(n14538), .ZN(n4774) );
  OAI22_X1 U7275 ( .A1(n8155), .A2(n14582), .B1(n8153), .B2(n14625), .ZN(n4777) );
  OAI22_X1 U7276 ( .A1(n8666), .A2(n14391), .B1(n8671), .B2(n14539), .ZN(n4810) );
  OAI22_X1 U7277 ( .A1(n8667), .A2(n14583), .B1(n8665), .B2(n14625), .ZN(n4813) );
  OAI22_X1 U7278 ( .A1(n9690), .A2(n14391), .B1(n9695), .B2(n14539), .ZN(n4818) );
  OAI22_X1 U7279 ( .A1(n9691), .A2(n14583), .B1(n9689), .B2(n14625), .ZN(n4821) );
  OAI22_X1 U7280 ( .A1(n6618), .A2(n14391), .B1(n6623), .B2(n14539), .ZN(n4826) );
  OAI22_X1 U7281 ( .A1(n6619), .A2(n14583), .B1(n6617), .B2(n14625), .ZN(n4829) );
  OAI22_X1 U7282 ( .A1(n7642), .A2(n14391), .B1(n7647), .B2(n14539), .ZN(n4834) );
  OAI22_X1 U7283 ( .A1(n7643), .A2(n14583), .B1(n7641), .B2(n14625), .ZN(n4837) );
  OAI22_X1 U7284 ( .A1(n8162), .A2(n14391), .B1(n8167), .B2(n14539), .ZN(n4846) );
  OAI22_X1 U7285 ( .A1(n8163), .A2(n14583), .B1(n8161), .B2(n14625), .ZN(n4849) );
  OAI22_X1 U7286 ( .A1(n9186), .A2(n14391), .B1(n9191), .B2(n14539), .ZN(n4854) );
  OAI22_X1 U7287 ( .A1(n9187), .A2(n14583), .B1(n9185), .B2(n14625), .ZN(n4857) );
  OAI22_X1 U7288 ( .A1(n6114), .A2(n14391), .B1(n6119), .B2(n14539), .ZN(n4862) );
  OAI22_X1 U7289 ( .A1(n6115), .A2(n14583), .B1(n6113), .B2(n14625), .ZN(n4865) );
  OAI22_X1 U7290 ( .A1(n7138), .A2(n14391), .B1(n7143), .B2(n14539), .ZN(n4870) );
  OAI22_X1 U7291 ( .A1(n7139), .A2(n14583), .B1(n7137), .B2(n14624), .ZN(n4873) );
  OAI22_X1 U7292 ( .A1(n8674), .A2(n14391), .B1(n8679), .B2(n14539), .ZN(n4882) );
  OAI22_X1 U7293 ( .A1(n8675), .A2(n14583), .B1(n8673), .B2(n14624), .ZN(n4885) );
  OAI22_X1 U7294 ( .A1(n9698), .A2(n14391), .B1(n9703), .B2(n14539), .ZN(n4890) );
  OAI22_X1 U7295 ( .A1(n9699), .A2(n14583), .B1(n9697), .B2(n14624), .ZN(n4893) );
  OAI22_X1 U7296 ( .A1(n6626), .A2(n14391), .B1(n6631), .B2(n14539), .ZN(n4898) );
  OAI22_X1 U7297 ( .A1(n6627), .A2(n14583), .B1(n6625), .B2(n14624), .ZN(n4901) );
  OAI22_X1 U7298 ( .A1(n7650), .A2(n14391), .B1(n7655), .B2(n14539), .ZN(n4906) );
  OAI22_X1 U7299 ( .A1(n7651), .A2(n14583), .B1(n7649), .B2(n14624), .ZN(n4909) );
  OAI22_X1 U7300 ( .A1(n8138), .A2(n14391), .B1(n8143), .B2(n14539), .ZN(n4923) );
  OAI22_X1 U7301 ( .A1(n8139), .A2(n14583), .B1(n8137), .B2(n14624), .ZN(n4926) );
  OAI22_X1 U7302 ( .A1(n8650), .A2(n14392), .B1(n8655), .B2(n14540), .ZN(n4959) );
  OAI22_X1 U7303 ( .A1(n8651), .A2(n14584), .B1(n8649), .B2(n14624), .ZN(n4962) );
  OAI22_X1 U7304 ( .A1(n9674), .A2(n14392), .B1(n9679), .B2(n14540), .ZN(n4967) );
  OAI22_X1 U7305 ( .A1(n9675), .A2(n14584), .B1(n9673), .B2(n14624), .ZN(n4970) );
  OAI22_X1 U7306 ( .A1(n6602), .A2(n14392), .B1(n6607), .B2(n14540), .ZN(n4975) );
  OAI22_X1 U7307 ( .A1(n6603), .A2(n14584), .B1(n6601), .B2(n14624), .ZN(n4978) );
  OAI22_X1 U7308 ( .A1(n7626), .A2(n14392), .B1(n7631), .B2(n14540), .ZN(n4983) );
  OAI22_X1 U7309 ( .A1(n7627), .A2(n14584), .B1(n7625), .B2(n14624), .ZN(n4986) );
  OAI22_X1 U7310 ( .A1(n8146), .A2(n14392), .B1(n8151), .B2(n14540), .ZN(n4995) );
  OAI22_X1 U7311 ( .A1(n8147), .A2(n14584), .B1(n8145), .B2(n14623), .ZN(n4998) );
  OAI22_X1 U7313 ( .A1(n9170), .A2(n14392), .B1(n9175), .B2(n14540), .ZN(n5003) );
  OAI22_X1 U7314 ( .A1(n9171), .A2(n14584), .B1(n9169), .B2(n14623), .ZN(n5006) );
  OAI22_X1 U7315 ( .A1(n6098), .A2(n14392), .B1(n6103), .B2(n14540), .ZN(n5011) );
  OAI22_X1 U7316 ( .A1(n6099), .A2(n14584), .B1(n6097), .B2(n14623), .ZN(n5014) );
  OAI22_X1 U7317 ( .A1(n7122), .A2(n14392), .B1(n7127), .B2(n14540), .ZN(n5019) );
  OAI22_X1 U7318 ( .A1(n7123), .A2(n14584), .B1(n7121), .B2(n14623), .ZN(n5022) );
  OAI22_X1 U7319 ( .A1(n8658), .A2(n14392), .B1(n8663), .B2(n14540), .ZN(n5031) );
  OAI22_X1 U7320 ( .A1(n8659), .A2(n14584), .B1(n8657), .B2(n14623), .ZN(n5034) );
  OAI22_X1 U7321 ( .A1(n9682), .A2(n14392), .B1(n9687), .B2(n14540), .ZN(n5039) );
  OAI22_X1 U7322 ( .A1(n9683), .A2(n14584), .B1(n9681), .B2(n14623), .ZN(n5042) );
  OAI22_X1 U7323 ( .A1(n6610), .A2(n14393), .B1(n6615), .B2(n14541), .ZN(n5047) );
  OAI22_X1 U7324 ( .A1(n6611), .A2(n14585), .B1(n6609), .B2(n14623), .ZN(n5050) );
  OAI22_X1 U7325 ( .A1(n7634), .A2(n14393), .B1(n7639), .B2(n14541), .ZN(n5055) );
  OAI22_X1 U7326 ( .A1(n7635), .A2(n14585), .B1(n7633), .B2(n14623), .ZN(n5058) );
  OAI22_X1 U7327 ( .A1(n8122), .A2(n14393), .B1(n8127), .B2(n14541), .ZN(n5072) );
  OAI22_X1 U7328 ( .A1(n8123), .A2(n14585), .B1(n8121), .B2(n14623), .ZN(n5075) );
  OAI22_X1 U7329 ( .A1(n8634), .A2(n14393), .B1(n8639), .B2(n14541), .ZN(n5108) );
  OAI22_X1 U7330 ( .A1(n8635), .A2(n14585), .B1(n8633), .B2(n14623), .ZN(n5111) );
  OAI22_X1 U7331 ( .A1(n9658), .A2(n14393), .B1(n9663), .B2(n14541), .ZN(n5116) );
  OAI22_X1 U7332 ( .A1(n9659), .A2(n14585), .B1(n9657), .B2(n14622), .ZN(n5119) );
  OAI22_X1 U7333 ( .A1(n6586), .A2(n14393), .B1(n6591), .B2(n14541), .ZN(n5124) );
  OAI22_X1 U7334 ( .A1(n6587), .A2(n14585), .B1(n6585), .B2(n14622), .ZN(n5127) );
  OAI22_X1 U7335 ( .A1(n7610), .A2(n14393), .B1(n7615), .B2(n14541), .ZN(n5132) );
  OAI22_X1 U7336 ( .A1(n7611), .A2(n14585), .B1(n7609), .B2(n14622), .ZN(n5135) );
  OAI22_X1 U7337 ( .A1(n8130), .A2(n14393), .B1(n8135), .B2(n14541), .ZN(n5144) );
  OAI22_X1 U7338 ( .A1(n8131), .A2(n14585), .B1(n8129), .B2(n14622), .ZN(n5147) );
  OAI22_X1 U7339 ( .A1(n9154), .A2(n14393), .B1(n9159), .B2(n14541), .ZN(n5152) );
  OAI22_X1 U7340 ( .A1(n9155), .A2(n14585), .B1(n9153), .B2(n14622), .ZN(n5155) );
  OAI22_X1 U7341 ( .A1(n6082), .A2(n14393), .B1(n6087), .B2(n14541), .ZN(n5160) );
  OAI22_X1 U7342 ( .A1(n6083), .A2(n14585), .B1(n6081), .B2(n14622), .ZN(n5163) );
  OAI22_X1 U7343 ( .A1(n7106), .A2(n14394), .B1(n7111), .B2(n14542), .ZN(n5168) );
  OAI22_X1 U7344 ( .A1(n7107), .A2(n14586), .B1(n7105), .B2(n14622), .ZN(n5171) );
  OAI22_X1 U7345 ( .A1(n8642), .A2(n14394), .B1(n8647), .B2(n14542), .ZN(n5180) );
  OAI22_X1 U7346 ( .A1(n8643), .A2(n14586), .B1(n8641), .B2(n14622), .ZN(n5183) );
  OAI22_X1 U7347 ( .A1(n9666), .A2(n14394), .B1(n9671), .B2(n14542), .ZN(n5188) );
  OAI22_X1 U7348 ( .A1(n9667), .A2(n14586), .B1(n9665), .B2(n14622), .ZN(n5191) );
  OAI22_X1 U7349 ( .A1(n6594), .A2(n14394), .B1(n6599), .B2(n14542), .ZN(n5196) );
  OAI22_X1 U7350 ( .A1(n6595), .A2(n14586), .B1(n6593), .B2(n14622), .ZN(n5199) );
  OAI22_X1 U7351 ( .A1(n7618), .A2(n14394), .B1(n7623), .B2(n14542), .ZN(n5204) );
  OAI22_X1 U7352 ( .A1(n7619), .A2(n14586), .B1(n7617), .B2(n14622), .ZN(n5207) );
  OAI22_X1 U7353 ( .A1(n8106), .A2(n14394), .B1(n8111), .B2(n14542), .ZN(n5221) );
  OAI22_X1 U7354 ( .A1(n8107), .A2(n14586), .B1(n8105), .B2(n14622), .ZN(n5224) );
  OAI22_X1 U7355 ( .A1(n8618), .A2(n14394), .B1(n8623), .B2(n14542), .ZN(n5257) );
  OAI22_X1 U7356 ( .A1(n8619), .A2(n14586), .B1(n8617), .B2(n14621), .ZN(n5260) );
  OAI22_X1 U7357 ( .A1(n9642), .A2(n14394), .B1(n9647), .B2(n14542), .ZN(n5265) );
  OAI22_X1 U7358 ( .A1(n9643), .A2(n14586), .B1(n9641), .B2(n14621), .ZN(n5268) );
  OAI22_X1 U7359 ( .A1(n6570), .A2(n14394), .B1(n6575), .B2(n14542), .ZN(n5273) );
  OAI22_X1 U7360 ( .A1(n6571), .A2(n14586), .B1(n6569), .B2(n14621), .ZN(n5276) );
  OAI22_X1 U7361 ( .A1(n7594), .A2(n14394), .B1(n7599), .B2(n14542), .ZN(n5281) );
  OAI22_X1 U7362 ( .A1(n7595), .A2(n14586), .B1(n7593), .B2(n14621), .ZN(n5284) );
  OAI22_X1 U7363 ( .A1(n8114), .A2(n14395), .B1(n8119), .B2(n14543), .ZN(n5293) );
  OAI22_X1 U7364 ( .A1(n8115), .A2(n14587), .B1(n8113), .B2(n14621), .ZN(n5296) );
  OAI22_X1 U7365 ( .A1(n9138), .A2(n14395), .B1(n9143), .B2(n14543), .ZN(n5301) );
  OAI22_X1 U7366 ( .A1(n9139), .A2(n14587), .B1(n9137), .B2(n14621), .ZN(n5304) );
  OAI22_X1 U7367 ( .A1(n6066), .A2(n14395), .B1(n6071), .B2(n14543), .ZN(n5309) );
  OAI22_X1 U7368 ( .A1(n6067), .A2(n14587), .B1(n6065), .B2(n14621), .ZN(n5312) );
  OAI22_X1 U7369 ( .A1(n7090), .A2(n14395), .B1(n7095), .B2(n14543), .ZN(n5317) );
  OAI22_X1 U7370 ( .A1(n7091), .A2(n14587), .B1(n7089), .B2(n14621), .ZN(n5320) );
  OAI22_X1 U7371 ( .A1(n8626), .A2(n14395), .B1(n8631), .B2(n14543), .ZN(n5329) );
  OAI22_X1 U7372 ( .A1(n8627), .A2(n14587), .B1(n8625), .B2(n14621), .ZN(n5332) );
  OAI22_X1 U7373 ( .A1(n9650), .A2(n14395), .B1(n9655), .B2(n14543), .ZN(n5337) );
  OAI22_X1 U7374 ( .A1(n9651), .A2(n14587), .B1(n9649), .B2(n14621), .ZN(n5340) );
  OAI22_X1 U7375 ( .A1(n6578), .A2(n14395), .B1(n6583), .B2(n14543), .ZN(n5345) );
  OAI22_X1 U7376 ( .A1(n6579), .A2(n14587), .B1(n6577), .B2(n14621), .ZN(n5348) );
  OAI22_X1 U7377 ( .A1(n7602), .A2(n14395), .B1(n7607), .B2(n14543), .ZN(n5353) );
  OAI22_X1 U7378 ( .A1(n7603), .A2(n14587), .B1(n7601), .B2(n14620), .ZN(n5356) );
  OAI22_X1 U7379 ( .A1(n8090), .A2(n14395), .B1(n8095), .B2(n14543), .ZN(n5370) );
  OAI22_X1 U7380 ( .A1(n8091), .A2(n14587), .B1(n8089), .B2(n14620), .ZN(n5373) );
  OAI22_X1 U7381 ( .A1(n8602), .A2(n14395), .B1(n8607), .B2(n14543), .ZN(n5406) );
  OAI22_X1 U7382 ( .A1(n8603), .A2(n14587), .B1(n8601), .B2(n14620), .ZN(n5409) );
  OAI22_X1 U7383 ( .A1(n9626), .A2(n14396), .B1(n9631), .B2(n14544), .ZN(n5414) );
  OAI22_X1 U7384 ( .A1(n9627), .A2(n14588), .B1(n9625), .B2(n14620), .ZN(n5417) );
  OAI22_X1 U7385 ( .A1(n6554), .A2(n14396), .B1(n6559), .B2(n14544), .ZN(n5422) );
  OAI22_X1 U7386 ( .A1(n6555), .A2(n14588), .B1(n6553), .B2(n14620), .ZN(n5425) );
  OAI22_X1 U7387 ( .A1(n7578), .A2(n14396), .B1(n7583), .B2(n14544), .ZN(n5430) );
  OAI22_X1 U7388 ( .A1(n7579), .A2(n14588), .B1(n7577), .B2(n14620), .ZN(n5433) );
  OAI22_X1 U7389 ( .A1(n8098), .A2(n14396), .B1(n8103), .B2(n14544), .ZN(n5442) );
  OAI22_X1 U7390 ( .A1(n8099), .A2(n14588), .B1(n8097), .B2(n14620), .ZN(n5445) );
  OAI22_X1 U7391 ( .A1(n9122), .A2(n14396), .B1(n9127), .B2(n14544), .ZN(n5450) );
  OAI22_X1 U7392 ( .A1(n9123), .A2(n14588), .B1(n9121), .B2(n14620), .ZN(n5453) );
  OAI22_X1 U7393 ( .A1(n6050), .A2(n14396), .B1(n6055), .B2(n14544), .ZN(n5458) );
  OAI22_X1 U7394 ( .A1(n6051), .A2(n14588), .B1(n6049), .B2(n14620), .ZN(n5461) );
  OAI22_X1 U7395 ( .A1(n7074), .A2(n14396), .B1(n7079), .B2(n14544), .ZN(n5466) );
  OAI22_X1 U7396 ( .A1(n7075), .A2(n14588), .B1(n7073), .B2(n14619), .ZN(n5469) );
  OAI22_X1 U7397 ( .A1(n8610), .A2(n14396), .B1(n8615), .B2(n14544), .ZN(n5478) );
  OAI22_X1 U7398 ( .A1(n8611), .A2(n14588), .B1(n8609), .B2(n14619), .ZN(n5481) );
  OAI22_X1 U7399 ( .A1(n9634), .A2(n14396), .B1(n9639), .B2(n14544), .ZN(n5486) );
  OAI22_X1 U7400 ( .A1(n9635), .A2(n14588), .B1(n9633), .B2(n14619), .ZN(n5489) );
  OAI22_X1 U7401 ( .A1(n6562), .A2(n14396), .B1(n6567), .B2(n14544), .ZN(n5494) );
  OAI22_X1 U7402 ( .A1(n6563), .A2(n14588), .B1(n6561), .B2(n14619), .ZN(n5497) );
  OAI22_X1 U7403 ( .A1(n7586), .A2(n14396), .B1(n7591), .B2(n14544), .ZN(n5502) );
  OAI22_X1 U7404 ( .A1(n7587), .A2(n14588), .B1(n7585), .B2(n14619), .ZN(n5505) );
  OAI22_X1 U7405 ( .A1(n8074), .A2(n14396), .B1(n8079), .B2(n14544), .ZN(n5519) );
  OAI22_X1 U7406 ( .A1(n8075), .A2(n14588), .B1(n8073), .B2(n14619), .ZN(n5522) );
  OAI22_X1 U7407 ( .A1(n8586), .A2(n14397), .B1(n8591), .B2(n14545), .ZN(n5555) );
  OAI22_X1 U7408 ( .A1(n8587), .A2(n14589), .B1(n8585), .B2(n14619), .ZN(n5558) );
  OAI22_X1 U7409 ( .A1(n9610), .A2(n14397), .B1(n9615), .B2(n14545), .ZN(n5563) );
  OAI22_X1 U7410 ( .A1(n9611), .A2(n14589), .B1(n9609), .B2(n14619), .ZN(n5566) );
  OAI22_X1 U7411 ( .A1(n6538), .A2(n14397), .B1(n6543), .B2(n14545), .ZN(n5571) );
  OAI22_X1 U7412 ( .A1(n6539), .A2(n14589), .B1(n6537), .B2(n14619), .ZN(n5574) );
  OAI22_X1 U7413 ( .A1(n7562), .A2(n14397), .B1(n7567), .B2(n14545), .ZN(n5579) );
  OAI22_X1 U7414 ( .A1(n7563), .A2(n14589), .B1(n7561), .B2(n14619), .ZN(n5582) );
  OAI22_X1 U7415 ( .A1(n8082), .A2(n14397), .B1(n8087), .B2(n14545), .ZN(n5591) );
  OAI22_X1 U7416 ( .A1(n8083), .A2(n14589), .B1(n8081), .B2(n14618), .ZN(n5594) );
  OAI22_X1 U7417 ( .A1(n9106), .A2(n14397), .B1(n9111), .B2(n14545), .ZN(n5599) );
  OAI22_X1 U7418 ( .A1(n9107), .A2(n14589), .B1(n9105), .B2(n14618), .ZN(n5602) );
  OAI22_X1 U7419 ( .A1(n6034), .A2(n14397), .B1(n6039), .B2(n14545), .ZN(n5607) );
  OAI22_X1 U7420 ( .A1(n6035), .A2(n14589), .B1(n6033), .B2(n14618), .ZN(n5610) );
  OAI22_X1 U7421 ( .A1(n7058), .A2(n14397), .B1(n7063), .B2(n14545), .ZN(n5615) );
  OAI22_X1 U7422 ( .A1(n7059), .A2(n14589), .B1(n7057), .B2(n14618), .ZN(n5618) );
  OAI22_X1 U7423 ( .A1(n8594), .A2(n14397), .B1(n8599), .B2(n14545), .ZN(n5627) );
  OAI22_X1 U7424 ( .A1(n8595), .A2(n14589), .B1(n8593), .B2(n14618), .ZN(n5630) );
  OAI22_X1 U7425 ( .A1(n9618), .A2(n14397), .B1(n9623), .B2(n14545), .ZN(n5635) );
  OAI22_X1 U7426 ( .A1(n9619), .A2(n14589), .B1(n9617), .B2(n14618), .ZN(n5638) );
  OAI22_X1 U7427 ( .A1(n6546), .A2(n14397), .B1(n6551), .B2(n14545), .ZN(n5643) );
  OAI22_X1 U7428 ( .A1(n6547), .A2(n14589), .B1(n6545), .B2(n14618), .ZN(n5646) );
  OAI22_X1 U7429 ( .A1(n7570), .A2(n14398), .B1(n7575), .B2(n14546), .ZN(n5651) );
  OAI22_X1 U7430 ( .A1(n7571), .A2(n14590), .B1(n7569), .B2(n14618), .ZN(n5654) );
  OAI22_X1 U7431 ( .A1(n8058), .A2(n14398), .B1(n8063), .B2(n14546), .ZN(n5668) );
  OAI22_X1 U7432 ( .A1(n8059), .A2(n14590), .B1(n8057), .B2(n14618), .ZN(n5671) );
  OAI22_X1 U7433 ( .A1(n8570), .A2(n14398), .B1(n8575), .B2(n14546), .ZN(n5704) );
  OAI22_X1 U7434 ( .A1(n8571), .A2(n14590), .B1(n8569), .B2(n14618), .ZN(n5707) );
  OAI22_X1 U7435 ( .A1(n9594), .A2(n14398), .B1(n9599), .B2(n14546), .ZN(n5712) );
  OAI22_X1 U7436 ( .A1(n9595), .A2(n14590), .B1(n9593), .B2(n14617), .ZN(n5715) );
  OAI22_X1 U7437 ( .A1(n6522), .A2(n14398), .B1(n6527), .B2(n14546), .ZN(n5720) );
  OAI22_X1 U7438 ( .A1(n6523), .A2(n14590), .B1(n6521), .B2(n14617), .ZN(n5723) );
  OAI22_X1 U7439 ( .A1(n7546), .A2(n14398), .B1(n7551), .B2(n14546), .ZN(n5728) );
  OAI22_X1 U7440 ( .A1(n7547), .A2(n14590), .B1(n7545), .B2(n14617), .ZN(n5731) );
  OAI22_X1 U7441 ( .A1(n8066), .A2(n14398), .B1(n8071), .B2(n14546), .ZN(n5740) );
  OAI22_X1 U7442 ( .A1(n8067), .A2(n14590), .B1(n8065), .B2(n14617), .ZN(n5743) );
  OAI22_X1 U7443 ( .A1(n9090), .A2(n14398), .B1(n9095), .B2(n14546), .ZN(n5748) );
  OAI22_X1 U7444 ( .A1(n9091), .A2(n14590), .B1(n9089), .B2(n14617), .ZN(n5751) );
  OAI22_X1 U7445 ( .A1(n6018), .A2(n14398), .B1(n6023), .B2(n14546), .ZN(n5756) );
  OAI22_X1 U7446 ( .A1(n6019), .A2(n14590), .B1(n6017), .B2(n14617), .ZN(n5759) );
  OAI22_X1 U7447 ( .A1(n7042), .A2(n14398), .B1(n7047), .B2(n14546), .ZN(n5764) );
  OAI22_X1 U7448 ( .A1(n7043), .A2(n14590), .B1(n7041), .B2(n14617), .ZN(n5767) );
  OAI22_X1 U7449 ( .A1(n8578), .A2(n14399), .B1(n8583), .B2(n14547), .ZN(n5776) );
  OAI22_X1 U7450 ( .A1(n8579), .A2(n14591), .B1(n8577), .B2(n14617), .ZN(n5779) );
  OAI22_X1 U7451 ( .A1(n9602), .A2(n14399), .B1(n9607), .B2(n14547), .ZN(n5784) );
  OAI22_X1 U7452 ( .A1(n9603), .A2(n14591), .B1(n9601), .B2(n14617), .ZN(n5787) );
  OAI22_X1 U7453 ( .A1(n6530), .A2(n14399), .B1(n6535), .B2(n14547), .ZN(n5792) );
  OAI22_X1 U7454 ( .A1(n6531), .A2(n14591), .B1(n6529), .B2(n14617), .ZN(n5795) );
  OAI22_X1 U7455 ( .A1(n7554), .A2(n14399), .B1(n7559), .B2(n14547), .ZN(n5800) );
  OAI22_X1 U7456 ( .A1(n7555), .A2(n14591), .B1(n7553), .B2(n14617), .ZN(n5803) );
  OAI22_X1 U7457 ( .A1(n7018), .A2(n14399), .B1(n7023), .B2(n14547), .ZN(n5841) );
  OAI22_X1 U7458 ( .A1(n7019), .A2(n14591), .B1(n7017), .B2(n14616), .ZN(n5844) );
  OAI22_X1 U7459 ( .A1(n8554), .A2(n14399), .B1(n8559), .B2(n14547), .ZN(n5853) );
  OAI22_X1 U7460 ( .A1(n8555), .A2(n14591), .B1(n8553), .B2(n14616), .ZN(n5856) );
  OAI22_X1 U7461 ( .A1(n9578), .A2(n14399), .B1(n9583), .B2(n14547), .ZN(n5861) );
  OAI22_X1 U7462 ( .A1(n9579), .A2(n14591), .B1(n9577), .B2(n14616), .ZN(n5864) );
  OAI22_X1 U7463 ( .A1(n6506), .A2(n14399), .B1(n6511), .B2(n14547), .ZN(n5869) );
  OAI22_X1 U7465 ( .A1(n6507), .A2(n14591), .B1(n6505), .B2(n14616), .ZN(n5872) );
  OAI22_X1 U7466 ( .A1(n7530), .A2(n14399), .B1(n7535), .B2(n14547), .ZN(n5877) );
  OAI22_X1 U7467 ( .A1(n7531), .A2(n14591), .B1(n7529), .B2(n14616), .ZN(n5880) );
  OAI22_X1 U7468 ( .A1(n8050), .A2(n14399), .B1(n8055), .B2(n14547), .ZN(n5891) );
  OAI22_X1 U7469 ( .A1(n8051), .A2(n14591), .B1(n8049), .B2(n14616), .ZN(n5894) );
  OAI22_X1 U7470 ( .A1(n9075), .A2(n14592), .B1(n9073), .B2(n14616), .ZN(n5902) );
  OAI22_X1 U7471 ( .A1(n6003), .A2(n14592), .B1(n6001), .B2(n14616), .ZN(n5910) );
  OAI22_X1 U7472 ( .A1(n7027), .A2(n14592), .B1(n7025), .B2(n14616), .ZN(n5918) );
  OAI22_X1 U7473 ( .A1(n8563), .A2(n14592), .B1(n8561), .B2(n14616), .ZN(n5930) );
  OAI22_X1 U7474 ( .A1(n9587), .A2(n14592), .B1(n9585), .B2(n14616), .ZN(n5938) );
  OAI22_X1 U7475 ( .A1(n6515), .A2(n14592), .B1(n6513), .B2(n14620), .ZN(n5946) );
  OAI22_X1 U7476 ( .A1(n7539), .A2(n14592), .B1(n7537), .B2(n14625), .ZN(n5958) );
  AOI21_X1 U7477 ( .B1(n1178), .B2(n1179), .A(n14303), .ZN(n1177) );
  AOI221_X1 U7478 ( .B1(n14450), .B2(n3790), .C1(n14493), .C2(n1406), .A(n1186), .ZN(n1178) );
  AOI221_X1 U7479 ( .B1(n14351), .B2(n3792), .C1(n5816), .C2(n1408), .A(n1183), 
        .ZN(n1179) );
  AOI21_X1 U7480 ( .B1(n1218), .B2(n1219), .A(n14291), .ZN(n1217) );
  AOI221_X1 U7481 ( .B1(n14450), .B2(n3793), .C1(n14493), .C2(n1409), .A(n1226), .ZN(n1218) );
  AOI221_X1 U7482 ( .B1(n14351), .B2(n3801), .C1(n5851), .C2(n1417), .A(n1223), 
        .ZN(n1219) );
  AOI21_X1 U7483 ( .B1(n1258), .B2(n1259), .A(n5957), .ZN(n1257) );
  AOI221_X1 U7484 ( .B1(n14449), .B2(n3802), .C1(n14492), .C2(n1418), .A(n1266), .ZN(n1258) );
  AOI221_X1 U7485 ( .B1(n14350), .B2(n3804), .C1(n5801), .C2(n1420), .A(n1263), 
        .ZN(n1259) );
  AOI21_X1 U7486 ( .B1(n1298), .B2(n1299), .A(n5934), .ZN(n1297) );
  AOI221_X1 U7487 ( .B1(n14449), .B2(n3805), .C1(n14492), .C2(n1421), .A(n1306), .ZN(n1298) );
  AOI221_X1 U7488 ( .B1(n14350), .B2(n3809), .C1(n5801), .C2(n1425), .A(n1303), 
        .ZN(n1299) );
  AOI21_X1 U7489 ( .B1(n1343), .B2(n1344), .A(n14303), .ZN(n1342) );
  AOI221_X1 U7490 ( .B1(n14449), .B2(n3810), .C1(n14492), .C2(n1426), .A(n1350), .ZN(n1343) );
  AOI221_X1 U7491 ( .B1(n14350), .B2(n3812), .C1(n5799), .C2(n1428), .A(n1347), 
        .ZN(n1344) );
  AOI21_X1 U7492 ( .B1(n1379), .B2(n1380), .A(n14291), .ZN(n1378) );
  AOI221_X1 U7493 ( .B1(n14448), .B2(n3813), .C1(n14491), .C2(n1429), .A(n1386), .ZN(n1379) );
  AOI221_X1 U7494 ( .B1(n14349), .B2(n3817), .C1(n5802), .C2(n1433), .A(n1383), 
        .ZN(n1380) );
  AOI21_X1 U7495 ( .B1(n1415), .B2(n1416), .A(n5957), .ZN(n1414) );
  AOI221_X1 U7496 ( .B1(n14448), .B2(n3818), .C1(n14491), .C2(n1434), .A(n1422), .ZN(n1415) );
  AOI221_X1 U7497 ( .B1(n14349), .B2(n3820), .C1(n5802), .C2(n1436), .A(n1419), 
        .ZN(n1416) );
  AOI21_X1 U7498 ( .B1(n1451), .B2(n1452), .A(n5934), .ZN(n1450) );
  AOI221_X1 U7499 ( .B1(n14448), .B2(n3821), .C1(n14491), .C2(n1437), .A(n1458), .ZN(n1451) );
  AOI221_X1 U7500 ( .B1(n14349), .B2(n3825), .C1(n5801), .C2(n1441), .A(n1455), 
        .ZN(n1452) );
  AOI21_X1 U7501 ( .B1(n1492), .B2(n1493), .A(n14303), .ZN(n1491) );
  AOI221_X1 U7502 ( .B1(n14447), .B2(n3826), .C1(n14490), .C2(n1442), .A(n1499), .ZN(n1492) );
  AOI221_X1 U7503 ( .B1(n14348), .B2(n3828), .C1(n5801), .C2(n1444), .A(n1496), 
        .ZN(n1493) );
  AOI21_X1 U7504 ( .B1(n1528), .B2(n1529), .A(n14291), .ZN(n1527) );
  AOI221_X1 U7505 ( .B1(n14447), .B2(n3829), .C1(n14490), .C2(n1445), .A(n1535), .ZN(n1528) );
  AOI221_X1 U7506 ( .B1(n14348), .B2(n3837), .C1(n5815), .C2(n1453), .A(n1532), 
        .ZN(n1529) );
  AOI21_X1 U7507 ( .B1(n1564), .B2(n1565), .A(n5957), .ZN(n1563) );
  AOI221_X1 U7508 ( .B1(n14447), .B2(n3838), .C1(n14490), .C2(n1454), .A(n1571), .ZN(n1564) );
  AOI221_X1 U7509 ( .B1(n14348), .B2(n3840), .C1(n5802), .C2(n1456), .A(n1568), 
        .ZN(n1565) );
  AOI21_X1 U7510 ( .B1(n1600), .B2(n1601), .A(n5934), .ZN(n1599) );
  AOI221_X1 U7511 ( .B1(n14446), .B2(n3841), .C1(n14489), .C2(n1457), .A(n1607), .ZN(n1600) );
  AOI221_X1 U7512 ( .B1(n14347), .B2(n3845), .C1(n5802), .C2(n1461), .A(n1604), 
        .ZN(n1601) );
  AOI21_X1 U7513 ( .B1(n1641), .B2(n1642), .A(n14303), .ZN(n1640) );
  AOI221_X1 U7514 ( .B1(n14446), .B2(n3846), .C1(n14489), .C2(n1462), .A(n1648), .ZN(n1641) );
  AOI221_X1 U7515 ( .B1(n14347), .B2(n3848), .C1(n5816), .C2(n1464), .A(n1645), 
        .ZN(n1642) );
  AOI21_X1 U7516 ( .B1(n1677), .B2(n1678), .A(n14291), .ZN(n1676) );
  AOI221_X1 U7517 ( .B1(n14446), .B2(n3849), .C1(n14489), .C2(n1465), .A(n1684), .ZN(n1677) );
  AOI221_X1 U7518 ( .B1(n14347), .B2(n3853), .C1(n5816), .C2(n1469), .A(n1681), 
        .ZN(n1678) );
  AOI21_X1 U7519 ( .B1(n1713), .B2(n1714), .A(n5957), .ZN(n1712) );
  AOI221_X1 U7520 ( .B1(n14446), .B2(n3854), .C1(n14489), .C2(n1470), .A(n1720), .ZN(n1713) );
  AOI221_X1 U7521 ( .B1(n14347), .B2(n3856), .C1(n5815), .C2(n1472), .A(n1717), 
        .ZN(n1714) );
  AOI21_X1 U7522 ( .B1(n1749), .B2(n1750), .A(n5934), .ZN(n1748) );
  AOI221_X1 U7523 ( .B1(n14445), .B2(n3857), .C1(n14488), .C2(n1473), .A(n1756), .ZN(n1749) );
  AOI221_X1 U7524 ( .B1(n14346), .B2(n3861), .C1(n5818), .C2(n1477), .A(n1753), 
        .ZN(n1750) );
  AOI21_X1 U7525 ( .B1(n1790), .B2(n1791), .A(n14303), .ZN(n1789) );
  AOI221_X1 U7526 ( .B1(n14445), .B2(n3862), .C1(n14488), .C2(n1478), .A(n1797), .ZN(n1790) );
  AOI221_X1 U7527 ( .B1(n14346), .B2(n3864), .C1(n5818), .C2(n1480), .A(n1794), 
        .ZN(n1791) );
  AOI21_X1 U7528 ( .B1(n1826), .B2(n1827), .A(n14291), .ZN(n1825) );
  AOI221_X1 U7529 ( .B1(n14445), .B2(n3865), .C1(n14488), .C2(n1481), .A(n1833), .ZN(n1826) );
  AOI221_X1 U7530 ( .B1(n14346), .B2(n3878), .C1(n5816), .C2(n1494), .A(n1830), 
        .ZN(n1827) );
  AOI21_X1 U7531 ( .B1(n1862), .B2(n1863), .A(n5957), .ZN(n1861) );
  AOI221_X1 U7532 ( .B1(n14444), .B2(n3879), .C1(n14487), .C2(n1495), .A(n1869), .ZN(n1862) );
  AOI221_X1 U7533 ( .B1(n14345), .B2(n3881), .C1(n5819), .C2(n1497), .A(n1866), 
        .ZN(n1863) );
  AOI21_X1 U7534 ( .B1(n1898), .B2(n1899), .A(n5934), .ZN(n1897) );
  AOI221_X1 U7535 ( .B1(n14444), .B2(n3882), .C1(n14487), .C2(n1498), .A(n1905), .ZN(n1898) );
  AOI221_X1 U7536 ( .B1(n14345), .B2(n3886), .C1(n5819), .C2(n1502), .A(n1902), 
        .ZN(n1899) );
  AOI21_X1 U7537 ( .B1(n1939), .B2(n1940), .A(n14303), .ZN(n1938) );
  AOI221_X1 U7538 ( .B1(n14444), .B2(n3887), .C1(n14487), .C2(n1503), .A(n1946), .ZN(n1939) );
  AOI221_X1 U7539 ( .B1(n14345), .B2(n3889), .C1(n5818), .C2(n1505), .A(n1943), 
        .ZN(n1940) );
  AOI21_X1 U7540 ( .B1(n1975), .B2(n1976), .A(n14291), .ZN(n1974) );
  AOI221_X1 U7541 ( .B1(n14443), .B2(n3890), .C1(n14486), .C2(n1506), .A(n1982), .ZN(n1975) );
  AOI221_X1 U7542 ( .B1(n14344), .B2(n3894), .C1(n5818), .C2(n1510), .A(n1979), 
        .ZN(n1976) );
  AOI21_X1 U7543 ( .B1(n2011), .B2(n2012), .A(n5957), .ZN(n2010) );
  AOI221_X1 U7544 ( .B1(n14443), .B2(n3895), .C1(n14486), .C2(n1511), .A(n2018), .ZN(n2011) );
  AOI221_X1 U7545 ( .B1(n14344), .B2(n3897), .C1(n5823), .C2(n1513), .A(n2015), 
        .ZN(n2012) );
  AOI21_X1 U7546 ( .B1(n2047), .B2(n2048), .A(n5934), .ZN(n2046) );
  AOI221_X1 U7547 ( .B1(n14443), .B2(n3898), .C1(n14486), .C2(n1514), .A(n2054), .ZN(n2047) );
  AOI221_X1 U7548 ( .B1(n14344), .B2(n3902), .C1(n5823), .C2(n1518), .A(n2051), 
        .ZN(n2048) );
  AOI21_X1 U7549 ( .B1(n2088), .B2(n2089), .A(n14303), .ZN(n2087) );
  AOI221_X1 U7550 ( .B1(n14442), .B2(n3903), .C1(n14485), .C2(n1519), .A(n2095), .ZN(n2088) );
  AOI221_X1 U7551 ( .B1(n14343), .B2(n3905), .C1(n5819), .C2(n1521), .A(n2092), 
        .ZN(n2089) );
  AOI21_X1 U7552 ( .B1(n2124), .B2(n2125), .A(n14291), .ZN(n2123) );
  AOI221_X1 U7553 ( .B1(n14442), .B2(n3906), .C1(n14485), .C2(n1522), .A(n2131), .ZN(n2124) );
  AOI221_X1 U7554 ( .B1(n14343), .B2(n3914), .C1(n5824), .C2(n1530), .A(n2128), 
        .ZN(n2125) );
  AOI21_X1 U7555 ( .B1(n2160), .B2(n2161), .A(n5957), .ZN(n2159) );
  AOI221_X1 U7556 ( .B1(n14442), .B2(n3915), .C1(n14485), .C2(n1531), .A(n2167), .ZN(n2160) );
  AOI221_X1 U7557 ( .B1(n14343), .B2(n3917), .C1(n5824), .C2(n1533), .A(n2164), 
        .ZN(n2161) );
  AOI21_X1 U7558 ( .B1(n2196), .B2(n2197), .A(n5934), .ZN(n2195) );
  AOI221_X1 U7559 ( .B1(n14442), .B2(n3918), .C1(n14485), .C2(n1534), .A(n2203), .ZN(n2196) );
  AOI221_X1 U7560 ( .B1(n14343), .B2(n3922), .C1(n5823), .C2(n1538), .A(n2200), 
        .ZN(n2197) );
  AOI21_X1 U7561 ( .B1(n2237), .B2(n2238), .A(n14303), .ZN(n2236) );
  AOI221_X1 U7562 ( .B1(n14441), .B2(n3923), .C1(n14484), .C2(n1539), .A(n2244), .ZN(n2237) );
  AOI221_X1 U7563 ( .B1(n14342), .B2(n3925), .C1(n5826), .C2(n1541), .A(n2241), 
        .ZN(n2238) );
  AOI21_X1 U7564 ( .B1(n2273), .B2(n2274), .A(n14291), .ZN(n2272) );
  AOI221_X1 U7565 ( .B1(n14441), .B2(n3926), .C1(n14484), .C2(n1542), .A(n2280), .ZN(n2273) );
  AOI221_X1 U7566 ( .B1(n14342), .B2(n3930), .C1(n5826), .C2(n1546), .A(n2277), 
        .ZN(n2274) );
  AOI21_X1 U7567 ( .B1(n2309), .B2(n2310), .A(n5957), .ZN(n2308) );
  AOI221_X1 U7568 ( .B1(n14441), .B2(n3931), .C1(n14484), .C2(n1547), .A(n2316), .ZN(n2309) );
  AOI221_X1 U7569 ( .B1(n14342), .B2(n3933), .C1(n5824), .C2(n1549), .A(n2313), 
        .ZN(n2310) );
  AOI21_X1 U7570 ( .B1(n2345), .B2(n2346), .A(n5934), .ZN(n2344) );
  AOI221_X1 U7571 ( .B1(n14440), .B2(n3934), .C1(n14483), .C2(n1550), .A(n2352), .ZN(n2345) );
  AOI221_X1 U7572 ( .B1(n14341), .B2(n3938), .C1(n5871), .C2(n1554), .A(n2349), 
        .ZN(n2346) );
  AOI21_X1 U7573 ( .B1(n2386), .B2(n2387), .A(n14303), .ZN(n2385) );
  AOI221_X1 U7574 ( .B1(n14440), .B2(n3939), .C1(n14483), .C2(n1555), .A(n2393), .ZN(n2386) );
  AOI221_X1 U7575 ( .B1(n14341), .B2(n3941), .C1(n5827), .C2(n1557), .A(n2390), 
        .ZN(n2387) );
  AOI21_X1 U7576 ( .B1(n2422), .B2(n2423), .A(n14291), .ZN(n2421) );
  AOI221_X1 U7577 ( .B1(n14440), .B2(n3942), .C1(n14483), .C2(n1558), .A(n2429), .ZN(n2422) );
  AOI221_X1 U7578 ( .B1(n14341), .B2(n3950), .C1(n5835), .C2(n1566), .A(n2426), 
        .ZN(n2423) );
  AOI21_X1 U7579 ( .B1(n2458), .B2(n2459), .A(n5957), .ZN(n2457) );
  AOI221_X1 U7580 ( .B1(n14439), .B2(n3951), .C1(n14482), .C2(n1567), .A(n2465), .ZN(n2458) );
  AOI221_X1 U7581 ( .B1(n14340), .B2(n3953), .C1(n5827), .C2(n1569), .A(n2462), 
        .ZN(n2459) );
  AOI21_X1 U7582 ( .B1(n2494), .B2(n2495), .A(n5934), .ZN(n2493) );
  AOI221_X1 U7583 ( .B1(n14439), .B2(n3954), .C1(n14482), .C2(n1570), .A(n2501), .ZN(n2494) );
  AOI221_X1 U7584 ( .B1(n14340), .B2(n3958), .C1(n5827), .C2(n1574), .A(n2498), 
        .ZN(n2495) );
  AOI21_X1 U7585 ( .B1(n2535), .B2(n2536), .A(n14303), .ZN(n2534) );
  AOI221_X1 U7586 ( .B1(n14439), .B2(n3959), .C1(n14482), .C2(n1575), .A(n2542), .ZN(n2535) );
  AOI221_X1 U7587 ( .B1(n14340), .B2(n3961), .C1(n5827), .C2(n1577), .A(n2539), 
        .ZN(n2536) );
  AOI21_X1 U7588 ( .B1(n2571), .B2(n2572), .A(n14291), .ZN(n2570) );
  AOI221_X1 U7589 ( .B1(n14438), .B2(n3962), .C1(n14481), .C2(n1578), .A(n2578), .ZN(n2571) );
  AOI221_X1 U7590 ( .B1(n14339), .B2(n3966), .C1(n5832), .C2(n1582), .A(n2575), 
        .ZN(n2572) );
  AOI21_X1 U7591 ( .B1(n2607), .B2(n2608), .A(n5957), .ZN(n2606) );
  AOI221_X1 U7592 ( .B1(n14438), .B2(n3967), .C1(n14481), .C2(n1583), .A(n2614), .ZN(n2607) );
  AOI221_X1 U7593 ( .B1(n14339), .B2(n3969), .C1(n5831), .C2(n1585), .A(n2611), 
        .ZN(n2608) );
  AOI21_X1 U7594 ( .B1(n2643), .B2(n2644), .A(n5934), .ZN(n2642) );
  AOI221_X1 U7595 ( .B1(n14438), .B2(n3970), .C1(n14481), .C2(n1586), .A(n2650), .ZN(n2643) );
  AOI221_X1 U7596 ( .B1(n14339), .B2(n3974), .C1(n5831), .C2(n1590), .A(n2647), 
        .ZN(n2644) );
  AOI21_X1 U7597 ( .B1(n2684), .B2(n2685), .A(n14303), .ZN(n2683) );
  AOI221_X1 U7598 ( .B1(n14438), .B2(n3975), .C1(n14481), .C2(n1591), .A(n2691), .ZN(n2684) );
  AOI221_X1 U7599 ( .B1(n14339), .B2(n3977), .C1(n5834), .C2(n1593), .A(n2688), 
        .ZN(n2685) );
  AOI21_X1 U7600 ( .B1(n2720), .B2(n2721), .A(n14291), .ZN(n2719) );
  AOI221_X1 U7601 ( .B1(n14437), .B2(n3978), .C1(n14480), .C2(n1594), .A(n2727), .ZN(n2720) );
  AOI221_X1 U7602 ( .B1(n14338), .B2(n3986), .C1(n5832), .C2(n1602), .A(n2724), 
        .ZN(n2721) );
  AOI21_X1 U7603 ( .B1(n2756), .B2(n2757), .A(n5957), .ZN(n2755) );
  AOI221_X1 U7604 ( .B1(n14437), .B2(n3987), .C1(n14480), .C2(n1603), .A(n2763), .ZN(n2756) );
  AOI221_X1 U7605 ( .B1(n14338), .B2(n3989), .C1(n5832), .C2(n1605), .A(n2760), 
        .ZN(n2757) );
  AOI21_X1 U7606 ( .B1(n2792), .B2(n2793), .A(n5934), .ZN(n2791) );
  AOI221_X1 U7607 ( .B1(n14437), .B2(n3990), .C1(n14480), .C2(n1606), .A(n2799), .ZN(n2792) );
  AOI221_X1 U7608 ( .B1(n14338), .B2(n3994), .C1(n5832), .C2(n1610), .A(n2796), 
        .ZN(n2793) );
  AOI21_X1 U7609 ( .B1(n2833), .B2(n2834), .A(n14303), .ZN(n2832) );
  AOI221_X1 U7610 ( .B1(n14436), .B2(n3995), .C1(n14479), .C2(n1611), .A(n2840), .ZN(n2833) );
  AOI221_X1 U7611 ( .B1(n14337), .B2(n3997), .C1(n5834), .C2(n1613), .A(n2837), 
        .ZN(n2834) );
  AOI21_X1 U7612 ( .B1(n2869), .B2(n2870), .A(n14291), .ZN(n2868) );
  AOI221_X1 U7613 ( .B1(n14436), .B2(n3998), .C1(n14479), .C2(n1614), .A(n2876), .ZN(n2869) );
  AOI221_X1 U7614 ( .B1(n14337), .B2(n4002), .C1(n5834), .C2(n1618), .A(n2873), 
        .ZN(n2870) );
  AOI21_X1 U7615 ( .B1(n2905), .B2(n2906), .A(n5957), .ZN(n2904) );
  AOI221_X1 U7617 ( .B1(n14436), .B2(n4003), .C1(n14479), .C2(n1619), .A(n2912), .ZN(n2905) );
  AOI221_X1 U7618 ( .B1(n14337), .B2(n4005), .C1(n5834), .C2(n1621), .A(n2909), 
        .ZN(n2906) );
  AOI21_X1 U7619 ( .B1(n2941), .B2(n2942), .A(n5934), .ZN(n2940) );
  AOI221_X1 U7620 ( .B1(n14435), .B2(n4006), .C1(n14478), .C2(n1622), .A(n2948), .ZN(n2941) );
  AOI221_X1 U7621 ( .B1(n14336), .B2(n4010), .C1(n5839), .C2(n1626), .A(n2945), 
        .ZN(n2942) );
  AOI21_X1 U7622 ( .B1(n2982), .B2(n2983), .A(n14303), .ZN(n2981) );
  AOI221_X1 U7623 ( .B1(n14435), .B2(n4011), .C1(n14478), .C2(n1627), .A(n2989), .ZN(n2982) );
  AOI221_X1 U7624 ( .B1(n14336), .B2(n4013), .C1(n5835), .C2(n1629), .A(n2986), 
        .ZN(n2983) );
  AOI21_X1 U7625 ( .B1(n3018), .B2(n3019), .A(n14291), .ZN(n3017) );
  AOI221_X1 U7626 ( .B1(n14435), .B2(n4014), .C1(n14478), .C2(n1630), .A(n3025), .ZN(n3018) );
  AOI221_X1 U7627 ( .B1(n14336), .B2(n4027), .C1(n5835), .C2(n1643), .A(n3022), 
        .ZN(n3019) );
  AOI21_X1 U7628 ( .B1(n3054), .B2(n3055), .A(n5957), .ZN(n3053) );
  AOI221_X1 U7629 ( .B1(n14434), .B2(n4028), .C1(n14477), .C2(n1644), .A(n3061), .ZN(n3054) );
  AOI221_X1 U7630 ( .B1(n14335), .B2(n4030), .C1(n5839), .C2(n1646), .A(n3058), 
        .ZN(n3055) );
  AOI21_X1 U7631 ( .B1(n3090), .B2(n3091), .A(n5934), .ZN(n3089) );
  AOI221_X1 U7632 ( .B1(n14434), .B2(n4031), .C1(n14477), .C2(n1647), .A(n3097), .ZN(n3090) );
  AOI221_X1 U7633 ( .B1(n14335), .B2(n4035), .C1(n5839), .C2(n1651), .A(n3094), 
        .ZN(n3091) );
  AOI21_X1 U7634 ( .B1(n3131), .B2(n3132), .A(n14304), .ZN(n3130) );
  AOI221_X1 U7635 ( .B1(n14434), .B2(n4036), .C1(n14477), .C2(n1652), .A(n3138), .ZN(n3131) );
  AOI221_X1 U7636 ( .B1(n14335), .B2(n4038), .C1(n5839), .C2(n1654), .A(n3135), 
        .ZN(n3132) );
  AOI21_X1 U7637 ( .B1(n3167), .B2(n3168), .A(n14292), .ZN(n3166) );
  AOI221_X1 U7638 ( .B1(n14434), .B2(n4039), .C1(n14477), .C2(n1655), .A(n3174), .ZN(n3167) );
  AOI221_X1 U7639 ( .B1(n14335), .B2(n4043), .C1(n5842), .C2(n1659), .A(n3171), 
        .ZN(n3168) );
  AOI21_X1 U7640 ( .B1(n3203), .B2(n3204), .A(n14280), .ZN(n3202) );
  AOI221_X1 U7641 ( .B1(n14433), .B2(n4044), .C1(n14476), .C2(n1660), .A(n3210), .ZN(n3203) );
  AOI221_X1 U7642 ( .B1(n14334), .B2(n4046), .C1(n5840), .C2(n1662), .A(n3207), 
        .ZN(n3204) );
  AOI21_X1 U7643 ( .B1(n3239), .B2(n3240), .A(n5936), .ZN(n3238) );
  AOI221_X1 U7644 ( .B1(n14433), .B2(n4047), .C1(n14476), .C2(n1663), .A(n3246), .ZN(n3239) );
  AOI221_X1 U7645 ( .B1(n14334), .B2(n4051), .C1(n5840), .C2(n1667), .A(n3243), 
        .ZN(n3240) );
  AOI21_X1 U7646 ( .B1(n3280), .B2(n3281), .A(n14304), .ZN(n3279) );
  AOI221_X1 U7647 ( .B1(n14433), .B2(n4052), .C1(n14476), .C2(n1668), .A(n3287), .ZN(n3280) );
  AOI221_X1 U7648 ( .B1(n14334), .B2(n4054), .C1(n5843), .C2(n1670), .A(n3284), 
        .ZN(n3281) );
  AOI21_X1 U7649 ( .B1(n3316), .B2(n3317), .A(n14292), .ZN(n3315) );
  AOI221_X1 U7650 ( .B1(n14432), .B2(n4055), .C1(n14475), .C2(n1671), .A(n3323), .ZN(n3316) );
  AOI221_X1 U7651 ( .B1(n14333), .B2(n4063), .C1(n5842), .C2(n1679), .A(n3320), 
        .ZN(n3317) );
  AOI21_X1 U7652 ( .B1(n3352), .B2(n3353), .A(n14280), .ZN(n3351) );
  AOI221_X1 U7653 ( .B1(n14432), .B2(n4064), .C1(n14475), .C2(n1680), .A(n3359), .ZN(n3352) );
  AOI221_X1 U7654 ( .B1(n14333), .B2(n4066), .C1(n5842), .C2(n1682), .A(n3356), 
        .ZN(n3353) );
  AOI21_X1 U7655 ( .B1(n3388), .B2(n3389), .A(n5936), .ZN(n3387) );
  AOI221_X1 U7656 ( .B1(n14432), .B2(n4067), .C1(n14475), .C2(n1683), .A(n3395), .ZN(n3388) );
  AOI221_X1 U7657 ( .B1(n14333), .B2(n4071), .C1(n5851), .C2(n1687), .A(n3392), 
        .ZN(n3389) );
  AOI21_X1 U7658 ( .B1(n3429), .B2(n3430), .A(n14304), .ZN(n3428) );
  AOI221_X1 U7659 ( .B1(n14431), .B2(n4072), .C1(n14474), .C2(n1688), .A(n3436), .ZN(n3429) );
  AOI221_X1 U7660 ( .B1(n14332), .B2(n4074), .C1(n5843), .C2(n1690), .A(n3433), 
        .ZN(n3430) );
  AOI21_X1 U7661 ( .B1(n3465), .B2(n3466), .A(n14292), .ZN(n3464) );
  AOI221_X1 U7662 ( .B1(n14431), .B2(n4075), .C1(n14474), .C2(n1691), .A(n3472), .ZN(n3465) );
  AOI221_X1 U7663 ( .B1(n14332), .B2(n4079), .C1(n5843), .C2(n1695), .A(n3469), 
        .ZN(n3466) );
  AOI21_X1 U7664 ( .B1(n3501), .B2(n3502), .A(n14280), .ZN(n3500) );
  AOI221_X1 U7665 ( .B1(n14431), .B2(n4080), .C1(n14474), .C2(n1696), .A(n3508), .ZN(n3501) );
  AOI221_X1 U7666 ( .B1(n14332), .B2(n4082), .C1(n5843), .C2(n1698), .A(n3505), 
        .ZN(n3502) );
  AOI21_X1 U7667 ( .B1(n3537), .B2(n3538), .A(n5936), .ZN(n3536) );
  AOI221_X1 U7668 ( .B1(n14430), .B2(n4083), .C1(n14473), .C2(n1699), .A(n3544), .ZN(n3537) );
  AOI221_X1 U7669 ( .B1(n14331), .B2(n4087), .C1(n5799), .C2(n1703), .A(n3541), 
        .ZN(n3538) );
  AOI21_X1 U7670 ( .B1(n3578), .B2(n3579), .A(n14304), .ZN(n3577) );
  AOI221_X1 U7671 ( .B1(n14430), .B2(n4088), .C1(n14473), .C2(n1704), .A(n3585), .ZN(n3578) );
  AOI221_X1 U7672 ( .B1(n14331), .B2(n4090), .C1(n5852), .C2(n1706), .A(n3582), 
        .ZN(n3579) );
  AOI21_X1 U7673 ( .B1(n3614), .B2(n3615), .A(n14292), .ZN(n3613) );
  AOI221_X1 U7674 ( .B1(n14430), .B2(n4091), .C1(n14473), .C2(n1707), .A(n3621), .ZN(n3614) );
  AOI221_X1 U7675 ( .B1(n14331), .B2(n4099), .C1(n5852), .C2(n1715), .A(n3618), 
        .ZN(n3615) );
  AOI21_X1 U7676 ( .B1(n3650), .B2(n3651), .A(n14280), .ZN(n3649) );
  AOI221_X1 U7677 ( .B1(n14430), .B2(n4100), .C1(n14473), .C2(n1716), .A(n3657), .ZN(n3650) );
  AOI221_X1 U7678 ( .B1(n14331), .B2(n4102), .C1(n5851), .C2(n1718), .A(n3654), 
        .ZN(n3651) );
  AOI21_X1 U7679 ( .B1(n3686), .B2(n3687), .A(n5936), .ZN(n3685) );
  AOI221_X1 U7680 ( .B1(n14429), .B2(n4103), .C1(n14472), .C2(n1719), .A(n3693), .ZN(n3686) );
  AOI221_X1 U7681 ( .B1(n14330), .B2(n4107), .C1(n5854), .C2(n1723), .A(n3690), 
        .ZN(n3687) );
  AOI21_X1 U7682 ( .B1(n3727), .B2(n3728), .A(n14304), .ZN(n3726) );
  AOI221_X1 U7683 ( .B1(n14429), .B2(n4108), .C1(n14472), .C2(n1724), .A(n3734), .ZN(n3727) );
  AOI221_X1 U7684 ( .B1(n14330), .B2(n4110), .C1(n5854), .C2(n1726), .A(n3731), 
        .ZN(n3728) );
  AOI21_X1 U7685 ( .B1(n3763), .B2(n3764), .A(n14292), .ZN(n3762) );
  AOI221_X1 U7686 ( .B1(n14429), .B2(n4111), .C1(n14472), .C2(n1727), .A(n3770), .ZN(n3763) );
  AOI221_X1 U7687 ( .B1(n14330), .B2(n4115), .C1(n5852), .C2(n1731), .A(n3767), 
        .ZN(n3764) );
  AOI21_X1 U7688 ( .B1(n3799), .B2(n3800), .A(n14280), .ZN(n3798) );
  AOI221_X1 U7689 ( .B1(n14428), .B2(n4116), .C1(n14471), .C2(n1732), .A(n3806), .ZN(n3799) );
  AOI221_X1 U7690 ( .B1(n14329), .B2(n4118), .C1(n5855), .C2(n1734), .A(n3803), 
        .ZN(n3800) );
  AOI21_X1 U7691 ( .B1(n3835), .B2(n3836), .A(n5936), .ZN(n3834) );
  AOI221_X1 U7692 ( .B1(n14428), .B2(n4119), .C1(n14471), .C2(n1735), .A(n3842), .ZN(n3835) );
  AOI221_X1 U7693 ( .B1(n14329), .B2(n4123), .C1(n5855), .C2(n1739), .A(n3839), 
        .ZN(n3836) );
  AOI21_X1 U7694 ( .B1(n3876), .B2(n3877), .A(n14304), .ZN(n3875) );
  AOI221_X1 U7695 ( .B1(n14428), .B2(n4124), .C1(n14471), .C2(n1740), .A(n3883), .ZN(n3876) );
  AOI221_X1 U7696 ( .B1(n14329), .B2(n4126), .C1(n5854), .C2(n1742), .A(n3880), 
        .ZN(n3877) );
  AOI21_X1 U7697 ( .B1(n3912), .B2(n3913), .A(n14292), .ZN(n3911) );
  AOI221_X1 U7698 ( .B1(n14427), .B2(n4127), .C1(n14470), .C2(n1743), .A(n3919), .ZN(n3912) );
  AOI221_X1 U7699 ( .B1(n14328), .B2(n4135), .C1(n5854), .C2(n1751), .A(n3916), 
        .ZN(n3913) );
  AOI21_X1 U7700 ( .B1(n3948), .B2(n3949), .A(n14280), .ZN(n3947) );
  AOI221_X1 U7701 ( .B1(n14427), .B2(n4136), .C1(n14470), .C2(n1752), .A(n3955), .ZN(n3948) );
  AOI221_X1 U7702 ( .B1(n14328), .B2(n4138), .C1(n5859), .C2(n1754), .A(n3952), 
        .ZN(n3949) );
  AOI21_X1 U7703 ( .B1(n3984), .B2(n3985), .A(n5936), .ZN(n3983) );
  AOI221_X1 U7704 ( .B1(n14427), .B2(n4139), .C1(n14470), .C2(n1755), .A(n3991), .ZN(n3984) );
  AOI221_X1 U7705 ( .B1(n14328), .B2(n4143), .C1(n5859), .C2(n1759), .A(n3988), 
        .ZN(n3985) );
  AOI21_X1 U7706 ( .B1(n4025), .B2(n4026), .A(n14304), .ZN(n4024) );
  AOI221_X1 U7707 ( .B1(n14426), .B2(n4144), .C1(n14469), .C2(n1760), .A(n4032), .ZN(n4025) );
  AOI221_X1 U7708 ( .B1(n14327), .B2(n4146), .C1(n5855), .C2(n1762), .A(n4029), 
        .ZN(n4026) );
  AOI21_X1 U7709 ( .B1(n4061), .B2(n4062), .A(n14292), .ZN(n4060) );
  AOI221_X1 U7710 ( .B1(n14426), .B2(n4147), .C1(n14469), .C2(n1763), .A(n4068), .ZN(n4061) );
  AOI221_X1 U7711 ( .B1(n14327), .B2(n4151), .C1(n5860), .C2(n1767), .A(n4065), 
        .ZN(n4062) );
  AOI21_X1 U7712 ( .B1(n4097), .B2(n4098), .A(n14280), .ZN(n4096) );
  AOI221_X1 U7713 ( .B1(n14426), .B2(n4152), .C1(n14469), .C2(n1768), .A(n4104), .ZN(n4097) );
  AOI221_X1 U7714 ( .B1(n14327), .B2(n4154), .C1(n5860), .C2(n1770), .A(n4101), 
        .ZN(n4098) );
  AOI21_X1 U7715 ( .B1(n4133), .B2(n4134), .A(n5936), .ZN(n4132) );
  AOI221_X1 U7716 ( .B1(n14426), .B2(n4155), .C1(n14469), .C2(n1771), .A(n4140), .ZN(n4133) );
  AOI221_X1 U7717 ( .B1(n14327), .B2(n4159), .C1(n5859), .C2(n1775), .A(n4137), 
        .ZN(n4134) );
  AOI21_X1 U7718 ( .B1(n4174), .B2(n4175), .A(n14304), .ZN(n4173) );
  AOI221_X1 U7719 ( .B1(n14425), .B2(n4160), .C1(n14468), .C2(n1776), .A(n4181), .ZN(n4174) );
  AOI221_X1 U7720 ( .B1(n14326), .B2(n4162), .C1(n5862), .C2(n1778), .A(n4178), 
        .ZN(n4175) );
  AOI21_X1 U7721 ( .B1(n4210), .B2(n4211), .A(n14292), .ZN(n4209) );
  AOI221_X1 U7722 ( .B1(n14425), .B2(n4163), .C1(n14468), .C2(n1779), .A(n4217), .ZN(n4210) );
  AOI221_X1 U7723 ( .B1(n14326), .B2(n4176), .C1(n5862), .C2(n1792), .A(n4214), 
        .ZN(n4211) );
  AOI21_X1 U7724 ( .B1(n4246), .B2(n4247), .A(n14280), .ZN(n4245) );
  AOI221_X1 U7725 ( .B1(n14425), .B2(n4177), .C1(n14468), .C2(n1793), .A(n4253), .ZN(n4246) );
  AOI221_X1 U7726 ( .B1(n14326), .B2(n4179), .C1(n5860), .C2(n1795), .A(n4250), 
        .ZN(n4247) );
  AOI21_X1 U7727 ( .B1(n4282), .B2(n4283), .A(n5936), .ZN(n4281) );
  AOI221_X1 U7728 ( .B1(n14424), .B2(n4180), .C1(n14467), .C2(n1796), .A(n4289), .ZN(n4282) );
  AOI221_X1 U7729 ( .B1(n14325), .B2(n4184), .C1(n5863), .C2(n1800), .A(n4286), 
        .ZN(n4283) );
  AOI21_X1 U7730 ( .B1(n4323), .B2(n4324), .A(n14304), .ZN(n4322) );
  AOI221_X1 U7731 ( .B1(n14424), .B2(n4185), .C1(n14467), .C2(n1801), .A(n4330), .ZN(n4323) );
  AOI221_X1 U7732 ( .B1(n14325), .B2(n4187), .C1(n5863), .C2(n1803), .A(n4327), 
        .ZN(n4324) );
  AOI21_X1 U7733 ( .B1(n4359), .B2(n4360), .A(n14292), .ZN(n4358) );
  AOI221_X1 U7734 ( .B1(n14424), .B2(n4188), .C1(n14467), .C2(n1804), .A(n4366), .ZN(n4359) );
  AOI221_X1 U7735 ( .B1(n14325), .B2(n4192), .C1(n5862), .C2(n1808), .A(n4363), 
        .ZN(n4360) );
  AOI21_X1 U7736 ( .B1(n4395), .B2(n4396), .A(n14280), .ZN(n4394) );
  AOI221_X1 U7737 ( .B1(n14423), .B2(n4193), .C1(n14466), .C2(n1809), .A(n4402), .ZN(n4395) );
  AOI221_X1 U7738 ( .B1(n14324), .B2(n4195), .C1(n5867), .C2(n1811), .A(n4399), 
        .ZN(n4396) );
  AOI21_X1 U7739 ( .B1(n4431), .B2(n4432), .A(n5936), .ZN(n4430) );
  AOI221_X1 U7740 ( .B1(n14423), .B2(n4196), .C1(n14466), .C2(n1812), .A(n4438), .ZN(n4431) );
  AOI221_X1 U7741 ( .B1(n14324), .B2(n4200), .C1(n5867), .C2(n1816), .A(n4435), 
        .ZN(n4432) );
  AOI21_X1 U7742 ( .B1(n4472), .B2(n4473), .A(n14304), .ZN(n4471) );
  AOI221_X1 U7743 ( .B1(n14423), .B2(n4201), .C1(n14466), .C2(n1817), .A(n4479), .ZN(n4472) );
  AOI221_X1 U7744 ( .B1(n14324), .B2(n4203), .C1(n5867), .C2(n1819), .A(n4476), 
        .ZN(n4473) );
  AOI21_X1 U7745 ( .B1(n4508), .B2(n4509), .A(n14292), .ZN(n4507) );
  AOI221_X1 U7746 ( .B1(n14422), .B2(n4204), .C1(n14465), .C2(n1820), .A(n4515), .ZN(n4508) );
  AOI221_X1 U7747 ( .B1(n14323), .B2(n4212), .C1(n5863), .C2(n1828), .A(n4512), 
        .ZN(n4509) );
  AOI21_X1 U7748 ( .B1(n4544), .B2(n4545), .A(n14280), .ZN(n4543) );
  AOI221_X1 U7749 ( .B1(n14422), .B2(n4213), .C1(n14465), .C2(n1829), .A(n4551), .ZN(n4544) );
  AOI221_X1 U7750 ( .B1(n14323), .B2(n4215), .C1(n5868), .C2(n1831), .A(n4548), 
        .ZN(n4545) );
  AOI21_X1 U7751 ( .B1(n4580), .B2(n4581), .A(n5936), .ZN(n4579) );
  AOI221_X1 U7752 ( .B1(n14422), .B2(n4216), .C1(n14465), .C2(n1832), .A(n4587), .ZN(n4580) );
  AOI221_X1 U7753 ( .B1(n14323), .B2(n4220), .C1(n5868), .C2(n1836), .A(n4584), 
        .ZN(n4581) );
  AOI21_X1 U7754 ( .B1(n4621), .B2(n4622), .A(n14304), .ZN(n4620) );
  AOI221_X1 U7755 ( .B1(n14422), .B2(n4221), .C1(n14465), .C2(n1837), .A(n4628), .ZN(n4621) );
  AOI221_X1 U7756 ( .B1(n14323), .B2(n4223), .C1(n5867), .C2(n1839), .A(n4625), 
        .ZN(n4622) );
  AOI21_X1 U7757 ( .B1(n4657), .B2(n4658), .A(n14292), .ZN(n4656) );
  AOI221_X1 U7758 ( .B1(n14421), .B2(n4224), .C1(n14464), .C2(n1840), .A(n4664), .ZN(n4657) );
  AOI221_X1 U7759 ( .B1(n14322), .B2(n4228), .C1(n5870), .C2(n1844), .A(n4661), 
        .ZN(n4658) );
  AOI21_X1 U7760 ( .B1(n4693), .B2(n4694), .A(n14280), .ZN(n4692) );
  AOI221_X1 U7761 ( .B1(n14421), .B2(n4229), .C1(n14464), .C2(n1845), .A(n4700), .ZN(n4693) );
  AOI221_X1 U7762 ( .B1(n14322), .B2(n4231), .C1(n5870), .C2(n1847), .A(n4697), 
        .ZN(n4694) );
  AOI21_X1 U7763 ( .B1(n4729), .B2(n4730), .A(n5936), .ZN(n4728) );
  AOI221_X1 U7764 ( .B1(n14421), .B2(n4232), .C1(n14464), .C2(n1848), .A(n4736), .ZN(n4729) );
  AOI221_X1 U7765 ( .B1(n14322), .B2(n4236), .C1(n5868), .C2(n1852), .A(n4733), 
        .ZN(n4730) );
  AOI21_X1 U7766 ( .B1(n4770), .B2(n4771), .A(n14304), .ZN(n4769) );
  AOI221_X1 U7767 ( .B1(n14420), .B2(n4237), .C1(n14463), .C2(n1853), .A(n4777), .ZN(n4770) );
  AOI221_X1 U7769 ( .B1(n14321), .B2(n4239), .C1(n5870), .C2(n1855), .A(n4774), 
        .ZN(n4771) );
  AOI21_X1 U7770 ( .B1(n4806), .B2(n4807), .A(n14292), .ZN(n4805) );
  AOI221_X1 U7771 ( .B1(n14420), .B2(n4240), .C1(n14463), .C2(n1856), .A(n4813), .ZN(n4806) );
  AOI221_X1 U7772 ( .B1(n14321), .B2(n4248), .C1(n5826), .C2(n1864), .A(n4810), 
        .ZN(n4807) );
  AOI21_X1 U7773 ( .B1(n4842), .B2(n4843), .A(n14280), .ZN(n4841) );
  AOI221_X1 U7774 ( .B1(n14420), .B2(n4249), .C1(n14463), .C2(n1865), .A(n4849), .ZN(n4842) );
  AOI221_X1 U7775 ( .B1(n14321), .B2(n4251), .C1(n5875), .C2(n1867), .A(n4846), 
        .ZN(n4843) );
  AOI21_X1 U7776 ( .B1(n4878), .B2(n4879), .A(n5936), .ZN(n4877) );
  AOI221_X1 U7777 ( .B1(n14419), .B2(n4252), .C1(n14462), .C2(n1868), .A(n4885), .ZN(n4878) );
  AOI221_X1 U7778 ( .B1(n14320), .B2(n4256), .C1(n5871), .C2(n1872), .A(n4882), 
        .ZN(n4879) );
  AOI21_X1 U7779 ( .B1(n4919), .B2(n4920), .A(n14304), .ZN(n4918) );
  AOI221_X1 U7780 ( .B1(n14419), .B2(n4257), .C1(n14462), .C2(n1873), .A(n4926), .ZN(n4919) );
  AOI221_X1 U7781 ( .B1(n14320), .B2(n4259), .C1(n5871), .C2(n1875), .A(n4923), 
        .ZN(n4920) );
  AOI21_X1 U7782 ( .B1(n4955), .B2(n4956), .A(n14292), .ZN(n4954) );
  AOI221_X1 U7783 ( .B1(n14419), .B2(n4260), .C1(n14462), .C2(n1876), .A(n4962), .ZN(n4955) );
  AOI221_X1 U7784 ( .B1(n14320), .B2(n4264), .C1(n5871), .C2(n1880), .A(n4959), 
        .ZN(n4956) );
  AOI21_X1 U7785 ( .B1(n4991), .B2(n4992), .A(n14280), .ZN(n4990) );
  AOI221_X1 U7786 ( .B1(n14418), .B2(n4265), .C1(n14461), .C2(n1881), .A(n4998), .ZN(n4991) );
  AOI221_X1 U7787 ( .B1(n14319), .B2(n4267), .C1(n5875), .C2(n1883), .A(n4995), 
        .ZN(n4992) );
  AOI21_X1 U7788 ( .B1(n5027), .B2(n5028), .A(n5936), .ZN(n5026) );
  AOI221_X1 U7789 ( .B1(n14418), .B2(n4268), .C1(n14461), .C2(n1884), .A(n5034), .ZN(n5027) );
  AOI221_X1 U7790 ( .B1(n14319), .B2(n4272), .C1(n5875), .C2(n1888), .A(n5031), 
        .ZN(n5028) );
  AOI21_X1 U7791 ( .B1(n5068), .B2(n5069), .A(n14305), .ZN(n5067) );
  AOI221_X1 U7792 ( .B1(n14418), .B2(n4273), .C1(n14461), .C2(n1889), .A(n5075), .ZN(n5068) );
  AOI221_X1 U7793 ( .B1(n14319), .B2(n4275), .C1(n5875), .C2(n1891), .A(n5072), 
        .ZN(n5069) );
  AOI21_X1 U7794 ( .B1(n5104), .B2(n5105), .A(n14293), .ZN(n5103) );
  AOI221_X1 U7795 ( .B1(n14418), .B2(n4276), .C1(n14461), .C2(n1892), .A(n5111), .ZN(n5104) );
  AOI221_X1 U7796 ( .B1(n14319), .B2(n4284), .C1(n5878), .C2(n1900), .A(n5108), 
        .ZN(n5105) );
  AOI21_X1 U7797 ( .B1(n5140), .B2(n5141), .A(n14281), .ZN(n5139) );
  AOI221_X1 U7798 ( .B1(n14417), .B2(n4285), .C1(n14460), .C2(n1901), .A(n5147), .ZN(n5140) );
  AOI221_X1 U7799 ( .B1(n14318), .B2(n4287), .C1(n5876), .C2(n1903), .A(n5144), 
        .ZN(n5141) );
  AOI21_X1 U7800 ( .B1(n5176), .B2(n5177), .A(n5937), .ZN(n5175) );
  AOI221_X1 U7801 ( .B1(n14417), .B2(n4288), .C1(n14460), .C2(n1904), .A(n5183), .ZN(n5176) );
  AOI221_X1 U7802 ( .B1(n14318), .B2(n4292), .C1(n5876), .C2(n1908), .A(n5180), 
        .ZN(n5177) );
  AOI21_X1 U7803 ( .B1(n5217), .B2(n5218), .A(n14305), .ZN(n5216) );
  AOI221_X1 U7804 ( .B1(n14417), .B2(n4293), .C1(n14460), .C2(n1909), .A(n5224), .ZN(n5217) );
  AOI221_X1 U7805 ( .B1(n14318), .B2(n4295), .C1(n5879), .C2(n1911), .A(n5221), 
        .ZN(n5218) );
  AOI21_X1 U7806 ( .B1(n5253), .B2(n5254), .A(n14293), .ZN(n5252) );
  AOI221_X1 U7807 ( .B1(n14416), .B2(n4296), .C1(n14459), .C2(n1912), .A(n5260), .ZN(n5253) );
  AOI221_X1 U7808 ( .B1(n14317), .B2(n4300), .C1(n5878), .C2(n1916), .A(n5257), 
        .ZN(n5254) );
  AOI21_X1 U7809 ( .B1(n5289), .B2(n5290), .A(n14281), .ZN(n5288) );
  AOI221_X1 U7810 ( .B1(n14416), .B2(n4301), .C1(n14459), .C2(n1917), .A(n5296), .ZN(n5289) );
  AOI221_X1 U7811 ( .B1(n14317), .B2(n4303), .C1(n5878), .C2(n1919), .A(n5293), 
        .ZN(n5290) );
  AOI21_X1 U7812 ( .B1(n5325), .B2(n5326), .A(n5937), .ZN(n5324) );
  AOI221_X1 U7813 ( .B1(n14416), .B2(n4304), .C1(n14459), .C2(n1920), .A(n5332), .ZN(n5325) );
  AOI221_X1 U7814 ( .B1(n14317), .B2(n4308), .C1(n5889), .C2(n1924), .A(n5329), 
        .ZN(n5326) );
  AOI21_X1 U7815 ( .B1(n5366), .B2(n5367), .A(n14305), .ZN(n5365) );
  AOI221_X1 U7816 ( .B1(n14415), .B2(n4309), .C1(n14458), .C2(n1925), .A(n5373), .ZN(n5366) );
  AOI221_X1 U7817 ( .B1(n14316), .B2(n4311), .C1(n5879), .C2(n1927), .A(n5370), 
        .ZN(n5367) );
  AOI21_X1 U7818 ( .B1(n5402), .B2(n5403), .A(n14293), .ZN(n5401) );
  AOI221_X1 U7819 ( .B1(n14415), .B2(n4312), .C1(n14458), .C2(n1928), .A(n5409), .ZN(n5402) );
  AOI221_X1 U7820 ( .B1(n14316), .B2(n4325), .C1(n5879), .C2(n1941), .A(n5406), 
        .ZN(n5403) );
  AOI21_X1 U7821 ( .B1(n5438), .B2(n5439), .A(n14281), .ZN(n5437) );
  AOI221_X1 U7822 ( .B1(n14415), .B2(n4326), .C1(n14458), .C2(n1942), .A(n5445), .ZN(n5438) );
  AOI221_X1 U7823 ( .B1(n14316), .B2(n4328), .C1(n5890), .C2(n1944), .A(n5442), 
        .ZN(n5439) );
  AOI21_X1 U7824 ( .B1(n5474), .B2(n5475), .A(n5937), .ZN(n5473) );
  AOI221_X1 U7825 ( .B1(n14414), .B2(n4329), .C1(n14457), .C2(n1945), .A(n5481), .ZN(n5474) );
  AOI221_X1 U7826 ( .B1(n14315), .B2(n4333), .C1(n5889), .C2(n1949), .A(n5478), 
        .ZN(n5475) );
  AOI21_X1 U7827 ( .B1(n5515), .B2(n5516), .A(n14305), .ZN(n5514) );
  AOI221_X1 U7828 ( .B1(n14414), .B2(n4334), .C1(n14457), .C2(n1950), .A(n5522), .ZN(n5515) );
  AOI221_X1 U7829 ( .B1(n14315), .B2(n4336), .C1(n5889), .C2(n1952), .A(n5519), 
        .ZN(n5516) );
  AOI21_X1 U7830 ( .B1(n5551), .B2(n5552), .A(n14293), .ZN(n5550) );
  AOI221_X1 U7831 ( .B1(n14414), .B2(n4337), .C1(n14457), .C2(n1953), .A(n5558), .ZN(n5551) );
  AOI221_X1 U7832 ( .B1(n14315), .B2(n4341), .C1(n5889), .C2(n1957), .A(n5555), 
        .ZN(n5552) );
  AOI21_X1 U7833 ( .B1(n5587), .B2(n5588), .A(n14281), .ZN(n5586) );
  AOI221_X1 U7834 ( .B1(n14414), .B2(n4342), .C1(n14457), .C2(n1958), .A(n5594), .ZN(n5587) );
  AOI221_X1 U7835 ( .B1(n14315), .B2(n4344), .C1(n5892), .C2(n1960), .A(n5591), 
        .ZN(n5588) );
  AOI21_X1 U7836 ( .B1(n5623), .B2(n5624), .A(n5937), .ZN(n5622) );
  AOI221_X1 U7837 ( .B1(n14413), .B2(n4345), .C1(n14456), .C2(n1961), .A(n5630), .ZN(n5623) );
  AOI221_X1 U7838 ( .B1(n14314), .B2(n4349), .C1(n5890), .C2(n1965), .A(n5627), 
        .ZN(n5624) );
  AOI21_X1 U7839 ( .B1(n5664), .B2(n5665), .A(n14305), .ZN(n5663) );
  AOI221_X1 U7840 ( .B1(n14413), .B2(n4350), .C1(n14456), .C2(n1966), .A(n5671), .ZN(n5664) );
  AOI221_X1 U7841 ( .B1(n14314), .B2(n4352), .C1(n5890), .C2(n1968), .A(n5668), 
        .ZN(n5665) );
  AOI21_X1 U7842 ( .B1(n5700), .B2(n5701), .A(n14293), .ZN(n5699) );
  AOI221_X1 U7843 ( .B1(n14413), .B2(n4353), .C1(n14456), .C2(n1969), .A(n5707), .ZN(n5700) );
  AOI221_X1 U7844 ( .B1(n14314), .B2(n4361), .C1(n5893), .C2(n1977), .A(n5704), 
        .ZN(n5701) );
  AOI21_X1 U7845 ( .B1(n5736), .B2(n5737), .A(n14281), .ZN(n5735) );
  AOI221_X1 U7846 ( .B1(n14412), .B2(n4362), .C1(n14455), .C2(n1978), .A(n5743), .ZN(n5736) );
  AOI221_X1 U7847 ( .B1(n14313), .B2(n4364), .C1(n5892), .C2(n1980), .A(n5740), 
        .ZN(n5737) );
  AOI21_X1 U7848 ( .B1(n5772), .B2(n5773), .A(n5937), .ZN(n5771) );
  AOI221_X1 U7849 ( .B1(n14412), .B2(n4365), .C1(n14455), .C2(n1981), .A(n5779), .ZN(n5772) );
  AOI221_X1 U7850 ( .B1(n14313), .B2(n4369), .C1(n5892), .C2(n1985), .A(n5776), 
        .ZN(n5773) );
  AOI21_X1 U7851 ( .B1(n5849), .B2(n5850), .A(n14293), .ZN(n5848) );
  AOI221_X1 U7852 ( .B1(n14411), .B2(n4370), .C1(n14454), .C2(n1986), .A(n5856), .ZN(n5849) );
  AOI221_X1 U7853 ( .B1(n14312), .B2(n4372), .C1(n5893), .C2(n1988), .A(n5853), 
        .ZN(n5850) );
  AOI21_X1 U7854 ( .B1(n5885), .B2(n5886), .A(n14281), .ZN(n5884) );
  AOI221_X1 U7855 ( .B1(n14411), .B2(n4373), .C1(n14454), .C2(n1989), .A(n5894), .ZN(n5885) );
  AOI221_X1 U7856 ( .B1(n14312), .B2(n4377), .C1(n5893), .C2(n1993), .A(n5891), 
        .ZN(n5886) );
  AOI21_X1 U7857 ( .B1(n5923), .B2(n5924), .A(n5937), .ZN(n5922) );
  AOI221_X1 U7858 ( .B1(n14411), .B2(n4378), .C1(n14454), .C2(n1994), .A(n5930), .ZN(n5923) );
  AOI221_X1 U7859 ( .B1(n14312), .B2(n4380), .C1(n5852), .C2(n1996), .A(n5927), 
        .ZN(n5924) );
  AOI21_X1 U7860 ( .B1(n1227), .B2(n1228), .A(n14288), .ZN(n1216) );
  AOI221_X1 U7861 ( .B1(n14449), .B2(n4381), .C1(n14492), .C2(n1997), .A(n1235), .ZN(n1227) );
  AOI221_X1 U7862 ( .B1(n14350), .B2(n4385), .C1(n5851), .C2(n2001), .A(n1232), 
        .ZN(n1228) );
  AOI21_X1 U7863 ( .B1(n1267), .B2(n1268), .A(n5954), .ZN(n1256) );
  AOI221_X1 U7864 ( .B1(n14449), .B2(n4386), .C1(n14492), .C2(n2002), .A(n1275), .ZN(n1267) );
  AOI221_X1 U7865 ( .B1(n14350), .B2(n4388), .C1(n5801), .C2(n2004), .A(n1272), 
        .ZN(n1268) );
  AOI21_X1 U7866 ( .B1(n1307), .B2(n1308), .A(n5928), .ZN(n1296) );
  AOI221_X1 U7867 ( .B1(n14449), .B2(n4389), .C1(n14492), .C2(n2005), .A(n1315), .ZN(n1307) );
  AOI221_X1 U7868 ( .B1(n14350), .B2(n4397), .C1(n5801), .C2(n2013), .A(n1312), 
        .ZN(n1308) );
  AOI21_X1 U7869 ( .B1(n1387), .B2(n1388), .A(n14288), .ZN(n1377) );
  AOI221_X1 U7870 ( .B1(n14448), .B2(n4398), .C1(n14491), .C2(n2014), .A(n1394), .ZN(n1387) );
  AOI221_X1 U7871 ( .B1(n14349), .B2(n4400), .C1(n5802), .C2(n2016), .A(n1391), 
        .ZN(n1388) );
  AOI21_X1 U7872 ( .B1(n1423), .B2(n1424), .A(n5954), .ZN(n1413) );
  AOI221_X1 U7873 ( .B1(n14448), .B2(n4401), .C1(n14491), .C2(n2017), .A(n1430), .ZN(n1423) );
  AOI221_X1 U7874 ( .B1(n14349), .B2(n4405), .C1(n5802), .C2(n2021), .A(n1427), 
        .ZN(n1424) );
  AOI21_X1 U7875 ( .B1(n1459), .B2(n1460), .A(n5928), .ZN(n1449) );
  AOI221_X1 U7876 ( .B1(n14448), .B2(n4406), .C1(n14491), .C2(n2022), .A(n1466), .ZN(n1459) );
  AOI221_X1 U7877 ( .B1(n14349), .B2(n4408), .C1(n5801), .C2(n2024), .A(n1463), 
        .ZN(n1460) );
  AOI21_X1 U7878 ( .B1(n1536), .B2(n1537), .A(n14288), .ZN(n1526) );
  AOI221_X1 U7879 ( .B1(n14447), .B2(n4409), .C1(n14490), .C2(n2025), .A(n1543), .ZN(n1536) );
  AOI221_X1 U7880 ( .B1(n14348), .B2(n4413), .C1(n5815), .C2(n2029), .A(n1540), 
        .ZN(n1537) );
  AOI21_X1 U7881 ( .B1(n1572), .B2(n1573), .A(n5954), .ZN(n1562) );
  AOI221_X1 U7882 ( .B1(n14447), .B2(n4414), .C1(n14490), .C2(n2030), .A(n1579), .ZN(n1572) );
  AOI221_X1 U7883 ( .B1(n14348), .B2(n4416), .C1(n5802), .C2(n2032), .A(n1576), 
        .ZN(n1573) );
  AOI21_X1 U7884 ( .B1(n1608), .B2(n1609), .A(n5928), .ZN(n1598) );
  AOI221_X1 U7885 ( .B1(n14446), .B2(n4417), .C1(n14489), .C2(n2033), .A(n1615), .ZN(n1608) );
  AOI221_X1 U7886 ( .B1(n14347), .B2(n4421), .C1(n5802), .C2(n2037), .A(n1612), 
        .ZN(n1609) );
  AOI21_X1 U7887 ( .B1(n1685), .B2(n1686), .A(n14288), .ZN(n1675) );
  AOI221_X1 U7888 ( .B1(n14446), .B2(n4422), .C1(n14489), .C2(n2038), .A(n1692), .ZN(n1685) );
  AOI221_X1 U7889 ( .B1(n14347), .B2(n4424), .C1(n5815), .C2(n2040), .A(n1689), 
        .ZN(n1686) );
  AOI21_X1 U7890 ( .B1(n1721), .B2(n1722), .A(n5954), .ZN(n1711) );
  AOI221_X1 U7891 ( .B1(n14445), .B2(n4425), .C1(n14488), .C2(n2041), .A(n1728), .ZN(n1721) );
  AOI221_X1 U7892 ( .B1(n14346), .B2(n4433), .C1(n5815), .C2(n2049), .A(n1725), 
        .ZN(n1722) );
  AOI21_X1 U7893 ( .B1(n1757), .B2(n1758), .A(n5928), .ZN(n1747) );
  AOI221_X1 U7894 ( .B1(n14445), .B2(n4434), .C1(n14488), .C2(n2050), .A(n1764), .ZN(n1757) );
  AOI221_X1 U7895 ( .B1(n14346), .B2(n4436), .C1(n5818), .C2(n2052), .A(n1761), 
        .ZN(n1758) );
  AOI21_X1 U7896 ( .B1(n1834), .B2(n1835), .A(n14288), .ZN(n1824) );
  AOI221_X1 U7897 ( .B1(n14445), .B2(n4437), .C1(n14488), .C2(n2053), .A(n1841), .ZN(n1834) );
  AOI221_X1 U7898 ( .B1(n14346), .B2(n4441), .C1(n5816), .C2(n2057), .A(n1838), 
        .ZN(n1835) );
  AOI21_X1 U7899 ( .B1(n1870), .B2(n1871), .A(n5954), .ZN(n1860) );
  AOI221_X1 U7900 ( .B1(n14444), .B2(n4442), .C1(n14487), .C2(n2058), .A(n1877), .ZN(n1870) );
  AOI221_X1 U7901 ( .B1(n14345), .B2(n4444), .C1(n5819), .C2(n2060), .A(n1874), 
        .ZN(n1871) );
  AOI21_X1 U7902 ( .B1(n1906), .B2(n1907), .A(n5928), .ZN(n1896) );
  AOI221_X1 U7903 ( .B1(n14444), .B2(n4445), .C1(n14487), .C2(n2061), .A(n1913), .ZN(n1906) );
  AOI221_X1 U7904 ( .B1(n14345), .B2(n4449), .C1(n5819), .C2(n2065), .A(n1910), 
        .ZN(n1907) );
  AOI21_X1 U7905 ( .B1(n1983), .B2(n1984), .A(n14288), .ZN(n1973) );
  AOI221_X1 U7906 ( .B1(n14443), .B2(n4450), .C1(n14486), .C2(n2066), .A(n1990), .ZN(n1983) );
  AOI221_X1 U7907 ( .B1(n14344), .B2(n4452), .C1(n5823), .C2(n2068), .A(n1987), 
        .ZN(n1984) );
  AOI21_X1 U7908 ( .B1(n2019), .B2(n2020), .A(n5954), .ZN(n2009) );
  AOI221_X1 U7909 ( .B1(n14443), .B2(n4453), .C1(n14486), .C2(n2069), .A(n2026), .ZN(n2019) );
  AOI221_X1 U7910 ( .B1(n14344), .B2(n4457), .C1(n5823), .C2(n2073), .A(n2023), 
        .ZN(n2020) );
  AOI21_X1 U7911 ( .B1(n2055), .B2(n2056), .A(n5928), .ZN(n2045) );
  AOI221_X1 U7912 ( .B1(n14443), .B2(n4458), .C1(n14486), .C2(n2074), .A(n2062), .ZN(n2055) );
  AOI221_X1 U7913 ( .B1(n14344), .B2(n4460), .C1(n5819), .C2(n2076), .A(n2059), 
        .ZN(n2056) );
  AOI21_X1 U7914 ( .B1(n2132), .B2(n2133), .A(n14288), .ZN(n2122) );
  AOI221_X1 U7915 ( .B1(n14442), .B2(n4461), .C1(n14485), .C2(n2077), .A(n2139), .ZN(n2132) );
  AOI221_X1 U7916 ( .B1(n14343), .B2(n4474), .C1(n5824), .C2(n2090), .A(n2136), 
        .ZN(n2133) );
  AOI21_X1 U7917 ( .B1(n2168), .B2(n2169), .A(n5954), .ZN(n2158) );
  AOI221_X1 U7918 ( .B1(n14442), .B2(n4475), .C1(n14485), .C2(n2091), .A(n2175), .ZN(n2168) );
  AOI221_X1 U7919 ( .B1(n14343), .B2(n4477), .C1(n5824), .C2(n2093), .A(n2172), 
        .ZN(n2169) );
  AOI21_X1 U7921 ( .B1(n2204), .B2(n2205), .A(n5928), .ZN(n2194) );
  AOI221_X1 U7922 ( .B1(n14441), .B2(n4478), .C1(n14484), .C2(n2094), .A(n2211), .ZN(n2204) );
  AOI221_X1 U7923 ( .B1(n14342), .B2(n4482), .C1(n5823), .C2(n2098), .A(n2208), 
        .ZN(n2205) );
  AOI21_X1 U7924 ( .B1(n2281), .B2(n2282), .A(n14288), .ZN(n2271) );
  AOI221_X1 U7925 ( .B1(n14441), .B2(n4483), .C1(n14484), .C2(n2099), .A(n2288), .ZN(n2281) );
  AOI221_X1 U7926 ( .B1(n14342), .B2(n4485), .C1(n5826), .C2(n2101), .A(n2285), 
        .ZN(n2282) );
  AOI21_X1 U7927 ( .B1(n2317), .B2(n2318), .A(n5954), .ZN(n2307) );
  AOI221_X1 U7928 ( .B1(n14441), .B2(n4486), .C1(n14484), .C2(n2102), .A(n2324), .ZN(n2317) );
  AOI221_X1 U7929 ( .B1(n14342), .B2(n4490), .C1(n5824), .C2(n2106), .A(n2321), 
        .ZN(n2318) );
  AOI21_X1 U7930 ( .B1(n2353), .B2(n2354), .A(n5928), .ZN(n2343) );
  AOI221_X1 U7931 ( .B1(n14440), .B2(n4491), .C1(n14483), .C2(n2107), .A(n2360), .ZN(n2353) );
  AOI221_X1 U7932 ( .B1(n14341), .B2(n4493), .C1(n5871), .C2(n2109), .A(n2357), 
        .ZN(n2354) );
  AOI21_X1 U7933 ( .B1(n2430), .B2(n2431), .A(n14288), .ZN(n2420) );
  AOI221_X1 U7934 ( .B1(n14440), .B2(n4494), .C1(n14483), .C2(n2110), .A(n2437), .ZN(n2430) );
  AOI221_X1 U7935 ( .B1(n14341), .B2(n4498), .C1(n5831), .C2(n2114), .A(n2434), 
        .ZN(n2431) );
  AOI21_X1 U7936 ( .B1(n2466), .B2(n2467), .A(n5954), .ZN(n2456) );
  AOI221_X1 U7937 ( .B1(n14439), .B2(n4499), .C1(n14482), .C2(n2115), .A(n2473), .ZN(n2466) );
  AOI221_X1 U7938 ( .B1(n14340), .B2(n4501), .C1(n5827), .C2(n2117), .A(n2470), 
        .ZN(n2467) );
  AOI21_X1 U7939 ( .B1(n2502), .B2(n2503), .A(n5928), .ZN(n2492) );
  AOI221_X1 U7940 ( .B1(n14439), .B2(n4502), .C1(n14482), .C2(n2118), .A(n2509), .ZN(n2502) );
  AOI221_X1 U7941 ( .B1(n14340), .B2(n4510), .C1(n5827), .C2(n2126), .A(n2506), 
        .ZN(n2503) );
  AOI21_X1 U7942 ( .B1(n2579), .B2(n2580), .A(n14288), .ZN(n2569) );
  AOI221_X1 U7943 ( .B1(n14438), .B2(n4511), .C1(n14481), .C2(n2127), .A(n2586), .ZN(n2579) );
  AOI221_X1 U7944 ( .B1(n14339), .B2(n4513), .C1(n5831), .C2(n2129), .A(n2583), 
        .ZN(n2580) );
  AOI21_X1 U7945 ( .B1(n2615), .B2(n2616), .A(n5954), .ZN(n2605) );
  AOI221_X1 U7946 ( .B1(n14438), .B2(n4514), .C1(n14481), .C2(n2130), .A(n2622), .ZN(n2615) );
  AOI221_X1 U7947 ( .B1(n14339), .B2(n4518), .C1(n5831), .C2(n2134), .A(n2619), 
        .ZN(n2616) );
  AOI21_X1 U7948 ( .B1(n2651), .B2(n2652), .A(n5928), .ZN(n2641) );
  AOI221_X1 U7949 ( .B1(n14438), .B2(n4519), .C1(n14481), .C2(n2135), .A(n2658), .ZN(n2651) );
  AOI221_X1 U7950 ( .B1(n14339), .B2(n4521), .C1(n5831), .C2(n2137), .A(n2655), 
        .ZN(n2652) );
  AOI21_X1 U7951 ( .B1(n2728), .B2(n2729), .A(n14288), .ZN(n2718) );
  AOI221_X1 U7952 ( .B1(n14437), .B2(n4522), .C1(n14480), .C2(n2138), .A(n2735), .ZN(n2728) );
  AOI221_X1 U7953 ( .B1(n14338), .B2(n4526), .C1(n5832), .C2(n2142), .A(n2732), 
        .ZN(n2729) );
  AOI21_X1 U7954 ( .B1(n2764), .B2(n2765), .A(n5954), .ZN(n2754) );
  AOI221_X1 U7955 ( .B1(n14437), .B2(n4527), .C1(n14480), .C2(n2143), .A(n2771), .ZN(n2764) );
  AOI221_X1 U7956 ( .B1(n14338), .B2(n4529), .C1(n5832), .C2(n2145), .A(n2768), 
        .ZN(n2765) );
  AOI21_X1 U7957 ( .B1(n2800), .B2(n2801), .A(n5928), .ZN(n2790) );
  AOI221_X1 U7958 ( .B1(n14437), .B2(n4530), .C1(n14480), .C2(n2146), .A(n2807), .ZN(n2800) );
  AOI221_X1 U7959 ( .B1(n14338), .B2(n4534), .C1(n5834), .C2(n2150), .A(n2804), 
        .ZN(n2801) );
  AOI21_X1 U7960 ( .B1(n2877), .B2(n2878), .A(n14288), .ZN(n2867) );
  AOI221_X1 U7961 ( .B1(n14436), .B2(n4535), .C1(n14479), .C2(n2151), .A(n2884), .ZN(n2877) );
  AOI221_X1 U7962 ( .B1(n14337), .B2(n4537), .C1(n5834), .C2(n2153), .A(n2881), 
        .ZN(n2878) );
  AOI21_X1 U7963 ( .B1(n2913), .B2(n2914), .A(n5954), .ZN(n2903) );
  AOI221_X1 U7964 ( .B1(n14436), .B2(n4538), .C1(n14479), .C2(n2154), .A(n2920), .ZN(n2913) );
  AOI221_X1 U7965 ( .B1(n14337), .B2(n4546), .C1(n5839), .C2(n2162), .A(n2917), 
        .ZN(n2914) );
  AOI21_X1 U7966 ( .B1(n2949), .B2(n2950), .A(n5928), .ZN(n2939) );
  AOI221_X1 U7967 ( .B1(n14435), .B2(n4547), .C1(n14478), .C2(n2163), .A(n2956), .ZN(n2949) );
  AOI221_X1 U7968 ( .B1(n14336), .B2(n4549), .C1(n5835), .C2(n2165), .A(n2953), 
        .ZN(n2950) );
  AOI21_X1 U7969 ( .B1(n3026), .B2(n3027), .A(n14288), .ZN(n3016) );
  AOI221_X1 U7970 ( .B1(n14435), .B2(n4550), .C1(n14478), .C2(n2166), .A(n3033), .ZN(n3026) );
  AOI221_X1 U7971 ( .B1(n14336), .B2(n4554), .C1(n5840), .C2(n2170), .A(n3030), 
        .ZN(n3027) );
  AOI21_X1 U7972 ( .B1(n3062), .B2(n3063), .A(n5954), .ZN(n3052) );
  AOI221_X1 U7973 ( .B1(n14434), .B2(n4555), .C1(n14477), .C2(n2171), .A(n3069), .ZN(n3062) );
  AOI221_X1 U7974 ( .B1(n14335), .B2(n4557), .C1(n5839), .C2(n2173), .A(n3066), 
        .ZN(n3063) );
  AOI21_X1 U7975 ( .B1(n3098), .B2(n3099), .A(n5928), .ZN(n3088) );
  AOI221_X1 U7976 ( .B1(n14434), .B2(n4558), .C1(n14477), .C2(n2174), .A(n3105), .ZN(n3098) );
  AOI221_X1 U7977 ( .B1(n14335), .B2(n4562), .C1(n5839), .C2(n2178), .A(n3102), 
        .ZN(n3099) );
  AOI21_X1 U7978 ( .B1(n3175), .B2(n3176), .A(n14289), .ZN(n3165) );
  AOI221_X1 U7979 ( .B1(n14433), .B2(n4563), .C1(n14476), .C2(n2179), .A(n3182), .ZN(n3175) );
  AOI221_X1 U7980 ( .B1(n14334), .B2(n4565), .C1(n5840), .C2(n2181), .A(n3179), 
        .ZN(n3176) );
  AOI21_X1 U7981 ( .B1(n3211), .B2(n3212), .A(n5955), .ZN(n3201) );
  AOI221_X1 U7982 ( .B1(n14433), .B2(n4566), .C1(n14476), .C2(n2182), .A(n3218), .ZN(n3211) );
  AOI221_X1 U7983 ( .B1(n14334), .B2(n4570), .C1(n5840), .C2(n2186), .A(n3215), 
        .ZN(n3212) );
  AOI21_X1 U7984 ( .B1(n3247), .B2(n3248), .A(n5929), .ZN(n3237) );
  AOI221_X1 U7985 ( .B1(n14433), .B2(n4571), .C1(n14476), .C2(n2187), .A(n3254), .ZN(n3247) );
  AOI221_X1 U7986 ( .B1(n14334), .B2(n4573), .C1(n5840), .C2(n2189), .A(n3251), 
        .ZN(n3248) );
  AOI21_X1 U7987 ( .B1(n3324), .B2(n3325), .A(n14289), .ZN(n3314) );
  AOI221_X1 U7988 ( .B1(n14432), .B2(n4574), .C1(n14475), .C2(n2190), .A(n3331), .ZN(n3324) );
  AOI221_X1 U7989 ( .B1(n14333), .B2(n4582), .C1(n5842), .C2(n2198), .A(n3328), 
        .ZN(n3325) );
  AOI21_X1 U7990 ( .B1(n3360), .B2(n3361), .A(n5955), .ZN(n3350) );
  AOI221_X1 U7991 ( .B1(n14432), .B2(n4583), .C1(n14475), .C2(n2199), .A(n3367), .ZN(n3360) );
  AOI221_X1 U7992 ( .B1(n14333), .B2(n4585), .C1(n5842), .C2(n2201), .A(n3364), 
        .ZN(n3361) );
  AOI21_X1 U7993 ( .B1(n3396), .B2(n3397), .A(n5929), .ZN(n3386) );
  AOI221_X1 U7994 ( .B1(n14432), .B2(n4586), .C1(n14475), .C2(n2202), .A(n3403), .ZN(n3396) );
  AOI221_X1 U7995 ( .B1(n14333), .B2(n4590), .C1(n5851), .C2(n2206), .A(n3400), 
        .ZN(n3397) );
  AOI21_X1 U7996 ( .B1(n3473), .B2(n3474), .A(n14289), .ZN(n3463) );
  AOI221_X1 U7997 ( .B1(n14431), .B2(n4591), .C1(n14474), .C2(n2207), .A(n3480), .ZN(n3473) );
  AOI221_X1 U7998 ( .B1(n14332), .B2(n4593), .C1(n5843), .C2(n2209), .A(n3477), 
        .ZN(n3474) );
  AOI21_X1 U7999 ( .B1(n3509), .B2(n3510), .A(n5955), .ZN(n3499) );
  AOI221_X1 U8000 ( .B1(n14431), .B2(n4594), .C1(n14474), .C2(n2210), .A(n3516), .ZN(n3509) );
  AOI221_X1 U8001 ( .B1(n14332), .B2(n4598), .C1(n5799), .C2(n2214), .A(n3513), 
        .ZN(n3510) );
  AOI21_X1 U8002 ( .B1(n3545), .B2(n3546), .A(n5929), .ZN(n3535) );
  AOI221_X1 U8003 ( .B1(n14430), .B2(n4599), .C1(n14473), .C2(n2215), .A(n3552), .ZN(n3545) );
  AOI221_X1 U8004 ( .B1(n14331), .B2(n4601), .C1(n5799), .C2(n2217), .A(n3549), 
        .ZN(n3546) );
  AOI21_X1 U8005 ( .B1(n3622), .B2(n3623), .A(n14289), .ZN(n3612) );
  AOI221_X1 U8006 ( .B1(n14430), .B2(n4602), .C1(n14473), .C2(n2218), .A(n3629), .ZN(n3622) );
  AOI221_X1 U8007 ( .B1(n14331), .B2(n4606), .C1(n5852), .C2(n2222), .A(n3626), 
        .ZN(n3623) );
  AOI21_X1 U8008 ( .B1(n3658), .B2(n3659), .A(n5955), .ZN(n3648) );
  AOI221_X1 U8009 ( .B1(n14429), .B2(n4607), .C1(n14472), .C2(n2223), .A(n3665), .ZN(n3658) );
  AOI221_X1 U8010 ( .B1(n14330), .B2(n4609), .C1(n5860), .C2(n2225), .A(n3662), 
        .ZN(n3659) );
  AOI21_X1 U8011 ( .B1(n3694), .B2(n3695), .A(n5929), .ZN(n3684) );
  AOI221_X1 U8012 ( .B1(n14429), .B2(n4610), .C1(n14472), .C2(n2226), .A(n3701), .ZN(n3694) );
  AOI221_X1 U8013 ( .B1(n14330), .B2(n4623), .C1(n5854), .C2(n2239), .A(n3698), 
        .ZN(n3695) );
  AOI21_X1 U8014 ( .B1(n3771), .B2(n3772), .A(n14289), .ZN(n3761) );
  AOI221_X1 U8015 ( .B1(n14429), .B2(n4624), .C1(n14472), .C2(n2240), .A(n3778), .ZN(n3771) );
  AOI221_X1 U8016 ( .B1(n14330), .B2(n4626), .C1(n5852), .C2(n2242), .A(n3775), 
        .ZN(n3772) );
  AOI21_X1 U8017 ( .B1(n3807), .B2(n3808), .A(n5955), .ZN(n3797) );
  AOI221_X1 U8018 ( .B1(n14428), .B2(n4627), .C1(n14471), .C2(n2243), .A(n3814), .ZN(n3807) );
  AOI221_X1 U8019 ( .B1(n14329), .B2(n4631), .C1(n5855), .C2(n2247), .A(n3811), 
        .ZN(n3808) );
  AOI21_X1 U8020 ( .B1(n3843), .B2(n3844), .A(n5929), .ZN(n3833) );
  AOI221_X1 U8021 ( .B1(n14428), .B2(n4632), .C1(n14471), .C2(n2248), .A(n3850), .ZN(n3843) );
  AOI221_X1 U8022 ( .B1(n14329), .B2(n4634), .C1(n5855), .C2(n2250), .A(n3847), 
        .ZN(n3844) );
  AOI21_X1 U8023 ( .B1(n3920), .B2(n3921), .A(n14289), .ZN(n3910) );
  AOI221_X1 U8024 ( .B1(n14427), .B2(n4635), .C1(n14470), .C2(n2251), .A(n3927), .ZN(n3920) );
  AOI221_X1 U8025 ( .B1(n14328), .B2(n4639), .C1(n5859), .C2(n2255), .A(n3924), 
        .ZN(n3921) );
  AOI21_X1 U8026 ( .B1(n3956), .B2(n3957), .A(n5955), .ZN(n3946) );
  AOI221_X1 U8027 ( .B1(n14427), .B2(n4640), .C1(n14470), .C2(n2256), .A(n3963), .ZN(n3956) );
  AOI221_X1 U8028 ( .B1(n14328), .B2(n4642), .C1(n5859), .C2(n2258), .A(n3960), 
        .ZN(n3957) );
  AOI21_X1 U8029 ( .B1(n3992), .B2(n3993), .A(n5929), .ZN(n3982) );
  AOI221_X1 U8030 ( .B1(n14427), .B2(n4643), .C1(n14470), .C2(n2259), .A(n3999), .ZN(n3992) );
  AOI221_X1 U8031 ( .B1(n14328), .B2(n4647), .C1(n5855), .C2(n2263), .A(n3996), 
        .ZN(n3993) );
  AOI21_X1 U8032 ( .B1(n4069), .B2(n4070), .A(n14289), .ZN(n4059) );
  AOI221_X1 U8033 ( .B1(n14426), .B2(n4648), .C1(n14469), .C2(n2264), .A(n4076), .ZN(n4069) );
  AOI221_X1 U8034 ( .B1(n14327), .B2(n4650), .C1(n5860), .C2(n2266), .A(n4073), 
        .ZN(n4070) );
  AOI21_X1 U8035 ( .B1(n4105), .B2(n4106), .A(n5955), .ZN(n4095) );
  AOI221_X1 U8036 ( .B1(n14426), .B2(n4651), .C1(n14469), .C2(n2267), .A(n4112), .ZN(n4105) );
  AOI221_X1 U8037 ( .B1(n14327), .B2(n4659), .C1(n5860), .C2(n2275), .A(n4109), 
        .ZN(n4106) );
  AOI21_X1 U8038 ( .B1(n4141), .B2(n4142), .A(n5929), .ZN(n4131) );
  AOI221_X1 U8039 ( .B1(n14425), .B2(n4660), .C1(n14468), .C2(n2276), .A(n4148), .ZN(n4141) );
  AOI221_X1 U8040 ( .B1(n14326), .B2(n4662), .C1(n5859), .C2(n2278), .A(n4145), 
        .ZN(n4142) );
  AOI21_X1 U8041 ( .B1(n4218), .B2(n4219), .A(n14289), .ZN(n4208) );
  AOI221_X1 U8042 ( .B1(n14425), .B2(n4663), .C1(n14468), .C2(n2279), .A(n4225), .ZN(n4218) );
  AOI221_X1 U8043 ( .B1(n14326), .B2(n4667), .C1(n5862), .C2(n2283), .A(n4222), 
        .ZN(n4219) );
  AOI21_X1 U8044 ( .B1(n4254), .B2(n4255), .A(n5955), .ZN(n4244) );
  AOI221_X1 U8045 ( .B1(n14425), .B2(n4668), .C1(n14468), .C2(n2284), .A(n4261), .ZN(n4254) );
  AOI221_X1 U8046 ( .B1(n14326), .B2(n4670), .C1(n5860), .C2(n2286), .A(n4258), 
        .ZN(n4255) );
  AOI21_X1 U8047 ( .B1(n4290), .B2(n4291), .A(n5929), .ZN(n4280) );
  AOI221_X1 U8048 ( .B1(n14424), .B2(n4671), .C1(n14467), .C2(n2287), .A(n4297), .ZN(n4290) );
  AOI221_X1 U8049 ( .B1(n14325), .B2(n4675), .C1(n5863), .C2(n2291), .A(n4294), 
        .ZN(n4291) );
  AOI21_X1 U8050 ( .B1(n4367), .B2(n4368), .A(n14289), .ZN(n4357) );
  AOI221_X1 U8051 ( .B1(n14424), .B2(n4676), .C1(n14467), .C2(n2292), .A(n4374), .ZN(n4367) );
  AOI221_X1 U8052 ( .B1(n14325), .B2(n4678), .C1(n5862), .C2(n2294), .A(n4371), 
        .ZN(n4368) );
  AOI21_X1 U8053 ( .B1(n4403), .B2(n4404), .A(n5955), .ZN(n4393) );
  AOI221_X1 U8054 ( .B1(n14423), .B2(n4679), .C1(n14466), .C2(n2295), .A(n4410), .ZN(n4403) );
  AOI221_X1 U8055 ( .B1(n14324), .B2(n4683), .C1(n5867), .C2(n2299), .A(n4407), 
        .ZN(n4404) );
  AOI21_X1 U8056 ( .B1(n4439), .B2(n4440), .A(n5929), .ZN(n4429) );
  AOI221_X1 U8057 ( .B1(n14423), .B2(n4684), .C1(n14466), .C2(n2300), .A(n4446), .ZN(n4439) );
  AOI221_X1 U8058 ( .B1(n14324), .B2(n4686), .C1(n5867), .C2(n2302), .A(n4443), 
        .ZN(n4440) );
  AOI21_X1 U8059 ( .B1(n4516), .B2(n4517), .A(n14289), .ZN(n4506) );
  AOI221_X1 U8060 ( .B1(n14422), .B2(n4687), .C1(n14465), .C2(n2303), .A(n4523), .ZN(n4516) );
  AOI221_X1 U8061 ( .B1(n14323), .B2(n4695), .C1(n5868), .C2(n2311), .A(n4520), 
        .ZN(n4517) );
  AOI21_X1 U8062 ( .B1(n4552), .B2(n4553), .A(n5955), .ZN(n4542) );
  AOI221_X1 U8063 ( .B1(n14422), .B2(n4696), .C1(n14465), .C2(n2312), .A(n4559), .ZN(n4552) );
  AOI221_X1 U8064 ( .B1(n14323), .B2(n4698), .C1(n5868), .C2(n2314), .A(n4556), 
        .ZN(n4553) );
  AOI21_X1 U8065 ( .B1(n4588), .B2(n4589), .A(n5929), .ZN(n4578) );
  AOI221_X1 U8066 ( .B1(n14422), .B2(n4699), .C1(n14465), .C2(n2315), .A(n4595), .ZN(n4588) );
  AOI221_X1 U8067 ( .B1(n14323), .B2(n4703), .C1(n5868), .C2(n2319), .A(n4592), 
        .ZN(n4589) );
  AOI21_X1 U8068 ( .B1(n4665), .B2(n4666), .A(n14289), .ZN(n4655) );
  AOI221_X1 U8069 ( .B1(n14421), .B2(n4704), .C1(n14464), .C2(n2320), .A(n4672), .ZN(n4665) );
  AOI221_X1 U8070 ( .B1(n14322), .B2(n4706), .C1(n5870), .C2(n2322), .A(n4669), 
        .ZN(n4666) );
  AOI21_X1 U8071 ( .B1(n4701), .B2(n4702), .A(n5955), .ZN(n4691) );
  AOI221_X1 U8073 ( .B1(n14421), .B2(n4707), .C1(n14464), .C2(n2323), .A(n4708), .ZN(n4701) );
  AOI221_X1 U8074 ( .B1(n14322), .B2(n4711), .C1(n5870), .C2(n2327), .A(n4705), 
        .ZN(n4702) );
  AOI21_X1 U8075 ( .B1(n4737), .B2(n4738), .A(n5929), .ZN(n4727) );
  AOI221_X1 U8076 ( .B1(n14421), .B2(n4712), .C1(n14464), .C2(n2328), .A(n4744), .ZN(n4737) );
  AOI221_X1 U8077 ( .B1(n14322), .B2(n4714), .C1(n5868), .C2(n2330), .A(n4741), 
        .ZN(n4738) );
  AOI21_X1 U8078 ( .B1(n4814), .B2(n4815), .A(n14289), .ZN(n4804) );
  AOI221_X1 U8079 ( .B1(n14420), .B2(n4715), .C1(n14463), .C2(n2331), .A(n4821), .ZN(n4814) );
  AOI221_X1 U8080 ( .B1(n14321), .B2(n4719), .C1(n5826), .C2(n2335), .A(n4818), 
        .ZN(n4815) );
  AOI21_X1 U8081 ( .B1(n4850), .B2(n4851), .A(n5955), .ZN(n4840) );
  AOI221_X1 U8082 ( .B1(n14420), .B2(n4720), .C1(n14463), .C2(n2336), .A(n4857), .ZN(n4850) );
  AOI221_X1 U8083 ( .B1(n14321), .B2(n4722), .C1(n5875), .C2(n2338), .A(n4854), 
        .ZN(n4851) );
  AOI21_X1 U8084 ( .B1(n4886), .B2(n4887), .A(n5929), .ZN(n4876) );
  AOI221_X1 U8085 ( .B1(n14419), .B2(n4723), .C1(n14462), .C2(n2339), .A(n4893), .ZN(n4886) );
  AOI221_X1 U8086 ( .B1(n14320), .B2(n4731), .C1(n5871), .C2(n2347), .A(n4890), 
        .ZN(n4887) );
  AOI21_X1 U8087 ( .B1(n4963), .B2(n4964), .A(n14289), .ZN(n4953) );
  AOI221_X1 U8088 ( .B1(n14419), .B2(n4732), .C1(n14462), .C2(n2348), .A(n4970), .ZN(n4963) );
  AOI221_X1 U8089 ( .B1(n14320), .B2(n4734), .C1(n5876), .C2(n2350), .A(n4967), 
        .ZN(n4964) );
  AOI21_X1 U8090 ( .B1(n4999), .B2(n5000), .A(n5955), .ZN(n4989) );
  AOI221_X1 U8091 ( .B1(n14418), .B2(n4735), .C1(n14461), .C2(n2351), .A(n5006), .ZN(n4999) );
  AOI221_X1 U8092 ( .B1(n14319), .B2(n4739), .C1(n5875), .C2(n2355), .A(n5003), 
        .ZN(n5000) );
  AOI21_X1 U8093 ( .B1(n5035), .B2(n5036), .A(n5929), .ZN(n5025) );
  AOI221_X1 U8094 ( .B1(n14418), .B2(n4740), .C1(n14461), .C2(n2356), .A(n5042), .ZN(n5035) );
  AOI221_X1 U8095 ( .B1(n14319), .B2(n4742), .C1(n5875), .C2(n2358), .A(n5039), 
        .ZN(n5036) );
  AOI21_X1 U8096 ( .B1(n5112), .B2(n5113), .A(n14290), .ZN(n5102) );
  AOI221_X1 U8097 ( .B1(n14417), .B2(n4743), .C1(n14460), .C2(n2359), .A(n5119), .ZN(n5112) );
  AOI221_X1 U8098 ( .B1(n14318), .B2(n4747), .C1(n5876), .C2(n2363), .A(n5116), 
        .ZN(n5113) );
  AOI21_X1 U8099 ( .B1(n5148), .B2(n5149), .A(n5956), .ZN(n5138) );
  AOI221_X1 U8100 ( .B1(n14417), .B2(n4748), .C1(n14460), .C2(n2364), .A(n5155), .ZN(n5148) );
  AOI221_X1 U8101 ( .B1(n14318), .B2(n4750), .C1(n5876), .C2(n2366), .A(n5152), 
        .ZN(n5149) );
  AOI21_X1 U8102 ( .B1(n5184), .B2(n5185), .A(n5933), .ZN(n5174) );
  AOI221_X1 U8103 ( .B1(n14417), .B2(n4751), .C1(n14460), .C2(n2367), .A(n5191), .ZN(n5184) );
  AOI221_X1 U8104 ( .B1(n14318), .B2(n4755), .C1(n5876), .C2(n2371), .A(n5188), 
        .ZN(n5185) );
  AOI21_X1 U8105 ( .B1(n5261), .B2(n5262), .A(n14290), .ZN(n5251) );
  AOI221_X1 U8106 ( .B1(n14416), .B2(n4756), .C1(n14459), .C2(n2372), .A(n5268), .ZN(n5261) );
  AOI221_X1 U8107 ( .B1(n14317), .B2(n4758), .C1(n5878), .C2(n2374), .A(n5265), 
        .ZN(n5262) );
  AOI21_X1 U8108 ( .B1(n5297), .B2(n5298), .A(n5956), .ZN(n5287) );
  AOI221_X1 U8109 ( .B1(n14416), .B2(n4759), .C1(n14459), .C2(n2375), .A(n5304), .ZN(n5297) );
  AOI221_X1 U8110 ( .B1(n14317), .B2(n4772), .C1(n5878), .C2(n2388), .A(n5301), 
        .ZN(n5298) );
  AOI21_X1 U8111 ( .B1(n5333), .B2(n5334), .A(n5933), .ZN(n5323) );
  AOI221_X1 U8112 ( .B1(n14416), .B2(n4773), .C1(n14459), .C2(n2389), .A(n5340), .ZN(n5333) );
  AOI221_X1 U8113 ( .B1(n14317), .B2(n4775), .C1(n5889), .C2(n2391), .A(n5337), 
        .ZN(n5334) );
  AOI21_X1 U8114 ( .B1(n5410), .B2(n5411), .A(n14290), .ZN(n5400) );
  AOI221_X1 U8115 ( .B1(n14415), .B2(n4776), .C1(n14458), .C2(n2392), .A(n5417), .ZN(n5410) );
  AOI221_X1 U8116 ( .B1(n14316), .B2(n4780), .C1(n5879), .C2(n2396), .A(n5414), 
        .ZN(n5411) );
  AOI21_X1 U8117 ( .B1(n5446), .B2(n5447), .A(n5956), .ZN(n5436) );
  AOI221_X1 U8118 ( .B1(n14415), .B2(n4781), .C1(n14458), .C2(n2397), .A(n5453), .ZN(n5446) );
  AOI221_X1 U8119 ( .B1(n14316), .B2(n4783), .C1(n5890), .C2(n2399), .A(n5450), 
        .ZN(n5447) );
  AOI21_X1 U8120 ( .B1(n5482), .B2(n5483), .A(n5933), .ZN(n5472) );
  AOI221_X1 U8121 ( .B1(n14414), .B2(n4784), .C1(n14457), .C2(n2400), .A(n5489), .ZN(n5482) );
  AOI221_X1 U8122 ( .B1(n14315), .B2(n4788), .C1(n5889), .C2(n2404), .A(n5486), 
        .ZN(n5483) );
  AOI21_X1 U8123 ( .B1(n5559), .B2(n5560), .A(n14290), .ZN(n5549) );
  AOI221_X1 U8124 ( .B1(n14414), .B2(n4789), .C1(n14457), .C2(n2405), .A(n5566), .ZN(n5559) );
  AOI221_X1 U8125 ( .B1(n14315), .B2(n4791), .C1(n5892), .C2(n2407), .A(n5563), 
        .ZN(n5560) );
  AOI21_X1 U8126 ( .B1(n5595), .B2(n5596), .A(n5956), .ZN(n5585) );
  AOI221_X1 U8127 ( .B1(n14413), .B2(n4792), .C1(n14456), .C2(n2408), .A(n5602), .ZN(n5595) );
  AOI221_X1 U8128 ( .B1(n14314), .B2(n4796), .C1(n5890), .C2(n2412), .A(n5599), 
        .ZN(n5596) );
  AOI21_X1 U8129 ( .B1(n5631), .B2(n5632), .A(n5933), .ZN(n5621) );
  AOI221_X1 U8130 ( .B1(n14413), .B2(n4797), .C1(n14456), .C2(n2413), .A(n5638), .ZN(n5631) );
  AOI221_X1 U8131 ( .B1(n14314), .B2(n4799), .C1(n5890), .C2(n2415), .A(n5635), 
        .ZN(n5632) );
  AOI21_X1 U8132 ( .B1(n5708), .B2(n5709), .A(n14290), .ZN(n5698) );
  AOI221_X1 U8133 ( .B1(n14413), .B2(n4800), .C1(n14456), .C2(n2416), .A(n5715), .ZN(n5708) );
  AOI221_X1 U8134 ( .B1(n14314), .B2(n4808), .C1(n5893), .C2(n2424), .A(n5712), 
        .ZN(n5709) );
  AOI21_X1 U8135 ( .B1(n5744), .B2(n5745), .A(n5956), .ZN(n5734) );
  AOI221_X1 U8136 ( .B1(n14412), .B2(n4809), .C1(n14455), .C2(n2425), .A(n5751), .ZN(n5744) );
  AOI221_X1 U8137 ( .B1(n14313), .B2(n4811), .C1(n5892), .C2(n2427), .A(n5748), 
        .ZN(n5745) );
  AOI21_X1 U8138 ( .B1(n5780), .B2(n5781), .A(n5933), .ZN(n5770) );
  AOI221_X1 U8139 ( .B1(n14412), .B2(n4812), .C1(n14455), .C2(n2428), .A(n5787), .ZN(n5780) );
  AOI221_X1 U8140 ( .B1(n14313), .B2(n4816), .C1(n5892), .C2(n2432), .A(n5784), 
        .ZN(n5781) );
  AOI21_X1 U8141 ( .B1(n5857), .B2(n5858), .A(n14290), .ZN(n5847) );
  AOI221_X1 U8142 ( .B1(n14411), .B2(n4817), .C1(n14454), .C2(n2433), .A(n5864), .ZN(n5857) );
  AOI221_X1 U8143 ( .B1(n14312), .B2(n4819), .C1(n5893), .C2(n2435), .A(n5861), 
        .ZN(n5858) );
  AOI21_X1 U8144 ( .B1(n5895), .B2(n5896), .A(n5956), .ZN(n5883) );
  AOI221_X1 U8145 ( .B1(n14411), .B2(n4820), .C1(n14454), .C2(n2436), .A(n5902), .ZN(n5895) );
  AOI221_X1 U8146 ( .B1(n14312), .B2(n4824), .C1(n5893), .C2(n2440), .A(n5899), 
        .ZN(n5896) );
  AOI21_X1 U8147 ( .B1(n5931), .B2(n5932), .A(n5933), .ZN(n5921) );
  AOI221_X1 U8148 ( .B1(n14411), .B2(n4825), .C1(n14454), .C2(n2441), .A(n5938), .ZN(n5931) );
  AOI221_X1 U8149 ( .B1(n14312), .B2(n4827), .C1(n5889), .C2(n2443), .A(n5935), 
        .ZN(n5932) );
  AOI21_X1 U8150 ( .B1(n1236), .B2(n1237), .A(n14285), .ZN(n1215) );
  AOI221_X1 U8151 ( .B1(n14449), .B2(n4828), .C1(n14492), .C2(n2444), .A(n1244), .ZN(n1236) );
  AOI221_X1 U8152 ( .B1(n14350), .B2(n4832), .C1(n5851), .C2(n2448), .A(n1241), 
        .ZN(n1237) );
  AOI21_X1 U8153 ( .B1(n1276), .B2(n1277), .A(n5945), .ZN(n1255) );
  AOI221_X1 U8154 ( .B1(n14449), .B2(n4833), .C1(n14492), .C2(n2449), .A(n1284), .ZN(n1276) );
  AOI221_X1 U8155 ( .B1(n14350), .B2(n4835), .C1(n5801), .C2(n2451), .A(n1281), 
        .ZN(n1277) );
  AOI21_X1 U8156 ( .B1(n1316), .B2(n1317), .A(n5917), .ZN(n1295) );
  AOI221_X1 U8157 ( .B1(n14449), .B2(n4836), .C1(n14492), .C2(n2452), .A(n1324), .ZN(n1316) );
  AOI221_X1 U8158 ( .B1(n14350), .B2(n4844), .C1(n5799), .C2(n2460), .A(n1321), 
        .ZN(n1317) );
  AOI21_X1 U8159 ( .B1(n1395), .B2(n1396), .A(n14285), .ZN(n1376) );
  AOI221_X1 U8160 ( .B1(n14448), .B2(n4845), .C1(n14491), .C2(n2461), .A(n1402), .ZN(n1395) );
  AOI221_X1 U8161 ( .B1(n14349), .B2(n4847), .C1(n5802), .C2(n2463), .A(n1399), 
        .ZN(n1396) );
  AOI21_X1 U8162 ( .B1(n1431), .B2(n1432), .A(n5945), .ZN(n1412) );
  AOI221_X1 U8163 ( .B1(n14448), .B2(n4848), .C1(n14491), .C2(n2464), .A(n1438), .ZN(n1431) );
  AOI221_X1 U8164 ( .B1(n14349), .B2(n4852), .C1(n5802), .C2(n2468), .A(n1435), 
        .ZN(n1432) );
  AOI21_X1 U8165 ( .B1(n1467), .B2(n1468), .A(n5917), .ZN(n1448) );
  AOI221_X1 U8166 ( .B1(n14448), .B2(n4853), .C1(n14491), .C2(n2469), .A(n1474), .ZN(n1467) );
  AOI221_X1 U8167 ( .B1(n14349), .B2(n4855), .C1(n5801), .C2(n2471), .A(n1471), 
        .ZN(n1468) );
  AOI21_X1 U8168 ( .B1(n1544), .B2(n1545), .A(n14285), .ZN(n1525) );
  AOI221_X1 U8169 ( .B1(n14447), .B2(n4856), .C1(n14490), .C2(n2472), .A(n1551), .ZN(n1544) );
  AOI221_X1 U8170 ( .B1(n14348), .B2(n4860), .C1(n5815), .C2(n2476), .A(n1548), 
        .ZN(n1545) );
  AOI21_X1 U8171 ( .B1(n1580), .B2(n1581), .A(n5945), .ZN(n1561) );
  AOI221_X1 U8172 ( .B1(n14447), .B2(n4861), .C1(n14490), .C2(n2477), .A(n1587), .ZN(n1580) );
  AOI221_X1 U8173 ( .B1(n14348), .B2(n4863), .C1(n5802), .C2(n2479), .A(n1584), 
        .ZN(n1581) );
  AOI21_X1 U8174 ( .B1(n1616), .B2(n1617), .A(n5917), .ZN(n1597) );
  AOI221_X1 U8175 ( .B1(n14446), .B2(n4864), .C1(n14489), .C2(n2480), .A(n1623), .ZN(n1616) );
  AOI221_X1 U8176 ( .B1(n14347), .B2(n4868), .C1(n5816), .C2(n2484), .A(n1620), 
        .ZN(n1617) );
  AOI21_X1 U8177 ( .B1(n1693), .B2(n1694), .A(n14285), .ZN(n1674) );
  AOI221_X1 U8178 ( .B1(n14446), .B2(n4869), .C1(n14489), .C2(n2485), .A(n1700), .ZN(n1693) );
  AOI221_X1 U8179 ( .B1(n14347), .B2(n4871), .C1(n5815), .C2(n2487), .A(n1697), 
        .ZN(n1694) );
  AOI21_X1 U8180 ( .B1(n1729), .B2(n1730), .A(n5945), .ZN(n1710) );
  AOI221_X1 U8181 ( .B1(n14445), .B2(n4872), .C1(n14488), .C2(n2488), .A(n1736), .ZN(n1729) );
  AOI221_X1 U8182 ( .B1(n14346), .B2(n4880), .C1(n5815), .C2(n2496), .A(n1733), 
        .ZN(n1730) );
  AOI21_X1 U8183 ( .B1(n1765), .B2(n1766), .A(n5917), .ZN(n1746) );
  AOI221_X1 U8184 ( .B1(n14445), .B2(n4881), .C1(n14488), .C2(n2497), .A(n1772), .ZN(n1765) );
  AOI221_X1 U8185 ( .B1(n14346), .B2(n4883), .C1(n5799), .C2(n2499), .A(n1769), 
        .ZN(n1766) );
  AOI21_X1 U8186 ( .B1(n1842), .B2(n1843), .A(n14285), .ZN(n1823) );
  AOI221_X1 U8187 ( .B1(n14444), .B2(n4884), .C1(n14487), .C2(n2500), .A(n1849), .ZN(n1842) );
  AOI221_X1 U8188 ( .B1(n14345), .B2(n4888), .C1(n5816), .C2(n2504), .A(n1846), 
        .ZN(n1843) );
  AOI21_X1 U8189 ( .B1(n1878), .B2(n1879), .A(n5945), .ZN(n1859) );
  AOI221_X1 U8190 ( .B1(n14444), .B2(n4889), .C1(n14487), .C2(n2505), .A(n1885), .ZN(n1878) );
  AOI221_X1 U8191 ( .B1(n14345), .B2(n4891), .C1(n5819), .C2(n2507), .A(n1882), 
        .ZN(n1879) );
  AOI21_X1 U8192 ( .B1(n1914), .B2(n1915), .A(n5917), .ZN(n1895) );
  AOI221_X1 U8193 ( .B1(n14444), .B2(n4892), .C1(n14487), .C2(n2508), .A(n1921), .ZN(n1914) );
  AOI221_X1 U8194 ( .B1(n14345), .B2(n4896), .C1(n5819), .C2(n2512), .A(n1918), 
        .ZN(n1915) );
  AOI21_X1 U8195 ( .B1(n1991), .B2(n1992), .A(n14285), .ZN(n1972) );
  AOI221_X1 U8196 ( .B1(n14443), .B2(n4897), .C1(n14486), .C2(n2513), .A(n1998), .ZN(n1991) );
  AOI221_X1 U8197 ( .B1(n14344), .B2(n4899), .C1(n5823), .C2(n2515), .A(n1995), 
        .ZN(n1992) );
  AOI21_X1 U8198 ( .B1(n2027), .B2(n2028), .A(n5945), .ZN(n2008) );
  AOI221_X1 U8199 ( .B1(n14443), .B2(n4900), .C1(n14486), .C2(n2516), .A(n2034), .ZN(n2027) );
  AOI221_X1 U8200 ( .B1(n14344), .B2(n4904), .C1(n5823), .C2(n2520), .A(n2031), 
        .ZN(n2028) );
  AOI21_X1 U8201 ( .B1(n2063), .B2(n2064), .A(n5917), .ZN(n2044) );
  AOI221_X1 U8202 ( .B1(n14443), .B2(n4905), .C1(n14486), .C2(n2521), .A(n2070), .ZN(n2063) );
  AOI221_X1 U8203 ( .B1(n14344), .B2(n4907), .C1(n5819), .C2(n2523), .A(n2067), 
        .ZN(n2064) );
  AOI21_X1 U8204 ( .B1(n2140), .B2(n2141), .A(n14285), .ZN(n2121) );
  AOI221_X1 U8205 ( .B1(n14442), .B2(n4908), .C1(n14485), .C2(n2524), .A(n2147), .ZN(n2140) );
  AOI221_X1 U8206 ( .B1(n14343), .B2(n4921), .C1(n5824), .C2(n2537), .A(n2144), 
        .ZN(n2141) );
  AOI21_X1 U8207 ( .B1(n2176), .B2(n2177), .A(n5945), .ZN(n2157) );
  AOI221_X1 U8208 ( .B1(n14442), .B2(n4922), .C1(n14485), .C2(n2538), .A(n2183), .ZN(n2176) );
  AOI221_X1 U8209 ( .B1(n14343), .B2(n4924), .C1(n5823), .C2(n2540), .A(n2180), 
        .ZN(n2177) );
  AOI21_X1 U8210 ( .B1(n2212), .B2(n2213), .A(n5917), .ZN(n2193) );
  AOI221_X1 U8211 ( .B1(n14441), .B2(n4925), .C1(n14484), .C2(n2541), .A(n2219), .ZN(n2212) );
  AOI221_X1 U8212 ( .B1(n14342), .B2(n4929), .C1(n5823), .C2(n2545), .A(n2216), 
        .ZN(n2213) );
  AOI21_X1 U8213 ( .B1(n2289), .B2(n2290), .A(n14285), .ZN(n2270) );
  AOI221_X1 U8214 ( .B1(n14441), .B2(n4930), .C1(n14484), .C2(n2546), .A(n2296), .ZN(n2289) );
  AOI221_X1 U8215 ( .B1(n14342), .B2(n4932), .C1(n5826), .C2(n2548), .A(n2293), 
        .ZN(n2290) );
  AOI21_X1 U8216 ( .B1(n2325), .B2(n2326), .A(n5945), .ZN(n2306) );
  AOI221_X1 U8217 ( .B1(n14440), .B2(n4933), .C1(n14483), .C2(n2549), .A(n2332), .ZN(n2325) );
  AOI221_X1 U8218 ( .B1(n14341), .B2(n4937), .C1(n5824), .C2(n2553), .A(n2329), 
        .ZN(n2326) );
  AOI21_X1 U8219 ( .B1(n2361), .B2(n2362), .A(n5917), .ZN(n2342) );
  AOI221_X1 U8220 ( .B1(n14440), .B2(n4938), .C1(n14483), .C2(n2554), .A(n2368), .ZN(n2361) );
  AOI221_X1 U8221 ( .B1(n14341), .B2(n4940), .C1(n5871), .C2(n2556), .A(n2365), 
        .ZN(n2362) );
  AOI21_X1 U8222 ( .B1(n2438), .B2(n2439), .A(n14285), .ZN(n2419) );
  AOI221_X1 U8223 ( .B1(n14440), .B2(n4941), .C1(n14483), .C2(n2557), .A(n2445), .ZN(n2438) );
  AOI221_X1 U8225 ( .B1(n14341), .B2(n4945), .C1(n5831), .C2(n2561), .A(n2442), 
        .ZN(n2439) );
  AOI21_X1 U8226 ( .B1(n2474), .B2(n2475), .A(n5945), .ZN(n2455) );
  AOI221_X1 U8227 ( .B1(n14439), .B2(n4946), .C1(n14482), .C2(n2562), .A(n2481), .ZN(n2474) );
  AOI221_X1 U8228 ( .B1(n14340), .B2(n4948), .C1(n5827), .C2(n2564), .A(n2478), 
        .ZN(n2475) );
  AOI21_X1 U8229 ( .B1(n2510), .B2(n2511), .A(n5917), .ZN(n2491) );
  AOI221_X1 U8230 ( .B1(n14439), .B2(n4949), .C1(n14482), .C2(n2565), .A(n2517), .ZN(n2510) );
  AOI221_X1 U8231 ( .B1(n14340), .B2(n4957), .C1(n5827), .C2(n2573), .A(n2514), 
        .ZN(n2511) );
  AOI21_X1 U8232 ( .B1(n2587), .B2(n2588), .A(n14285), .ZN(n2568) );
  AOI221_X1 U8233 ( .B1(n14438), .B2(n4958), .C1(n14481), .C2(n2574), .A(n2594), .ZN(n2587) );
  AOI221_X1 U8234 ( .B1(n14339), .B2(n4960), .C1(n5831), .C2(n2576), .A(n2591), 
        .ZN(n2588) );
  AOI21_X1 U8235 ( .B1(n2623), .B2(n2624), .A(n5945), .ZN(n2604) );
  AOI221_X1 U8236 ( .B1(n14438), .B2(n4961), .C1(n14481), .C2(n2577), .A(n2630), .ZN(n2623) );
  AOI221_X1 U8237 ( .B1(n14339), .B2(n4965), .C1(n5831), .C2(n2581), .A(n2627), 
        .ZN(n2624) );
  AOI21_X1 U8238 ( .B1(n2659), .B2(n2660), .A(n5917), .ZN(n2640) );
  AOI221_X1 U8239 ( .B1(n14438), .B2(n4966), .C1(n14481), .C2(n2582), .A(n2666), .ZN(n2659) );
  AOI221_X1 U8240 ( .B1(n14339), .B2(n4968), .C1(n5831), .C2(n2584), .A(n2663), 
        .ZN(n2660) );
  AOI21_X1 U8241 ( .B1(n2736), .B2(n2737), .A(n14285), .ZN(n2717) );
  AOI221_X1 U8242 ( .B1(n14437), .B2(n4969), .C1(n14480), .C2(n2585), .A(n2743), .ZN(n2736) );
  AOI221_X1 U8243 ( .B1(n14338), .B2(n4973), .C1(n5832), .C2(n2589), .A(n2740), 
        .ZN(n2737) );
  AOI21_X1 U8244 ( .B1(n2772), .B2(n2773), .A(n5945), .ZN(n2753) );
  AOI221_X1 U8245 ( .B1(n14437), .B2(n4974), .C1(n14480), .C2(n2590), .A(n2779), .ZN(n2772) );
  AOI221_X1 U8246 ( .B1(n14338), .B2(n4976), .C1(n5832), .C2(n2592), .A(n2776), 
        .ZN(n2773) );
  AOI21_X1 U8247 ( .B1(n2808), .B2(n2809), .A(n5917), .ZN(n2789) );
  AOI221_X1 U8248 ( .B1(n14436), .B2(n4977), .C1(n14479), .C2(n2593), .A(n2815), .ZN(n2808) );
  AOI221_X1 U8249 ( .B1(n14337), .B2(n4981), .C1(n5835), .C2(n2597), .A(n2812), 
        .ZN(n2809) );
  AOI21_X1 U8250 ( .B1(n2885), .B2(n2886), .A(n14285), .ZN(n2866) );
  AOI221_X1 U8251 ( .B1(n14436), .B2(n4982), .C1(n14479), .C2(n2598), .A(n2892), .ZN(n2885) );
  AOI221_X1 U8252 ( .B1(n14337), .B2(n4984), .C1(n5834), .C2(n2600), .A(n2889), 
        .ZN(n2886) );
  AOI21_X1 U8253 ( .B1(n2921), .B2(n2922), .A(n5945), .ZN(n2902) );
  AOI221_X1 U8254 ( .B1(n14436), .B2(n4985), .C1(n14479), .C2(n2601), .A(n2928), .ZN(n2921) );
  AOI221_X1 U8255 ( .B1(n14337), .B2(n4993), .C1(n5839), .C2(n2609), .A(n2925), 
        .ZN(n2922) );
  AOI21_X1 U8256 ( .B1(n2957), .B2(n2958), .A(n5917), .ZN(n2938) );
  AOI221_X1 U8257 ( .B1(n14435), .B2(n4994), .C1(n14478), .C2(n2610), .A(n2964), .ZN(n2957) );
  AOI221_X1 U8258 ( .B1(n14336), .B2(n4996), .C1(n5835), .C2(n2612), .A(n2961), 
        .ZN(n2958) );
  AOI21_X1 U8259 ( .B1(n3034), .B2(n3035), .A(n14285), .ZN(n3015) );
  AOI221_X1 U8260 ( .B1(n14435), .B2(n4997), .C1(n14478), .C2(n2613), .A(n3041), .ZN(n3034) );
  AOI221_X1 U8261 ( .B1(n14336), .B2(n5001), .C1(n5840), .C2(n2617), .A(n3038), 
        .ZN(n3035) );
  AOI21_X1 U8262 ( .B1(n3070), .B2(n3071), .A(n5945), .ZN(n3051) );
  AOI221_X1 U8263 ( .B1(n14434), .B2(n5002), .C1(n14477), .C2(n2618), .A(n3077), .ZN(n3070) );
  AOI221_X1 U8264 ( .B1(n14335), .B2(n5004), .C1(n5839), .C2(n2620), .A(n3074), 
        .ZN(n3071) );
  AOI21_X1 U8265 ( .B1(n3106), .B2(n3107), .A(n5917), .ZN(n3087) );
  AOI221_X1 U8266 ( .B1(n14434), .B2(n5005), .C1(n14477), .C2(n2621), .A(n3113), .ZN(n3106) );
  AOI221_X1 U8267 ( .B1(n14335), .B2(n5009), .C1(n5839), .C2(n2625), .A(n3110), 
        .ZN(n3107) );
  AOI21_X1 U8268 ( .B1(n3183), .B2(n3184), .A(n14286), .ZN(n3164) );
  AOI221_X1 U8269 ( .B1(n14433), .B2(n5010), .C1(n14476), .C2(n2626), .A(n3190), .ZN(n3183) );
  AOI221_X1 U8270 ( .B1(n14334), .B2(n5012), .C1(n5840), .C2(n2628), .A(n3187), 
        .ZN(n3184) );
  AOI21_X1 U8271 ( .B1(n3219), .B2(n3220), .A(n5949), .ZN(n3200) );
  AOI221_X1 U8272 ( .B1(n14433), .B2(n5013), .C1(n14476), .C2(n2629), .A(n3226), .ZN(n3219) );
  AOI221_X1 U8273 ( .B1(n14334), .B2(n5017), .C1(n5840), .C2(n2633), .A(n3223), 
        .ZN(n3220) );
  AOI21_X1 U8274 ( .B1(n3255), .B2(n3256), .A(n5925), .ZN(n3236) );
  AOI221_X1 U8275 ( .B1(n14433), .B2(n5018), .C1(n14476), .C2(n2634), .A(n3262), .ZN(n3255) );
  AOI221_X1 U8276 ( .B1(n14334), .B2(n5020), .C1(n5840), .C2(n2636), .A(n3259), 
        .ZN(n3256) );
  AOI21_X1 U8277 ( .B1(n3332), .B2(n3333), .A(n14286), .ZN(n3313) );
  AOI221_X1 U8278 ( .B1(n14432), .B2(n5021), .C1(n14475), .C2(n2637), .A(n3339), .ZN(n3332) );
  AOI221_X1 U8279 ( .B1(n14333), .B2(n5029), .C1(n5842), .C2(n2645), .A(n3336), 
        .ZN(n3333) );
  AOI21_X1 U8280 ( .B1(n3368), .B2(n3369), .A(n5949), .ZN(n3349) );
  AOI221_X1 U8281 ( .B1(n14432), .B2(n5030), .C1(n14475), .C2(n2646), .A(n3375), .ZN(n3368) );
  AOI221_X1 U8282 ( .B1(n14333), .B2(n5032), .C1(n5842), .C2(n2648), .A(n3372), 
        .ZN(n3369) );
  AOI21_X1 U8283 ( .B1(n3404), .B2(n3405), .A(n5925), .ZN(n3385) );
  AOI221_X1 U8284 ( .B1(n14432), .B2(n5033), .C1(n14475), .C2(n2649), .A(n3411), .ZN(n3404) );
  AOI221_X1 U8285 ( .B1(n14333), .B2(n5037), .C1(n5851), .C2(n2653), .A(n3408), 
        .ZN(n3405) );
  AOI21_X1 U8286 ( .B1(n3481), .B2(n3482), .A(n14286), .ZN(n3462) );
  AOI221_X1 U8287 ( .B1(n14431), .B2(n5038), .C1(n14474), .C2(n2654), .A(n3488), .ZN(n3481) );
  AOI221_X1 U8288 ( .B1(n14332), .B2(n5040), .C1(n5843), .C2(n2656), .A(n3485), 
        .ZN(n3482) );
  AOI21_X1 U8289 ( .B1(n3517), .B2(n3518), .A(n5949), .ZN(n3498) );
  AOI221_X1 U8290 ( .B1(n14431), .B2(n5041), .C1(n14474), .C2(n2657), .A(n3524), .ZN(n3517) );
  AOI221_X1 U8291 ( .B1(n14332), .B2(n5045), .C1(n5799), .C2(n2661), .A(n3521), 
        .ZN(n3518) );
  AOI21_X1 U8292 ( .B1(n3553), .B2(n3554), .A(n5925), .ZN(n3534) );
  AOI221_X1 U8293 ( .B1(n14430), .B2(n5046), .C1(n14473), .C2(n2662), .A(n3560), .ZN(n3553) );
  AOI221_X1 U8294 ( .B1(n14331), .B2(n5048), .C1(n5835), .C2(n2664), .A(n3557), 
        .ZN(n3554) );
  AOI21_X1 U8295 ( .B1(n3630), .B2(n3631), .A(n14286), .ZN(n3611) );
  AOI221_X1 U8296 ( .B1(n14430), .B2(n5049), .C1(n14473), .C2(n2665), .A(n3637), .ZN(n3630) );
  AOI221_X1 U8297 ( .B1(n14331), .B2(n5053), .C1(n5851), .C2(n2669), .A(n3634), 
        .ZN(n3631) );
  AOI21_X1 U8298 ( .B1(n3702), .B2(n3703), .A(n5925), .ZN(n3683) );
  AOI221_X1 U8299 ( .B1(n14429), .B2(n5054), .C1(n14472), .C2(n2670), .A(n3709), .ZN(n3702) );
  AOI221_X1 U8300 ( .B1(n14330), .B2(n5056), .C1(n5854), .C2(n2672), .A(n3706), 
        .ZN(n3703) );
  AOI21_X1 U8301 ( .B1(n3779), .B2(n3780), .A(n14286), .ZN(n3760) );
  AOI221_X1 U8302 ( .B1(n14428), .B2(n5057), .C1(n14471), .C2(n2673), .A(n3786), .ZN(n3779) );
  AOI221_X1 U8303 ( .B1(n14329), .B2(n5070), .C1(n5852), .C2(n2686), .A(n3783), 
        .ZN(n3780) );
  AOI21_X1 U8304 ( .B1(n3815), .B2(n3816), .A(n5949), .ZN(n3796) );
  AOI221_X1 U8305 ( .B1(n14428), .B2(n5071), .C1(n14471), .C2(n2687), .A(n3822), .ZN(n3815) );
  AOI221_X1 U8306 ( .B1(n14329), .B2(n5073), .C1(n5855), .C2(n2689), .A(n3819), 
        .ZN(n3816) );
  AOI21_X1 U8307 ( .B1(n3851), .B2(n3852), .A(n5925), .ZN(n3832) );
  AOI221_X1 U8308 ( .B1(n14428), .B2(n5074), .C1(n14471), .C2(n2690), .A(n3858), .ZN(n3851) );
  AOI221_X1 U8309 ( .B1(n14329), .B2(n5078), .C1(n5855), .C2(n2694), .A(n3855), 
        .ZN(n3852) );
  AOI21_X1 U8310 ( .B1(n3928), .B2(n3929), .A(n14286), .ZN(n3909) );
  AOI221_X1 U8311 ( .B1(n14427), .B2(n5079), .C1(n14470), .C2(n2695), .A(n3935), .ZN(n3928) );
  AOI221_X1 U8312 ( .B1(n14328), .B2(n5081), .C1(n5859), .C2(n2697), .A(n3932), 
        .ZN(n3929) );
  AOI21_X1 U8313 ( .B1(n3964), .B2(n3965), .A(n5949), .ZN(n3945) );
  AOI221_X1 U8314 ( .B1(n14427), .B2(n5082), .C1(n14470), .C2(n2698), .A(n3971), .ZN(n3964) );
  AOI221_X1 U8315 ( .B1(n14328), .B2(n5086), .C1(n5859), .C2(n2702), .A(n3968), 
        .ZN(n3965) );
  AOI21_X1 U8316 ( .B1(n4000), .B2(n4001), .A(n5925), .ZN(n3981) );
  AOI221_X1 U8317 ( .B1(n14427), .B2(n5087), .C1(n14470), .C2(n2703), .A(n4007), .ZN(n4000) );
  AOI221_X1 U8318 ( .B1(n14328), .B2(n5089), .C1(n5855), .C2(n2705), .A(n4004), 
        .ZN(n4001) );
  AOI21_X1 U8319 ( .B1(n4077), .B2(n4078), .A(n14286), .ZN(n4058) );
  AOI221_X1 U8320 ( .B1(n14426), .B2(n5090), .C1(n14469), .C2(n2706), .A(n4084), .ZN(n4077) );
  AOI221_X1 U8321 ( .B1(n14327), .B2(n5094), .C1(n5860), .C2(n2710), .A(n4081), 
        .ZN(n4078) );
  AOI21_X1 U8322 ( .B1(n4113), .B2(n4114), .A(n5949), .ZN(n4094) );
  AOI221_X1 U8323 ( .B1(n14426), .B2(n5095), .C1(n14469), .C2(n2711), .A(n4120), .ZN(n4113) );
  AOI221_X1 U8324 ( .B1(n14327), .B2(n5097), .C1(n5859), .C2(n2713), .A(n4117), 
        .ZN(n4114) );
  AOI21_X1 U8325 ( .B1(n4149), .B2(n4150), .A(n5925), .ZN(n4130) );
  AOI221_X1 U8326 ( .B1(n14425), .B2(n5098), .C1(n14468), .C2(n2714), .A(n4156), .ZN(n4149) );
  AOI221_X1 U8327 ( .B1(n14326), .B2(n5106), .C1(n5859), .C2(n2722), .A(n4153), 
        .ZN(n4150) );
  AOI21_X1 U8328 ( .B1(n4226), .B2(n4227), .A(n14286), .ZN(n4207) );
  AOI221_X1 U8329 ( .B1(n14425), .B2(n5107), .C1(n14468), .C2(n2723), .A(n4233), .ZN(n4226) );
  AOI221_X1 U8330 ( .B1(n14326), .B2(n5109), .C1(n5862), .C2(n2725), .A(n4230), 
        .ZN(n4227) );
  AOI21_X1 U8331 ( .B1(n4262), .B2(n4263), .A(n5949), .ZN(n4243) );
  AOI221_X1 U8332 ( .B1(n14424), .B2(n5110), .C1(n14467), .C2(n2726), .A(n4269), .ZN(n4262) );
  AOI221_X1 U8333 ( .B1(n14325), .B2(n5114), .C1(n5860), .C2(n2730), .A(n4266), 
        .ZN(n4263) );
  AOI21_X1 U8334 ( .B1(n4298), .B2(n4299), .A(n5925), .ZN(n4279) );
  AOI221_X1 U8335 ( .B1(n14424), .B2(n5115), .C1(n14467), .C2(n2731), .A(n4305), .ZN(n4298) );
  AOI221_X1 U8336 ( .B1(n14325), .B2(n5117), .C1(n5863), .C2(n2733), .A(n4302), 
        .ZN(n4299) );
  AOI21_X1 U8337 ( .B1(n4375), .B2(n4376), .A(n14286), .ZN(n4356) );
  AOI221_X1 U8338 ( .B1(n14424), .B2(n5118), .C1(n14467), .C2(n2734), .A(n4382), .ZN(n4375) );
  AOI221_X1 U8339 ( .B1(n14325), .B2(n5122), .C1(n5862), .C2(n2738), .A(n4379), 
        .ZN(n4376) );
  AOI21_X1 U8340 ( .B1(n4411), .B2(n4412), .A(n5949), .ZN(n4392) );
  AOI221_X1 U8341 ( .B1(n14423), .B2(n5123), .C1(n14466), .C2(n2739), .A(n4418), .ZN(n4411) );
  AOI221_X1 U8342 ( .B1(n14324), .B2(n5125), .C1(n5867), .C2(n2741), .A(n4415), 
        .ZN(n4412) );
  AOI21_X1 U8343 ( .B1(n4447), .B2(n4448), .A(n5925), .ZN(n4428) );
  AOI221_X1 U8344 ( .B1(n14423), .B2(n5126), .C1(n14466), .C2(n2742), .A(n4454), .ZN(n4447) );
  AOI221_X1 U8345 ( .B1(n14324), .B2(n5130), .C1(n5867), .C2(n2746), .A(n4451), 
        .ZN(n4448) );
  AOI21_X1 U8346 ( .B1(n4524), .B2(n4525), .A(n14286), .ZN(n4505) );
  AOI221_X1 U8347 ( .B1(n14422), .B2(n5131), .C1(n14465), .C2(n2747), .A(n4531), .ZN(n4524) );
  AOI221_X1 U8348 ( .B1(n14323), .B2(n5133), .C1(n5868), .C2(n2749), .A(n4528), 
        .ZN(n4525) );
  AOI21_X1 U8349 ( .B1(n4560), .B2(n4561), .A(n5949), .ZN(n4541) );
  AOI221_X1 U8350 ( .B1(n14422), .B2(n5134), .C1(n14465), .C2(n2750), .A(n4567), .ZN(n4560) );
  AOI221_X1 U8351 ( .B1(n14323), .B2(n5142), .C1(n5868), .C2(n2758), .A(n4564), 
        .ZN(n4561) );
  AOI21_X1 U8352 ( .B1(n4596), .B2(n4597), .A(n5925), .ZN(n4577) );
  AOI221_X1 U8353 ( .B1(n14422), .B2(n5143), .C1(n14465), .C2(n2759), .A(n4603), .ZN(n4596) );
  AOI221_X1 U8354 ( .B1(n14323), .B2(n5145), .C1(n5867), .C2(n2761), .A(n4600), 
        .ZN(n4597) );
  AOI21_X1 U8355 ( .B1(n4673), .B2(n4674), .A(n14286), .ZN(n4654) );
  AOI221_X1 U8356 ( .B1(n14421), .B2(n5146), .C1(n14464), .C2(n2762), .A(n4680), .ZN(n4673) );
  AOI221_X1 U8357 ( .B1(n14322), .B2(n5150), .C1(n5870), .C2(n2766), .A(n4677), 
        .ZN(n4674) );
  AOI21_X1 U8358 ( .B1(n4709), .B2(n4710), .A(n5949), .ZN(n4690) );
  AOI221_X1 U8359 ( .B1(n14421), .B2(n5151), .C1(n14464), .C2(n2767), .A(n4716), .ZN(n4709) );
  AOI221_X1 U8360 ( .B1(n14322), .B2(n5153), .C1(n5870), .C2(n2769), .A(n4713), 
        .ZN(n4710) );
  AOI21_X1 U8361 ( .B1(n4745), .B2(n4746), .A(n5925), .ZN(n4726) );
  AOI221_X1 U8362 ( .B1(n14420), .B2(n5154), .C1(n14463), .C2(n2770), .A(n4752), .ZN(n4745) );
  AOI221_X1 U8363 ( .B1(n14321), .B2(n5158), .C1(n5862), .C2(n2774), .A(n4749), 
        .ZN(n4746) );
  AOI21_X1 U8364 ( .B1(n4822), .B2(n4823), .A(n14286), .ZN(n4803) );
  AOI221_X1 U8365 ( .B1(n14420), .B2(n5159), .C1(n14463), .C2(n2775), .A(n4829), .ZN(n4822) );
  AOI221_X1 U8366 ( .B1(n14321), .B2(n5161), .C1(n5826), .C2(n2777), .A(n4826), 
        .ZN(n4823) );
  AOI21_X1 U8367 ( .B1(n4858), .B2(n4859), .A(n5949), .ZN(n4839) );
  AOI221_X1 U8368 ( .B1(n14420), .B2(n5162), .C1(n14463), .C2(n2778), .A(n4865), .ZN(n4858) );
  AOI221_X1 U8369 ( .B1(n14321), .B2(n5166), .C1(n5875), .C2(n2782), .A(n4862), 
        .ZN(n4859) );
  AOI21_X1 U8370 ( .B1(n4894), .B2(n4895), .A(n5925), .ZN(n4875) );
  AOI221_X1 U8371 ( .B1(n14419), .B2(n5167), .C1(n14462), .C2(n2783), .A(n4901), .ZN(n4894) );
  AOI221_X1 U8372 ( .B1(n14320), .B2(n5169), .C1(n5871), .C2(n2785), .A(n4898), 
        .ZN(n4895) );
  AOI21_X1 U8373 ( .B1(n4971), .B2(n4972), .A(n14286), .ZN(n4952) );
  AOI221_X1 U8374 ( .B1(n14419), .B2(n5170), .C1(n14462), .C2(n2786), .A(n4978), .ZN(n4971) );
  AOI221_X1 U8375 ( .B1(n14320), .B2(n5178), .C1(n5876), .C2(n2794), .A(n4975), 
        .ZN(n4972) );
  AOI21_X1 U8377 ( .B1(n5007), .B2(n5008), .A(n5949), .ZN(n4988) );
  AOI221_X1 U8378 ( .B1(n14418), .B2(n5179), .C1(n14461), .C2(n2795), .A(n5014), .ZN(n5007) );
  AOI221_X1 U8379 ( .B1(n14319), .B2(n5181), .C1(n5875), .C2(n2797), .A(n5011), 
        .ZN(n5008) );
  AOI21_X1 U8380 ( .B1(n5043), .B2(n5044), .A(n5925), .ZN(n5024) );
  AOI221_X1 U8381 ( .B1(n14418), .B2(n5182), .C1(n14461), .C2(n2798), .A(n5050), .ZN(n5043) );
  AOI221_X1 U8382 ( .B1(n14319), .B2(n5186), .C1(n5875), .C2(n2802), .A(n5047), 
        .ZN(n5044) );
  AOI21_X1 U8383 ( .B1(n5120), .B2(n5121), .A(n14287), .ZN(n5101) );
  AOI221_X1 U8384 ( .B1(n14417), .B2(n5187), .C1(n14460), .C2(n2803), .A(n5127), .ZN(n5120) );
  AOI221_X1 U8385 ( .B1(n14318), .B2(n5189), .C1(n5876), .C2(n2805), .A(n5124), 
        .ZN(n5121) );
  AOI21_X1 U8386 ( .B1(n5156), .B2(n5157), .A(n5950), .ZN(n5137) );
  AOI221_X1 U8387 ( .B1(n14417), .B2(n5190), .C1(n14460), .C2(n2806), .A(n5163), .ZN(n5156) );
  AOI221_X1 U8388 ( .B1(n14318), .B2(n5194), .C1(n5876), .C2(n2810), .A(n5160), 
        .ZN(n5157) );
  AOI21_X1 U8389 ( .B1(n5192), .B2(n5193), .A(n5926), .ZN(n5173) );
  AOI221_X1 U8390 ( .B1(n14417), .B2(n5195), .C1(n14460), .C2(n2811), .A(n5199), .ZN(n5192) );
  AOI221_X1 U8391 ( .B1(n14318), .B2(n5197), .C1(n5876), .C2(n2813), .A(n5196), 
        .ZN(n5193) );
  AOI21_X1 U8392 ( .B1(n5269), .B2(n5270), .A(n14287), .ZN(n5250) );
  AOI221_X1 U8393 ( .B1(n14416), .B2(n5198), .C1(n14459), .C2(n2814), .A(n5276), .ZN(n5269) );
  AOI221_X1 U8394 ( .B1(n14317), .B2(n5202), .C1(n5878), .C2(n2818), .A(n5273), 
        .ZN(n5270) );
  AOI21_X1 U8395 ( .B1(n5305), .B2(n5306), .A(n5950), .ZN(n5286) );
  AOI221_X1 U8396 ( .B1(n14416), .B2(n5203), .C1(n14459), .C2(n2819), .A(n5312), .ZN(n5305) );
  AOI221_X1 U8397 ( .B1(n14317), .B2(n5205), .C1(n5878), .C2(n2821), .A(n5309), 
        .ZN(n5306) );
  AOI21_X1 U8398 ( .B1(n5341), .B2(n5342), .A(n5926), .ZN(n5322) );
  AOI221_X1 U8399 ( .B1(n14416), .B2(n5206), .C1(n14459), .C2(n2822), .A(n5348), .ZN(n5341) );
  AOI221_X1 U8400 ( .B1(n14317), .B2(n5219), .C1(n5889), .C2(n2835), .A(n5345), 
        .ZN(n5342) );
  AOI21_X1 U8401 ( .B1(n5418), .B2(n5419), .A(n14287), .ZN(n5399) );
  AOI221_X1 U8402 ( .B1(n14415), .B2(n5220), .C1(n14458), .C2(n2836), .A(n5425), .ZN(n5418) );
  AOI221_X1 U8403 ( .B1(n14316), .B2(n5222), .C1(n5879), .C2(n2838), .A(n5422), 
        .ZN(n5419) );
  AOI21_X1 U8404 ( .B1(n5454), .B2(n5455), .A(n5950), .ZN(n5435) );
  AOI221_X1 U8405 ( .B1(n14415), .B2(n5223), .C1(n14458), .C2(n2839), .A(n5461), .ZN(n5454) );
  AOI221_X1 U8406 ( .B1(n14316), .B2(n5227), .C1(n5890), .C2(n2843), .A(n5458), 
        .ZN(n5455) );
  AOI21_X1 U8407 ( .B1(n5490), .B2(n5491), .A(n5926), .ZN(n5471) );
  AOI221_X1 U8408 ( .B1(n14414), .B2(n5228), .C1(n14457), .C2(n2844), .A(n5497), .ZN(n5490) );
  AOI221_X1 U8409 ( .B1(n14315), .B2(n5230), .C1(n5889), .C2(n2846), .A(n5494), 
        .ZN(n5491) );
  AOI21_X1 U8410 ( .B1(n5567), .B2(n5568), .A(n14287), .ZN(n5548) );
  AOI221_X1 U8411 ( .B1(n14414), .B2(n5231), .C1(n14457), .C2(n2847), .A(n5574), .ZN(n5567) );
  AOI221_X1 U8412 ( .B1(n14315), .B2(n5235), .C1(n5892), .C2(n2851), .A(n5571), 
        .ZN(n5568) );
  AOI21_X1 U8413 ( .B1(n5603), .B2(n5604), .A(n5950), .ZN(n5584) );
  AOI221_X1 U8414 ( .B1(n14413), .B2(n5236), .C1(n14456), .C2(n2852), .A(n5610), .ZN(n5603) );
  AOI221_X1 U8415 ( .B1(n14314), .B2(n5238), .C1(n5890), .C2(n2854), .A(n5607), 
        .ZN(n5604) );
  AOI21_X1 U8416 ( .B1(n5639), .B2(n5640), .A(n5926), .ZN(n5620) );
  AOI221_X1 U8417 ( .B1(n14413), .B2(n5239), .C1(n14456), .C2(n2855), .A(n5646), .ZN(n5639) );
  AOI221_X1 U8418 ( .B1(n14314), .B2(n5243), .C1(n5890), .C2(n2859), .A(n5643), 
        .ZN(n5640) );
  AOI21_X1 U8419 ( .B1(n5716), .B2(n5717), .A(n14287), .ZN(n5697) );
  AOI221_X1 U8420 ( .B1(n14412), .B2(n5244), .C1(n14455), .C2(n2860), .A(n5723), .ZN(n5716) );
  AOI221_X1 U8421 ( .B1(n14313), .B2(n5246), .C1(n5892), .C2(n2862), .A(n5720), 
        .ZN(n5717) );
  AOI21_X1 U8422 ( .B1(n5752), .B2(n5753), .A(n5950), .ZN(n5733) );
  AOI221_X1 U8423 ( .B1(n14412), .B2(n5247), .C1(n14455), .C2(n2863), .A(n5759), .ZN(n5752) );
  AOI221_X1 U8424 ( .B1(n14313), .B2(n5255), .C1(n5892), .C2(n2871), .A(n5756), 
        .ZN(n5753) );
  AOI21_X1 U8425 ( .B1(n5788), .B2(n5789), .A(n5926), .ZN(n5769) );
  AOI221_X1 U8426 ( .B1(n14412), .B2(n5256), .C1(n14455), .C2(n2872), .A(n5795), .ZN(n5788) );
  AOI221_X1 U8427 ( .B1(n14313), .B2(n5258), .C1(n5892), .C2(n2874), .A(n5792), 
        .ZN(n5789) );
  AOI21_X1 U8428 ( .B1(n5865), .B2(n5866), .A(n14287), .ZN(n5846) );
  AOI221_X1 U8429 ( .B1(n14411), .B2(n5259), .C1(n14454), .C2(n2875), .A(n5872), .ZN(n5865) );
  AOI221_X1 U8430 ( .B1(n14312), .B2(n5263), .C1(n5893), .C2(n2879), .A(n5869), 
        .ZN(n5866) );
  AOI21_X1 U8431 ( .B1(n5903), .B2(n5904), .A(n5950), .ZN(n5882) );
  AOI221_X1 U8432 ( .B1(n14411), .B2(n5264), .C1(n14454), .C2(n2880), .A(n5910), .ZN(n5903) );
  AOI221_X1 U8433 ( .B1(n14312), .B2(n5266), .C1(n5893), .C2(n2882), .A(n5907), 
        .ZN(n5904) );
  AOI21_X1 U8434 ( .B1(n5939), .B2(n5940), .A(n5926), .ZN(n5920) );
  AOI221_X1 U8435 ( .B1(n14411), .B2(n5267), .C1(n14454), .C2(n2883), .A(n5946), .ZN(n5939) );
  AOI221_X1 U8436 ( .B1(n14312), .B2(n5271), .C1(n5868), .C2(n2887), .A(n5943), 
        .ZN(n5940) );
  AOI21_X1 U8437 ( .B1(n1245), .B2(n1246), .A(n14282), .ZN(n1214) );
  AOI221_X1 U8438 ( .B1(n14449), .B2(n5272), .C1(n14492), .C2(n2888), .A(n1253), .ZN(n1245) );
  AOI221_X1 U8439 ( .B1(n14350), .B2(n5274), .C1(n5801), .C2(n2890), .A(n1250), 
        .ZN(n1246) );
  AOI21_X1 U8440 ( .B1(n1285), .B2(n1286), .A(n5941), .ZN(n1254) );
  AOI221_X1 U8441 ( .B1(n14449), .B2(n5275), .C1(n14492), .C2(n2891), .A(n1293), .ZN(n1285) );
  AOI221_X1 U8442 ( .B1(n14350), .B2(n5279), .C1(n5801), .C2(n2895), .A(n1290), 
        .ZN(n1286) );
  AOI21_X1 U8443 ( .B1(n1325), .B2(n1326), .A(n5913), .ZN(n1294) );
  AOI221_X1 U8444 ( .B1(n14449), .B2(n5280), .C1(n14492), .C2(n2896), .A(n1333), .ZN(n1325) );
  AOI221_X1 U8445 ( .B1(n14350), .B2(n5282), .C1(n5799), .C2(n2898), .A(n1330), 
        .ZN(n1326) );
  AOI21_X1 U8446 ( .B1(n1403), .B2(n1404), .A(n14282), .ZN(n1375) );
  AOI221_X1 U8447 ( .B1(n14448), .B2(n5283), .C1(n14491), .C2(n2899), .A(n1410), .ZN(n1403) );
  AOI221_X1 U8448 ( .B1(n14349), .B2(n5291), .C1(n5802), .C2(n2907), .A(n1407), 
        .ZN(n1404) );
  AOI21_X1 U8449 ( .B1(n1439), .B2(n1440), .A(n5941), .ZN(n1411) );
  AOI221_X1 U8450 ( .B1(n14448), .B2(n5292), .C1(n14491), .C2(n2908), .A(n1446), .ZN(n1439) );
  AOI221_X1 U8451 ( .B1(n14349), .B2(n5294), .C1(n5801), .C2(n2910), .A(n1443), 
        .ZN(n1440) );
  AOI21_X1 U8452 ( .B1(n1475), .B2(n1476), .A(n5913), .ZN(n1447) );
  AOI221_X1 U8453 ( .B1(n14447), .B2(n5295), .C1(n14490), .C2(n2911), .A(n1482), .ZN(n1475) );
  AOI221_X1 U8454 ( .B1(n14348), .B2(n5299), .C1(n5801), .C2(n2915), .A(n1479), 
        .ZN(n1476) );
  AOI21_X1 U8455 ( .B1(n1552), .B2(n1553), .A(n14282), .ZN(n1524) );
  AOI221_X1 U8456 ( .B1(n14447), .B2(n5300), .C1(n14490), .C2(n2916), .A(n1559), .ZN(n1552) );
  AOI221_X1 U8457 ( .B1(n14348), .B2(n5302), .C1(n5815), .C2(n2918), .A(n1556), 
        .ZN(n1553) );
  AOI21_X1 U8458 ( .B1(n1588), .B2(n1589), .A(n5941), .ZN(n1560) );
  AOI221_X1 U8459 ( .B1(n14447), .B2(n5303), .C1(n14490), .C2(n2919), .A(n1595), .ZN(n1588) );
  AOI221_X1 U8460 ( .B1(n14348), .B2(n5307), .C1(n5802), .C2(n2923), .A(n1592), 
        .ZN(n1589) );
  AOI21_X1 U8461 ( .B1(n1624), .B2(n1625), .A(n5913), .ZN(n1596) );
  AOI221_X1 U8462 ( .B1(n14446), .B2(n5308), .C1(n14489), .C2(n2924), .A(n1631), .ZN(n1624) );
  AOI221_X1 U8463 ( .B1(n14347), .B2(n5310), .C1(n5816), .C2(n2926), .A(n1628), 
        .ZN(n1625) );
  AOI21_X1 U8464 ( .B1(n1701), .B2(n1702), .A(n14282), .ZN(n1673) );
  AOI221_X1 U8465 ( .B1(n14446), .B2(n5311), .C1(n14489), .C2(n2927), .A(n1708), .ZN(n1701) );
  AOI221_X1 U8466 ( .B1(n14347), .B2(n5315), .C1(n5815), .C2(n2931), .A(n1705), 
        .ZN(n1702) );
  AOI21_X1 U8467 ( .B1(n1737), .B2(n1738), .A(n5941), .ZN(n1709) );
  AOI221_X1 U8468 ( .B1(n14445), .B2(n5316), .C1(n14488), .C2(n2932), .A(n1744), .ZN(n1737) );
  AOI221_X1 U8469 ( .B1(n14346), .B2(n5318), .C1(n5818), .C2(n2934), .A(n1741), 
        .ZN(n1738) );
  AOI21_X1 U8470 ( .B1(n1773), .B2(n1774), .A(n5913), .ZN(n1745) );
  AOI221_X1 U8471 ( .B1(n14445), .B2(n5319), .C1(n14488), .C2(n2935), .A(n1780), .ZN(n1773) );
  AOI221_X1 U8472 ( .B1(n14346), .B2(n5327), .C1(n5818), .C2(n2943), .A(n1777), 
        .ZN(n1774) );
  AOI21_X1 U8473 ( .B1(n1850), .B2(n1851), .A(n14282), .ZN(n1822) );
  AOI221_X1 U8474 ( .B1(n14444), .B2(n5328), .C1(n14487), .C2(n2944), .A(n1857), .ZN(n1850) );
  AOI221_X1 U8475 ( .B1(n14345), .B2(n5330), .C1(n5816), .C2(n2946), .A(n1854), 
        .ZN(n1851) );
  AOI21_X1 U8476 ( .B1(n1886), .B2(n1887), .A(n5941), .ZN(n1858) );
  AOI221_X1 U8477 ( .B1(n14444), .B2(n5331), .C1(n14487), .C2(n2947), .A(n1893), .ZN(n1886) );
  AOI221_X1 U8478 ( .B1(n14345), .B2(n5335), .C1(n5819), .C2(n2951), .A(n1890), 
        .ZN(n1887) );
  AOI21_X1 U8479 ( .B1(n1922), .B2(n1923), .A(n5913), .ZN(n1894) );
  AOI221_X1 U8480 ( .B1(n14444), .B2(n5336), .C1(n14487), .C2(n2952), .A(n1929), .ZN(n1922) );
  AOI221_X1 U8481 ( .B1(n14345), .B2(n5338), .C1(n5819), .C2(n2954), .A(n1926), 
        .ZN(n1923) );
  AOI21_X1 U8482 ( .B1(n1999), .B2(n2000), .A(n14282), .ZN(n1971) );
  AOI221_X1 U8483 ( .B1(n14443), .B2(n5339), .C1(n14486), .C2(n2955), .A(n2006), .ZN(n1999) );
  AOI221_X1 U8484 ( .B1(n14344), .B2(n5343), .C1(n5823), .C2(n2959), .A(n2003), 
        .ZN(n2000) );
  AOI21_X1 U8485 ( .B1(n2035), .B2(n2036), .A(n5941), .ZN(n2007) );
  AOI221_X1 U8486 ( .B1(n14443), .B2(n5344), .C1(n14486), .C2(n2960), .A(n2042), .ZN(n2035) );
  AOI221_X1 U8487 ( .B1(n14344), .B2(n5346), .C1(n5823), .C2(n2962), .A(n2039), 
        .ZN(n2036) );
  AOI21_X1 U8488 ( .B1(n2071), .B2(n2072), .A(n5913), .ZN(n2043) );
  AOI221_X1 U8489 ( .B1(n14443), .B2(n5347), .C1(n14486), .C2(n2963), .A(n2078), .ZN(n2071) );
  AOI221_X1 U8490 ( .B1(n14344), .B2(n5351), .C1(n5819), .C2(n2967), .A(n2075), 
        .ZN(n2072) );
  AOI21_X1 U8491 ( .B1(n2148), .B2(n2149), .A(n14282), .ZN(n2120) );
  AOI221_X1 U8492 ( .B1(n14442), .B2(n5352), .C1(n14485), .C2(n2968), .A(n2155), .ZN(n2148) );
  AOI221_X1 U8493 ( .B1(n14343), .B2(n5354), .C1(n5824), .C2(n2970), .A(n2152), 
        .ZN(n2149) );
  AOI21_X1 U8494 ( .B1(n2184), .B2(n2185), .A(n5941), .ZN(n2156) );
  AOI221_X1 U8495 ( .B1(n14442), .B2(n5355), .C1(n14485), .C2(n2971), .A(n2191), .ZN(n2184) );
  AOI221_X1 U8496 ( .B1(n14343), .B2(n5368), .C1(n5823), .C2(n2984), .A(n2188), 
        .ZN(n2185) );
  AOI21_X1 U8497 ( .B1(n2220), .B2(n2221), .A(n5913), .ZN(n2192) );
  AOI221_X1 U8498 ( .B1(n14441), .B2(n5369), .C1(n14484), .C2(n2985), .A(n2227), .ZN(n2220) );
  AOI221_X1 U8499 ( .B1(n14342), .B2(n5371), .C1(n5826), .C2(n2987), .A(n2224), 
        .ZN(n2221) );
  AOI21_X1 U8500 ( .B1(n2297), .B2(n2298), .A(n14282), .ZN(n2269) );
  AOI221_X1 U8501 ( .B1(n14441), .B2(n5372), .C1(n14484), .C2(n2988), .A(n2304), .ZN(n2297) );
  AOI221_X1 U8502 ( .B1(n14342), .B2(n5376), .C1(n5824), .C2(n2992), .A(n2301), 
        .ZN(n2298) );
  AOI21_X1 U8503 ( .B1(n2333), .B2(n2334), .A(n5941), .ZN(n2305) );
  AOI221_X1 U8504 ( .B1(n14440), .B2(n5377), .C1(n14483), .C2(n2993), .A(n2340), .ZN(n2333) );
  AOI221_X1 U8505 ( .B1(n14341), .B2(n5379), .C1(n5824), .C2(n2995), .A(n2337), 
        .ZN(n2334) );
  AOI21_X1 U8506 ( .B1(n2369), .B2(n2370), .A(n5913), .ZN(n2341) );
  AOI221_X1 U8507 ( .B1(n14440), .B2(n5380), .C1(n14483), .C2(n2996), .A(n2376), .ZN(n2369) );
  AOI221_X1 U8508 ( .B1(n14341), .B2(n5384), .C1(n5818), .C2(n3000), .A(n2373), 
        .ZN(n2370) );
  AOI21_X1 U8509 ( .B1(n2446), .B2(n2447), .A(n14282), .ZN(n2418) );
  AOI221_X1 U8510 ( .B1(n14439), .B2(n5385), .C1(n14482), .C2(n3001), .A(n2453), .ZN(n2446) );
  AOI221_X1 U8511 ( .B1(n14340), .B2(n5387), .C1(n5827), .C2(n3003), .A(n2450), 
        .ZN(n2447) );
  AOI21_X1 U8512 ( .B1(n2482), .B2(n2483), .A(n5941), .ZN(n2454) );
  AOI221_X1 U8513 ( .B1(n14439), .B2(n5388), .C1(n14482), .C2(n3004), .A(n2489), .ZN(n2482) );
  AOI221_X1 U8514 ( .B1(n14340), .B2(n5392), .C1(n5827), .C2(n3008), .A(n2486), 
        .ZN(n2483) );
  AOI21_X1 U8515 ( .B1(n2518), .B2(n2519), .A(n5913), .ZN(n2490) );
  AOI221_X1 U8516 ( .B1(n14439), .B2(n5393), .C1(n14482), .C2(n3009), .A(n2525), .ZN(n2518) );
  AOI221_X1 U8517 ( .B1(n14340), .B2(n5395), .C1(n5827), .C2(n3011), .A(n2522), 
        .ZN(n2519) );
  AOI21_X1 U8518 ( .B1(n2595), .B2(n2596), .A(n14282), .ZN(n2567) );
  AOI221_X1 U8519 ( .B1(n14438), .B2(n5396), .C1(n14481), .C2(n3012), .A(n2602), .ZN(n2595) );
  AOI221_X1 U8520 ( .B1(n14339), .B2(n5404), .C1(n5831), .C2(n3020), .A(n2599), 
        .ZN(n2596) );
  AOI21_X1 U8521 ( .B1(n2631), .B2(n2632), .A(n5941), .ZN(n2603) );
  AOI221_X1 U8522 ( .B1(n14438), .B2(n5405), .C1(n14481), .C2(n3021), .A(n2638), .ZN(n2631) );
  AOI221_X1 U8523 ( .B1(n14339), .B2(n5407), .C1(n5831), .C2(n3023), .A(n2635), 
        .ZN(n2632) );
  AOI21_X1 U8524 ( .B1(n2667), .B2(n2668), .A(n5913), .ZN(n2639) );
  AOI221_X1 U8525 ( .B1(n14438), .B2(n5408), .C1(n14481), .C2(n3024), .A(n2674), .ZN(n2667) );
  AOI221_X1 U8526 ( .B1(n14339), .B2(n5412), .C1(n5834), .C2(n3028), .A(n2671), 
        .ZN(n2668) );
  AOI21_X1 U8527 ( .B1(n2744), .B2(n2745), .A(n14282), .ZN(n2716) );
  AOI221_X1 U8529 ( .B1(n14437), .B2(n5413), .C1(n14480), .C2(n3029), .A(n2751), .ZN(n2744) );
  AOI221_X1 U8530 ( .B1(n14338), .B2(n5415), .C1(n5832), .C2(n3031), .A(n2748), 
        .ZN(n2745) );
  AOI21_X1 U8531 ( .B1(n2780), .B2(n2781), .A(n5941), .ZN(n2752) );
  AOI221_X1 U8532 ( .B1(n14437), .B2(n5416), .C1(n14480), .C2(n3032), .A(n2787), .ZN(n2780) );
  AOI221_X1 U8533 ( .B1(n14338), .B2(n5420), .C1(n5835), .C2(n3036), .A(n2784), 
        .ZN(n2781) );
  AOI21_X1 U8534 ( .B1(n2816), .B2(n2817), .A(n5913), .ZN(n2788) );
  AOI221_X1 U8535 ( .B1(n14436), .B2(n5421), .C1(n14479), .C2(n3037), .A(n2823), .ZN(n2816) );
  AOI221_X1 U8536 ( .B1(n14337), .B2(n5423), .C1(n5834), .C2(n3039), .A(n2820), 
        .ZN(n2817) );
  AOI21_X1 U8537 ( .B1(n2893), .B2(n2894), .A(n14282), .ZN(n2865) );
  AOI221_X1 U8538 ( .B1(n14436), .B2(n5424), .C1(n14479), .C2(n3040), .A(n2900), .ZN(n2893) );
  AOI221_X1 U8539 ( .B1(n14337), .B2(n5428), .C1(n5834), .C2(n3044), .A(n2897), 
        .ZN(n2894) );
  AOI21_X1 U8540 ( .B1(n2929), .B2(n2930), .A(n5941), .ZN(n2901) );
  AOI221_X1 U8541 ( .B1(n14435), .B2(n5429), .C1(n14478), .C2(n3045), .A(n2936), .ZN(n2929) );
  AOI221_X1 U8542 ( .B1(n14336), .B2(n5431), .C1(n5835), .C2(n3047), .A(n2933), 
        .ZN(n2930) );
  AOI21_X1 U8543 ( .B1(n2965), .B2(n2966), .A(n5913), .ZN(n2937) );
  AOI221_X1 U8544 ( .B1(n14435), .B2(n5432), .C1(n14478), .C2(n3048), .A(n2972), .ZN(n2965) );
  AOI221_X1 U8545 ( .B1(n14336), .B2(n5440), .C1(n5835), .C2(n3056), .A(n2969), 
        .ZN(n2966) );
  AOI21_X1 U8546 ( .B1(n3042), .B2(n3043), .A(n14282), .ZN(n3014) );
  AOI221_X1 U8547 ( .B1(n14435), .B2(n5441), .C1(n14478), .C2(n3057), .A(n3049), .ZN(n3042) );
  AOI221_X1 U8548 ( .B1(n14336), .B2(n5443), .C1(n5840), .C2(n3059), .A(n3046), 
        .ZN(n3043) );
  AOI21_X1 U8549 ( .B1(n3078), .B2(n3079), .A(n5941), .ZN(n3050) );
  AOI221_X1 U8550 ( .B1(n14434), .B2(n5444), .C1(n14477), .C2(n3060), .A(n3085), .ZN(n3078) );
  AOI221_X1 U8551 ( .B1(n14335), .B2(n5448), .C1(n5839), .C2(n3064), .A(n3082), 
        .ZN(n3079) );
  AOI21_X1 U8552 ( .B1(n3114), .B2(n3115), .A(n5913), .ZN(n3086) );
  AOI221_X1 U8553 ( .B1(n14434), .B2(n5449), .C1(n14477), .C2(n3065), .A(n3121), .ZN(n3114) );
  AOI221_X1 U8554 ( .B1(n14335), .B2(n5451), .C1(n5839), .C2(n3067), .A(n3118), 
        .ZN(n3115) );
  AOI21_X1 U8555 ( .B1(n3191), .B2(n3192), .A(n14283), .ZN(n3163) );
  AOI221_X1 U8556 ( .B1(n14433), .B2(n5452), .C1(n14476), .C2(n3068), .A(n3198), .ZN(n3191) );
  AOI221_X1 U8557 ( .B1(n14334), .B2(n5456), .C1(n5840), .C2(n3072), .A(n3195), 
        .ZN(n3192) );
  AOI21_X1 U8558 ( .B1(n3227), .B2(n3228), .A(n5942), .ZN(n3199) );
  AOI221_X1 U8559 ( .B1(n14433), .B2(n5457), .C1(n14476), .C2(n3073), .A(n3234), .ZN(n3227) );
  AOI221_X1 U8560 ( .B1(n14334), .B2(n5459), .C1(n5840), .C2(n3075), .A(n3231), 
        .ZN(n3228) );
  AOI21_X1 U8561 ( .B1(n3263), .B2(n3264), .A(n5914), .ZN(n3235) );
  AOI221_X1 U8562 ( .B1(n14433), .B2(n5460), .C1(n14476), .C2(n3076), .A(n3270), .ZN(n3263) );
  AOI221_X1 U8563 ( .B1(n14334), .B2(n5464), .C1(n5843), .C2(n3080), .A(n3267), 
        .ZN(n3264) );
  AOI21_X1 U8564 ( .B1(n3340), .B2(n3341), .A(n14283), .ZN(n3312) );
  AOI221_X1 U8565 ( .B1(n14432), .B2(n5465), .C1(n14475), .C2(n3081), .A(n3347), .ZN(n3340) );
  AOI221_X1 U8566 ( .B1(n14333), .B2(n5467), .C1(n5842), .C2(n3083), .A(n3344), 
        .ZN(n3341) );
  AOI21_X1 U8567 ( .B1(n3376), .B2(n3377), .A(n5942), .ZN(n3348) );
  AOI221_X1 U8568 ( .B1(n14432), .B2(n5468), .C1(n14475), .C2(n3084), .A(n3383), .ZN(n3376) );
  AOI221_X1 U8569 ( .B1(n14333), .B2(n5476), .C1(n5842), .C2(n3092), .A(n3380), 
        .ZN(n3377) );
  AOI21_X1 U8570 ( .B1(n3412), .B2(n3413), .A(n5914), .ZN(n3384) );
  AOI221_X1 U8571 ( .B1(n14431), .B2(n5477), .C1(n14474), .C2(n3093), .A(n3419), .ZN(n3412) );
  AOI221_X1 U8572 ( .B1(n14332), .B2(n5479), .C1(n5843), .C2(n3095), .A(n3416), 
        .ZN(n3413) );
  AOI21_X1 U8573 ( .B1(n3489), .B2(n3490), .A(n14283), .ZN(n3461) );
  AOI221_X1 U8574 ( .B1(n14431), .B2(n5480), .C1(n14474), .C2(n3096), .A(n3496), .ZN(n3489) );
  AOI221_X1 U8575 ( .B1(n14332), .B2(n5484), .C1(n5843), .C2(n3100), .A(n3493), 
        .ZN(n3490) );
  AOI21_X1 U8576 ( .B1(n3525), .B2(n3526), .A(n5942), .ZN(n3497) );
  AOI221_X1 U8577 ( .B1(n14431), .B2(n5485), .C1(n14474), .C2(n3101), .A(n3532), .ZN(n3525) );
  AOI221_X1 U8578 ( .B1(n14332), .B2(n5487), .C1(n5799), .C2(n3103), .A(n3529), 
        .ZN(n3526) );
  AOI21_X1 U8579 ( .B1(n3561), .B2(n3562), .A(n5914), .ZN(n3533) );
  AOI221_X1 U8580 ( .B1(n14430), .B2(n5488), .C1(n14473), .C2(n3104), .A(n3568), .ZN(n3561) );
  AOI221_X1 U8581 ( .B1(n14331), .B2(n5492), .C1(n5852), .C2(n3108), .A(n3565), 
        .ZN(n3562) );
  AOI21_X1 U8582 ( .B1(n3638), .B2(n3639), .A(n14283), .ZN(n3610) );
  AOI221_X1 U8583 ( .B1(n14430), .B2(n5493), .C1(n14473), .C2(n3109), .A(n3645), .ZN(n3638) );
  AOI221_X1 U8584 ( .B1(n14331), .B2(n5495), .C1(n5851), .C2(n3111), .A(n3642), 
        .ZN(n3639) );
  AOI21_X1 U8585 ( .B1(n3674), .B2(n3675), .A(n5942), .ZN(n3646) );
  AOI221_X1 U8586 ( .B1(n14429), .B2(n5496), .C1(n14472), .C2(n3112), .A(n3681), .ZN(n3674) );
  AOI221_X1 U8587 ( .B1(n14330), .B2(n5500), .C1(n5854), .C2(n3116), .A(n3678), 
        .ZN(n3675) );
  AOI21_X1 U8588 ( .B1(n3710), .B2(n3711), .A(n5914), .ZN(n3682) );
  AOI221_X1 U8589 ( .B1(n14429), .B2(n5501), .C1(n14472), .C2(n3117), .A(n3717), .ZN(n3710) );
  AOI221_X1 U8590 ( .B1(n14330), .B2(n5503), .C1(n5854), .C2(n3119), .A(n3714), 
        .ZN(n3711) );
  AOI21_X1 U8591 ( .B1(n3787), .B2(n3788), .A(n14283), .ZN(n3759) );
  AOI221_X1 U8592 ( .B1(n14428), .B2(n5504), .C1(n14471), .C2(n3120), .A(n3794), .ZN(n3787) );
  AOI221_X1 U8593 ( .B1(n14329), .B2(n5517), .C1(n5852), .C2(n3133), .A(n3791), 
        .ZN(n3788) );
  AOI21_X1 U8594 ( .B1(n3823), .B2(n3824), .A(n5942), .ZN(n3795) );
  AOI221_X1 U8595 ( .B1(n14428), .B2(n5518), .C1(n14471), .C2(n3134), .A(n3830), .ZN(n3823) );
  AOI221_X1 U8596 ( .B1(n14329), .B2(n5520), .C1(n5855), .C2(n3136), .A(n3827), 
        .ZN(n3824) );
  AOI21_X1 U8597 ( .B1(n3859), .B2(n3860), .A(n5914), .ZN(n3831) );
  AOI221_X1 U8598 ( .B1(n14428), .B2(n5521), .C1(n14471), .C2(n3137), .A(n3866), .ZN(n3859) );
  AOI221_X1 U8599 ( .B1(n14329), .B2(n5525), .C1(n5855), .C2(n3141), .A(n3863), 
        .ZN(n3860) );
  AOI21_X1 U8600 ( .B1(n3936), .B2(n3937), .A(n14283), .ZN(n3908) );
  AOI221_X1 U8601 ( .B1(n14427), .B2(n5526), .C1(n14470), .C2(n3142), .A(n3943), .ZN(n3936) );
  AOI221_X1 U8602 ( .B1(n14328), .B2(n5528), .C1(n5859), .C2(n3144), .A(n3940), 
        .ZN(n3937) );
  AOI21_X1 U8603 ( .B1(n3972), .B2(n3973), .A(n5942), .ZN(n3944) );
  AOI221_X1 U8604 ( .B1(n14427), .B2(n5529), .C1(n14470), .C2(n3145), .A(n3979), .ZN(n3972) );
  AOI221_X1 U8605 ( .B1(n14328), .B2(n5533), .C1(n5859), .C2(n3149), .A(n3976), 
        .ZN(n3973) );
  AOI21_X1 U8606 ( .B1(n4008), .B2(n4009), .A(n5914), .ZN(n3980) );
  AOI221_X1 U8607 ( .B1(n14427), .B2(n5534), .C1(n14470), .C2(n3150), .A(n4015), .ZN(n4008) );
  AOI221_X1 U8608 ( .B1(n14328), .B2(n5536), .C1(n5855), .C2(n3152), .A(n4012), 
        .ZN(n4009) );
  AOI21_X1 U8609 ( .B1(n4085), .B2(n4086), .A(n14283), .ZN(n4057) );
  AOI221_X1 U8610 ( .B1(n14426), .B2(n5537), .C1(n14469), .C2(n3153), .A(n4092), .ZN(n4085) );
  AOI221_X1 U8611 ( .B1(n14327), .B2(n5541), .C1(n5860), .C2(n3157), .A(n4089), 
        .ZN(n4086) );
  AOI21_X1 U8612 ( .B1(n4121), .B2(n4122), .A(n5942), .ZN(n4093) );
  AOI221_X1 U8613 ( .B1(n14426), .B2(n5542), .C1(n14469), .C2(n3158), .A(n4128), .ZN(n4121) );
  AOI221_X1 U8614 ( .B1(n14327), .B2(n5544), .C1(n5859), .C2(n3160), .A(n4125), 
        .ZN(n4122) );
  AOI21_X1 U8615 ( .B1(n4157), .B2(n4158), .A(n5914), .ZN(n4129) );
  AOI221_X1 U8616 ( .B1(n14425), .B2(n5545), .C1(n14468), .C2(n3161), .A(n4164), .ZN(n4157) );
  AOI221_X1 U8617 ( .B1(n14326), .B2(n5553), .C1(n5862), .C2(n3169), .A(n4161), 
        .ZN(n4158) );
  AOI21_X1 U8618 ( .B1(n4234), .B2(n4235), .A(n14283), .ZN(n4206) );
  AOI221_X1 U8619 ( .B1(n14425), .B2(n5554), .C1(n14468), .C2(n3170), .A(n4241), .ZN(n4234) );
  AOI221_X1 U8620 ( .B1(n14326), .B2(n5556), .C1(n5860), .C2(n3172), .A(n4238), 
        .ZN(n4235) );
  AOI21_X1 U8621 ( .B1(n4270), .B2(n4271), .A(n5942), .ZN(n4242) );
  AOI221_X1 U8622 ( .B1(n14424), .B2(n5557), .C1(n14467), .C2(n3173), .A(n4277), .ZN(n4270) );
  AOI221_X1 U8623 ( .B1(n14325), .B2(n5561), .C1(n5863), .C2(n3177), .A(n4274), 
        .ZN(n4271) );
  AOI21_X1 U8624 ( .B1(n4306), .B2(n4307), .A(n5914), .ZN(n4278) );
  AOI221_X1 U8625 ( .B1(n14424), .B2(n5562), .C1(n14467), .C2(n3178), .A(n4313), .ZN(n4306) );
  AOI221_X1 U8626 ( .B1(n14325), .B2(n5564), .C1(n5863), .C2(n3180), .A(n4310), 
        .ZN(n4307) );
  AOI21_X1 U8627 ( .B1(n4383), .B2(n4384), .A(n14283), .ZN(n4355) );
  AOI221_X1 U8628 ( .B1(n14423), .B2(n5565), .C1(n14466), .C2(n3181), .A(n4390), .ZN(n4383) );
  AOI221_X1 U8629 ( .B1(n14324), .B2(n5569), .C1(n5862), .C2(n3185), .A(n4387), 
        .ZN(n4384) );
  AOI21_X1 U8630 ( .B1(n4419), .B2(n4420), .A(n5942), .ZN(n4391) );
  AOI221_X1 U8631 ( .B1(n14423), .B2(n5570), .C1(n14466), .C2(n3186), .A(n4426), .ZN(n4419) );
  AOI221_X1 U8632 ( .B1(n14324), .B2(n5572), .C1(n5867), .C2(n3188), .A(n4423), 
        .ZN(n4420) );
  AOI21_X1 U8633 ( .B1(n4455), .B2(n4456), .A(n5914), .ZN(n4427) );
  AOI221_X1 U8634 ( .B1(n14423), .B2(n5573), .C1(n14466), .C2(n3189), .A(n4462), .ZN(n4455) );
  AOI221_X1 U8635 ( .B1(n14324), .B2(n5577), .C1(n5867), .C2(n3193), .A(n4459), 
        .ZN(n4456) );
  AOI21_X1 U8636 ( .B1(n4532), .B2(n4533), .A(n14283), .ZN(n4504) );
  AOI221_X1 U8637 ( .B1(n14422), .B2(n5578), .C1(n14465), .C2(n3194), .A(n4539), .ZN(n4532) );
  AOI221_X1 U8638 ( .B1(n14323), .B2(n5580), .C1(n5868), .C2(n3196), .A(n4536), 
        .ZN(n4533) );
  AOI21_X1 U8639 ( .B1(n4568), .B2(n4569), .A(n5942), .ZN(n4540) );
  AOI221_X1 U8640 ( .B1(n14422), .B2(n5581), .C1(n14465), .C2(n3197), .A(n4575), .ZN(n4568) );
  AOI221_X1 U8641 ( .B1(n14323), .B2(n5589), .C1(n5868), .C2(n3205), .A(n4572), 
        .ZN(n4569) );
  AOI21_X1 U8642 ( .B1(n4604), .B2(n4605), .A(n5914), .ZN(n4576) );
  AOI221_X1 U8643 ( .B1(n14422), .B2(n5590), .C1(n14465), .C2(n3206), .A(n4611), .ZN(n4604) );
  AOI221_X1 U8644 ( .B1(n14323), .B2(n5592), .C1(n5867), .C2(n3208), .A(n4608), 
        .ZN(n4605) );
  AOI21_X1 U8645 ( .B1(n4681), .B2(n4682), .A(n14283), .ZN(n4653) );
  AOI221_X1 U8646 ( .B1(n14421), .B2(n5593), .C1(n14464), .C2(n3209), .A(n4688), .ZN(n4681) );
  AOI221_X1 U8647 ( .B1(n14322), .B2(n5597), .C1(n5870), .C2(n3213), .A(n4685), 
        .ZN(n4682) );
  AOI21_X1 U8648 ( .B1(n4717), .B2(n4718), .A(n5942), .ZN(n4689) );
  AOI221_X1 U8649 ( .B1(n14421), .B2(n5598), .C1(n14464), .C2(n3214), .A(n4724), .ZN(n4717) );
  AOI221_X1 U8650 ( .B1(n14322), .B2(n5600), .C1(n5868), .C2(n3216), .A(n4721), 
        .ZN(n4718) );
  AOI21_X1 U8651 ( .B1(n4753), .B2(n4754), .A(n5914), .ZN(n4725) );
  AOI221_X1 U8652 ( .B1(n14420), .B2(n5601), .C1(n14463), .C2(n3217), .A(n4760), .ZN(n4753) );
  AOI221_X1 U8653 ( .B1(n14321), .B2(n5605), .C1(n5870), .C2(n3221), .A(n4757), 
        .ZN(n4754) );
  AOI21_X1 U8654 ( .B1(n4830), .B2(n4831), .A(n14283), .ZN(n4802) );
  AOI221_X1 U8655 ( .B1(n14420), .B2(n5606), .C1(n14463), .C2(n3222), .A(n4837), .ZN(n4830) );
  AOI221_X1 U8656 ( .B1(n14321), .B2(n5608), .C1(n5826), .C2(n3224), .A(n4834), 
        .ZN(n4831) );
  AOI21_X1 U8657 ( .B1(n4866), .B2(n4867), .A(n5942), .ZN(n4838) );
  AOI221_X1 U8658 ( .B1(n14419), .B2(n5609), .C1(n14462), .C2(n3225), .A(n4873), .ZN(n4866) );
  AOI221_X1 U8659 ( .B1(n14320), .B2(n5613), .C1(n5871), .C2(n3229), .A(n4870), 
        .ZN(n4867) );
  AOI21_X1 U8660 ( .B1(n4902), .B2(n4903), .A(n5914), .ZN(n4874) );
  AOI221_X1 U8661 ( .B1(n14419), .B2(n5614), .C1(n14462), .C2(n3230), .A(n4909), .ZN(n4902) );
  AOI221_X1 U8662 ( .B1(n14320), .B2(n5616), .C1(n5871), .C2(n3232), .A(n4906), 
        .ZN(n4903) );
  AOI21_X1 U8663 ( .B1(n4979), .B2(n4980), .A(n14283), .ZN(n4951) );
  AOI221_X1 U8664 ( .B1(n14419), .B2(n5617), .C1(n14462), .C2(n3233), .A(n4986), .ZN(n4979) );
  AOI221_X1 U8665 ( .B1(n14320), .B2(n5625), .C1(n5876), .C2(n3241), .A(n4983), 
        .ZN(n4980) );
  AOI21_X1 U8666 ( .B1(n5015), .B2(n5016), .A(n5942), .ZN(n4987) );
  AOI221_X1 U8667 ( .B1(n14418), .B2(n5626), .C1(n14461), .C2(n3242), .A(n5022), .ZN(n5015) );
  AOI221_X1 U8668 ( .B1(n14319), .B2(n5628), .C1(n5875), .C2(n3244), .A(n5019), 
        .ZN(n5016) );
  AOI21_X1 U8669 ( .B1(n5051), .B2(n5052), .A(n5914), .ZN(n5023) );
  AOI221_X1 U8670 ( .B1(n14418), .B2(n5629), .C1(n14461), .C2(n3245), .A(n5058), .ZN(n5051) );
  AOI221_X1 U8671 ( .B1(n14319), .B2(n5633), .C1(n5875), .C2(n3249), .A(n5055), 
        .ZN(n5052) );
  AOI21_X1 U8672 ( .B1(n5128), .B2(n5129), .A(n14284), .ZN(n5100) );
  AOI221_X1 U8673 ( .B1(n14417), .B2(n5634), .C1(n14460), .C2(n3250), .A(n5135), .ZN(n5128) );
  AOI221_X1 U8674 ( .B1(n14318), .B2(n5636), .C1(n5876), .C2(n3252), .A(n5132), 
        .ZN(n5129) );
  AOI21_X1 U8675 ( .B1(n5164), .B2(n5165), .A(n5944), .ZN(n5136) );
  AOI221_X1 U8676 ( .B1(n14417), .B2(n5637), .C1(n14460), .C2(n3253), .A(n5171), .ZN(n5164) );
  AOI221_X1 U8677 ( .B1(n14318), .B2(n5641), .C1(n5876), .C2(n3257), .A(n5168), 
        .ZN(n5165) );
  AOI21_X1 U8678 ( .B1(n5200), .B2(n5201), .A(n5916), .ZN(n5172) );
  AOI221_X1 U8679 ( .B1(n14417), .B2(n5642), .C1(n14460), .C2(n3258), .A(n5207), .ZN(n5200) );
  AOI221_X1 U8681 ( .B1(n14318), .B2(n5644), .C1(n5879), .C2(n3260), .A(n5204), 
        .ZN(n5201) );
  AOI21_X1 U8682 ( .B1(n5277), .B2(n5278), .A(n14284), .ZN(n5249) );
  AOI221_X1 U8683 ( .B1(n14416), .B2(n5645), .C1(n14459), .C2(n3261), .A(n5284), .ZN(n5277) );
  AOI221_X1 U8684 ( .B1(n14317), .B2(n5649), .C1(n5878), .C2(n3265), .A(n5281), 
        .ZN(n5278) );
  AOI21_X1 U8685 ( .B1(n5313), .B2(n5314), .A(n5944), .ZN(n5285) );
  AOI221_X1 U8686 ( .B1(n14416), .B2(n5650), .C1(n14459), .C2(n3266), .A(n5320), .ZN(n5313) );
  AOI221_X1 U8687 ( .B1(n14317), .B2(n5652), .C1(n5878), .C2(n3268), .A(n5317), 
        .ZN(n5314) );
  AOI21_X1 U8688 ( .B1(n5349), .B2(n5350), .A(n5916), .ZN(n5321) );
  AOI221_X1 U8689 ( .B1(n14415), .B2(n5653), .C1(n14458), .C2(n3269), .A(n5356), .ZN(n5349) );
  AOI221_X1 U8690 ( .B1(n14316), .B2(n5666), .C1(n5879), .C2(n3282), .A(n5353), 
        .ZN(n5350) );
  AOI21_X1 U8691 ( .B1(n5426), .B2(n5427), .A(n14284), .ZN(n5398) );
  AOI221_X1 U8692 ( .B1(n14415), .B2(n5667), .C1(n14458), .C2(n3283), .A(n5433), .ZN(n5426) );
  AOI221_X1 U8693 ( .B1(n14316), .B2(n5669), .C1(n5879), .C2(n3285), .A(n5430), 
        .ZN(n5427) );
  AOI21_X1 U8694 ( .B1(n5462), .B2(n5463), .A(n5944), .ZN(n5434) );
  AOI221_X1 U8695 ( .B1(n14415), .B2(n5670), .C1(n14458), .C2(n3286), .A(n5469), .ZN(n5462) );
  AOI221_X1 U8696 ( .B1(n14316), .B2(n5674), .C1(n5890), .C2(n3290), .A(n5466), 
        .ZN(n5463) );
  AOI21_X1 U8697 ( .B1(n5498), .B2(n5499), .A(n5916), .ZN(n5470) );
  AOI221_X1 U8698 ( .B1(n14414), .B2(n5675), .C1(n14457), .C2(n3291), .A(n5505), .ZN(n5498) );
  AOI221_X1 U8699 ( .B1(n14315), .B2(n5677), .C1(n5889), .C2(n3293), .A(n5502), 
        .ZN(n5499) );
  AOI21_X1 U8700 ( .B1(n5575), .B2(n5576), .A(n14284), .ZN(n5547) );
  AOI221_X1 U8701 ( .B1(n14414), .B2(n5678), .C1(n14457), .C2(n3294), .A(n5582), .ZN(n5575) );
  AOI221_X1 U8702 ( .B1(n14315), .B2(n5682), .C1(n5892), .C2(n3298), .A(n5579), 
        .ZN(n5576) );
  AOI21_X1 U8703 ( .B1(n5611), .B2(n5612), .A(n5944), .ZN(n5583) );
  AOI221_X1 U8704 ( .B1(n14413), .B2(n5683), .C1(n14456), .C2(n3299), .A(n5618), .ZN(n5611) );
  AOI221_X1 U8705 ( .B1(n14314), .B2(n5685), .C1(n5890), .C2(n3301), .A(n5615), 
        .ZN(n5612) );
  AOI21_X1 U8706 ( .B1(n5647), .B2(n5648), .A(n5916), .ZN(n5619) );
  AOI221_X1 U8707 ( .B1(n14413), .B2(n5686), .C1(n14456), .C2(n3302), .A(n5654), .ZN(n5647) );
  AOI221_X1 U8708 ( .B1(n14314), .B2(n5690), .C1(n5890), .C2(n3306), .A(n5651), 
        .ZN(n5648) );
  AOI21_X1 U8709 ( .B1(n5724), .B2(n5725), .A(n14284), .ZN(n5696) );
  AOI221_X1 U8710 ( .B1(n14412), .B2(n5691), .C1(n14455), .C2(n3307), .A(n5731), .ZN(n5724) );
  AOI221_X1 U8711 ( .B1(n14313), .B2(n5693), .C1(n5892), .C2(n3309), .A(n5728), 
        .ZN(n5725) );
  AOI21_X1 U8712 ( .B1(n5760), .B2(n5761), .A(n5944), .ZN(n5732) );
  AOI221_X1 U8713 ( .B1(n14412), .B2(n5694), .C1(n14455), .C2(n3310), .A(n5767), .ZN(n5760) );
  AOI221_X1 U8714 ( .B1(n14313), .B2(n5702), .C1(n5892), .C2(n3318), .A(n5764), 
        .ZN(n5761) );
  AOI21_X1 U8715 ( .B1(n5837), .B2(n5838), .A(n14296), .ZN(n5809) );
  AOI221_X1 U8716 ( .B1(n14411), .B2(n5703), .C1(n14454), .C2(n3319), .A(n5844), .ZN(n5837) );
  AOI221_X1 U8717 ( .B1(n14312), .B2(n5705), .C1(n5893), .C2(n3321), .A(n5841), 
        .ZN(n5838) );
  AOI21_X1 U8718 ( .B1(n5873), .B2(n5874), .A(n14284), .ZN(n5845) );
  AOI221_X1 U8719 ( .B1(n14411), .B2(n5706), .C1(n14454), .C2(n3322), .A(n5880), .ZN(n5873) );
  AOI221_X1 U8720 ( .B1(n14312), .B2(n5710), .C1(n5893), .C2(n3326), .A(n5877), 
        .ZN(n5874) );
  AOI21_X1 U8721 ( .B1(n5911), .B2(n5912), .A(n5944), .ZN(n5881) );
  AOI221_X1 U8722 ( .B1(n14411), .B2(n5711), .C1(n14454), .C2(n3327), .A(n5918), .ZN(n5911) );
  AOI221_X1 U8723 ( .B1(n14312), .B2(n5713), .C1(n5893), .C2(n3329), .A(n5915), 
        .ZN(n5912) );
  AOI21_X1 U8724 ( .B1(n5947), .B2(n5948), .A(n5916), .ZN(n5919) );
  AOI221_X1 U8725 ( .B1(n14411), .B2(n5714), .C1(n14454), .C2(n3330), .A(n5958), .ZN(n5947) );
  AOI221_X1 U8726 ( .B1(n14312), .B2(n5718), .C1(n5870), .C2(n3334), .A(n5951), 
        .ZN(n5948) );
  AOI21_X1 U8727 ( .B1(n3666), .B2(n3667), .A(n5949), .ZN(n3647) );
  AOI221_X1 U8728 ( .B1(n14429), .B2(n5719), .C1(n14472), .C2(n3335), .A(n3673), .ZN(n3666) );
  AOI221_X1 U8729 ( .B1(n14330), .B2(n5721), .C1(n5897), .C2(n3337), .A(n3670), 
        .ZN(n3667) );
  AOI21_X1 U8730 ( .B1(n5796), .B2(n5797), .A(n5916), .ZN(n5768) );
  AOI221_X1 U8731 ( .B1(n14412), .B2(n5722), .C1(n14455), .C2(n3338), .A(n5803), .ZN(n5796) );
  AOI221_X1 U8732 ( .B1(n14313), .B2(n5726), .C1(n5897), .C2(n3342), .A(n5800), 
        .ZN(n5797) );
  CLKBUF_X1 U8733 ( .A(n239), .Z(n5799) );
  CLKBUF_X1 U8734 ( .A(n239), .Z(n5801) );
  CLKBUF_X1 U8735 ( .A(n239), .Z(n5802) );
  CLKBUF_X1 U8736 ( .A(n239), .Z(n5815) );
  CLKBUF_X1 U8737 ( .A(n239), .Z(n5816) );
  CLKBUF_X1 U8738 ( .A(n239), .Z(n5818) );
  CLKBUF_X1 U8739 ( .A(n239), .Z(n5819) );
  CLKBUF_X1 U8740 ( .A(n239), .Z(n5823) );
  CLKBUF_X1 U8741 ( .A(n239), .Z(n5824) );
  CLKBUF_X1 U8742 ( .A(n239), .Z(n5826) );
  CLKBUF_X1 U8743 ( .A(n239), .Z(n5827) );
  CLKBUF_X1 U8744 ( .A(n239), .Z(n5831) );
  CLKBUF_X1 U8745 ( .A(n239), .Z(n5832) );
  CLKBUF_X1 U8746 ( .A(n239), .Z(n5834) );
  CLKBUF_X1 U8747 ( .A(n239), .Z(n5835) );
  CLKBUF_X1 U8748 ( .A(n239), .Z(n5839) );
  CLKBUF_X1 U8749 ( .A(n239), .Z(n5840) );
  CLKBUF_X1 U8750 ( .A(n239), .Z(n5842) );
  CLKBUF_X1 U8751 ( .A(n239), .Z(n5843) );
  CLKBUF_X1 U8752 ( .A(n239), .Z(n5851) );
  CLKBUF_X1 U8753 ( .A(n239), .Z(n5852) );
  CLKBUF_X1 U8754 ( .A(n239), .Z(n5854) );
  CLKBUF_X1 U8755 ( .A(n239), .Z(n5855) );
  CLKBUF_X1 U8756 ( .A(n239), .Z(n5859) );
  CLKBUF_X1 U8757 ( .A(n239), .Z(n5860) );
  CLKBUF_X1 U8758 ( .A(n239), .Z(n5862) );
  CLKBUF_X1 U8759 ( .A(n239), .Z(n5863) );
  CLKBUF_X1 U8760 ( .A(n239), .Z(n5867) );
  CLKBUF_X1 U8761 ( .A(n239), .Z(n5868) );
  CLKBUF_X1 U8762 ( .A(n239), .Z(n5870) );
  CLKBUF_X1 U8763 ( .A(n239), .Z(n5871) );
  CLKBUF_X1 U8764 ( .A(n239), .Z(n5875) );
  CLKBUF_X1 U8765 ( .A(n239), .Z(n5876) );
  CLKBUF_X1 U8766 ( .A(n239), .Z(n5878) );
  CLKBUF_X1 U8767 ( .A(n239), .Z(n5879) );
  CLKBUF_X1 U8768 ( .A(n239), .Z(n5889) );
  CLKBUF_X1 U8769 ( .A(n239), .Z(n5890) );
  CLKBUF_X1 U8770 ( .A(n239), .Z(n5892) );
  CLKBUF_X1 U8771 ( .A(n239), .Z(n5893) );
  CLKBUF_X1 U8772 ( .A(n239), .Z(n5897) );
  CLKBUF_X1 U8773 ( .A(n5908), .Z(n14351) );
  CLKBUF_X1 U8774 ( .A(n14360), .Z(n14400) );
  CLKBUF_X1 U8775 ( .A(n5898), .Z(n14450) );
  CLKBUF_X1 U8776 ( .A(n5901), .Z(n14493) );
  CLKBUF_X1 U8777 ( .A(n14508), .Z(n14548) );
  CLKBUF_X1 U8778 ( .A(n5905), .Z(n14592) );
  CLKBUF_X1 U8779 ( .A(n5906), .Z(n14645) );
  CLKBUF_X1 U8780 ( .A(n75), .Z(n14689) );
  CLKBUF_X1 U8781 ( .A(n74), .Z(n14729) );
  CLKBUF_X1 U8782 ( .A(n73), .Z(n14769) );
  CLKBUF_X1 U8783 ( .A(n72), .Z(n14809) );
  CLKBUF_X1 U8784 ( .A(n71), .Z(n14849) );
  CLKBUF_X1 U8785 ( .A(n70), .Z(n14889) );
  CLKBUF_X1 U8786 ( .A(n69), .Z(n14929) );
  CLKBUF_X1 U8787 ( .A(n68), .Z(n14969) );
  INV_X1 U8788 ( .A(ADDR[2]), .ZN(n14988) );
endmodule


module CAM_TAG_BIT23_SET_BIT4 ( TAG_IN, TAG_OUT, SET_INDEX, COUNT, VALID, CLK, 
        RST, WE );
  input [22:0] TAG_IN;
  output [22:0] TAG_OUT;
  input [3:0] SET_INDEX;
  input [4:0] COUNT;
  input CLK, RST, WE;
  output VALID;
  wire   \CAM_MEM[15][22] , \CAM_MEM[15][21] , \CAM_MEM[15][20] ,
         \CAM_MEM[15][19] , \CAM_MEM[15][18] , \CAM_MEM[15][17] ,
         \CAM_MEM[15][16] , \CAM_MEM[15][15] , \CAM_MEM[15][14] ,
         \CAM_MEM[15][13] , \CAM_MEM[15][12] , \CAM_MEM[15][11] ,
         \CAM_MEM[15][10] , \CAM_MEM[15][9] , \CAM_MEM[15][8] ,
         \CAM_MEM[15][7] , \CAM_MEM[15][6] , \CAM_MEM[15][5] ,
         \CAM_MEM[15][4] , \CAM_MEM[15][3] , \CAM_MEM[15][2] ,
         \CAM_MEM[15][1] , \CAM_MEM[15][0] , \CAM_MEM[14][22] ,
         \CAM_MEM[14][21] , \CAM_MEM[14][20] , \CAM_MEM[14][19] ,
         \CAM_MEM[14][18] , \CAM_MEM[14][17] , \CAM_MEM[14][16] ,
         \CAM_MEM[14][15] , \CAM_MEM[14][14] , \CAM_MEM[14][13] ,
         \CAM_MEM[14][12] , \CAM_MEM[14][11] , \CAM_MEM[14][10] ,
         \CAM_MEM[14][9] , \CAM_MEM[14][8] , \CAM_MEM[14][7] ,
         \CAM_MEM[14][6] , \CAM_MEM[14][5] , \CAM_MEM[14][4] ,
         \CAM_MEM[14][3] , \CAM_MEM[14][2] , \CAM_MEM[14][1] ,
         \CAM_MEM[14][0] , \CAM_MEM[13][22] , \CAM_MEM[13][21] ,
         \CAM_MEM[13][20] , \CAM_MEM[13][19] , \CAM_MEM[13][18] ,
         \CAM_MEM[13][17] , \CAM_MEM[13][16] , \CAM_MEM[13][15] ,
         \CAM_MEM[13][14] , \CAM_MEM[13][13] , \CAM_MEM[13][12] ,
         \CAM_MEM[13][11] , \CAM_MEM[13][10] , \CAM_MEM[13][9] ,
         \CAM_MEM[13][8] , \CAM_MEM[13][7] , \CAM_MEM[13][6] ,
         \CAM_MEM[13][5] , \CAM_MEM[13][4] , \CAM_MEM[13][3] ,
         \CAM_MEM[13][2] , \CAM_MEM[13][1] , \CAM_MEM[13][0] ,
         \CAM_MEM[12][22] , \CAM_MEM[12][21] , \CAM_MEM[12][20] ,
         \CAM_MEM[12][19] , \CAM_MEM[12][18] , \CAM_MEM[12][17] ,
         \CAM_MEM[12][16] , \CAM_MEM[12][15] , \CAM_MEM[12][14] ,
         \CAM_MEM[12][13] , \CAM_MEM[12][12] , \CAM_MEM[12][11] ,
         \CAM_MEM[12][10] , \CAM_MEM[12][9] , \CAM_MEM[12][8] ,
         \CAM_MEM[12][7] , \CAM_MEM[12][6] , \CAM_MEM[12][5] ,
         \CAM_MEM[12][4] , \CAM_MEM[12][3] , \CAM_MEM[12][2] ,
         \CAM_MEM[12][1] , \CAM_MEM[12][0] , \CAM_MEM[11][22] ,
         \CAM_MEM[11][21] , \CAM_MEM[11][20] , \CAM_MEM[11][19] ,
         \CAM_MEM[11][18] , \CAM_MEM[11][17] , \CAM_MEM[11][16] ,
         \CAM_MEM[11][15] , \CAM_MEM[11][14] , \CAM_MEM[11][13] ,
         \CAM_MEM[11][12] , \CAM_MEM[11][11] , \CAM_MEM[11][10] ,
         \CAM_MEM[11][9] , \CAM_MEM[11][8] , \CAM_MEM[11][7] ,
         \CAM_MEM[11][6] , \CAM_MEM[11][5] , \CAM_MEM[11][4] ,
         \CAM_MEM[11][3] , \CAM_MEM[11][2] , \CAM_MEM[11][1] ,
         \CAM_MEM[11][0] , \CAM_MEM[10][22] , \CAM_MEM[10][21] ,
         \CAM_MEM[10][20] , \CAM_MEM[10][19] , \CAM_MEM[10][18] ,
         \CAM_MEM[10][17] , \CAM_MEM[10][16] , \CAM_MEM[10][15] ,
         \CAM_MEM[10][14] , \CAM_MEM[10][13] , \CAM_MEM[10][12] ,
         \CAM_MEM[10][11] , \CAM_MEM[10][10] , \CAM_MEM[10][9] ,
         \CAM_MEM[10][8] , \CAM_MEM[10][7] , \CAM_MEM[10][6] ,
         \CAM_MEM[10][5] , \CAM_MEM[10][4] , \CAM_MEM[10][3] ,
         \CAM_MEM[10][2] , \CAM_MEM[10][1] , \CAM_MEM[10][0] ,
         \CAM_MEM[9][22] , \CAM_MEM[9][21] , \CAM_MEM[9][20] ,
         \CAM_MEM[9][19] , \CAM_MEM[9][18] , \CAM_MEM[9][17] ,
         \CAM_MEM[9][16] , \CAM_MEM[9][15] , \CAM_MEM[9][14] ,
         \CAM_MEM[9][13] , \CAM_MEM[9][12] , \CAM_MEM[9][11] ,
         \CAM_MEM[9][10] , \CAM_MEM[9][9] , \CAM_MEM[9][8] , \CAM_MEM[9][7] ,
         \CAM_MEM[9][6] , \CAM_MEM[9][5] , \CAM_MEM[9][4] , \CAM_MEM[9][3] ,
         \CAM_MEM[9][2] , \CAM_MEM[9][1] , \CAM_MEM[9][0] , \CAM_MEM[8][22] ,
         \CAM_MEM[8][21] , \CAM_MEM[8][20] , \CAM_MEM[8][19] ,
         \CAM_MEM[8][18] , \CAM_MEM[8][17] , \CAM_MEM[8][16] ,
         \CAM_MEM[8][15] , \CAM_MEM[8][14] , \CAM_MEM[8][13] ,
         \CAM_MEM[8][12] , \CAM_MEM[8][11] , \CAM_MEM[8][10] , \CAM_MEM[8][9] ,
         \CAM_MEM[8][8] , \CAM_MEM[8][7] , \CAM_MEM[8][6] , \CAM_MEM[8][5] ,
         \CAM_MEM[8][4] , \CAM_MEM[8][3] , \CAM_MEM[8][2] , \CAM_MEM[8][1] ,
         \CAM_MEM[8][0] , \CAM_MEM[7][22] , \CAM_MEM[7][21] , \CAM_MEM[7][20] ,
         \CAM_MEM[7][19] , \CAM_MEM[7][18] , \CAM_MEM[7][17] ,
         \CAM_MEM[7][16] , \CAM_MEM[7][15] , \CAM_MEM[7][14] ,
         \CAM_MEM[7][13] , \CAM_MEM[7][12] , \CAM_MEM[7][11] ,
         \CAM_MEM[7][10] , \CAM_MEM[7][9] , \CAM_MEM[7][8] , \CAM_MEM[7][7] ,
         \CAM_MEM[7][6] , \CAM_MEM[7][5] , \CAM_MEM[7][4] , \CAM_MEM[7][3] ,
         \CAM_MEM[7][2] , \CAM_MEM[7][1] , \CAM_MEM[7][0] , \CAM_MEM[6][22] ,
         \CAM_MEM[6][21] , \CAM_MEM[6][20] , \CAM_MEM[6][19] ,
         \CAM_MEM[6][18] , \CAM_MEM[6][17] , \CAM_MEM[6][16] ,
         \CAM_MEM[6][15] , \CAM_MEM[6][14] , \CAM_MEM[6][13] ,
         \CAM_MEM[6][12] , \CAM_MEM[6][11] , \CAM_MEM[6][10] , \CAM_MEM[6][9] ,
         \CAM_MEM[6][8] , \CAM_MEM[6][7] , \CAM_MEM[6][6] , \CAM_MEM[6][5] ,
         \CAM_MEM[6][4] , \CAM_MEM[6][3] , \CAM_MEM[6][2] , \CAM_MEM[6][1] ,
         \CAM_MEM[6][0] , \CAM_MEM[5][22] , \CAM_MEM[5][21] , \CAM_MEM[5][20] ,
         \CAM_MEM[5][19] , \CAM_MEM[5][18] , \CAM_MEM[5][17] ,
         \CAM_MEM[5][16] , \CAM_MEM[5][15] , \CAM_MEM[5][14] ,
         \CAM_MEM[5][13] , \CAM_MEM[5][12] , \CAM_MEM[5][11] ,
         \CAM_MEM[5][10] , \CAM_MEM[5][9] , \CAM_MEM[5][8] , \CAM_MEM[5][7] ,
         \CAM_MEM[5][6] , \CAM_MEM[5][5] , \CAM_MEM[5][4] , \CAM_MEM[5][3] ,
         \CAM_MEM[5][2] , \CAM_MEM[5][1] , \CAM_MEM[5][0] , \CAM_MEM[4][22] ,
         \CAM_MEM[4][21] , \CAM_MEM[4][20] , \CAM_MEM[4][19] ,
         \CAM_MEM[4][18] , \CAM_MEM[4][17] , \CAM_MEM[4][16] ,
         \CAM_MEM[4][15] , \CAM_MEM[4][14] , \CAM_MEM[4][13] ,
         \CAM_MEM[4][12] , \CAM_MEM[4][11] , \CAM_MEM[4][10] , \CAM_MEM[4][9] ,
         \CAM_MEM[4][8] , \CAM_MEM[4][7] , \CAM_MEM[4][6] , \CAM_MEM[4][5] ,
         \CAM_MEM[4][4] , \CAM_MEM[4][3] , \CAM_MEM[4][2] , \CAM_MEM[4][1] ,
         \CAM_MEM[4][0] , \CAM_MEM[3][22] , \CAM_MEM[3][21] , \CAM_MEM[3][20] ,
         \CAM_MEM[3][19] , \CAM_MEM[3][18] , \CAM_MEM[3][17] ,
         \CAM_MEM[3][16] , \CAM_MEM[3][15] , \CAM_MEM[3][14] ,
         \CAM_MEM[3][13] , \CAM_MEM[3][12] , \CAM_MEM[3][11] ,
         \CAM_MEM[3][10] , \CAM_MEM[3][9] , \CAM_MEM[3][8] , \CAM_MEM[3][7] ,
         \CAM_MEM[3][6] , \CAM_MEM[3][5] , \CAM_MEM[3][4] , \CAM_MEM[3][3] ,
         \CAM_MEM[3][2] , \CAM_MEM[3][1] , \CAM_MEM[3][0] , \CAM_MEM[2][22] ,
         \CAM_MEM[2][21] , \CAM_MEM[2][20] , \CAM_MEM[2][19] ,
         \CAM_MEM[2][18] , \CAM_MEM[2][17] , \CAM_MEM[2][16] ,
         \CAM_MEM[2][15] , \CAM_MEM[2][14] , \CAM_MEM[2][13] ,
         \CAM_MEM[2][12] , \CAM_MEM[2][11] , \CAM_MEM[2][10] , \CAM_MEM[2][9] ,
         \CAM_MEM[2][8] , \CAM_MEM[2][7] , \CAM_MEM[2][6] , \CAM_MEM[2][5] ,
         \CAM_MEM[2][4] , \CAM_MEM[2][3] , \CAM_MEM[2][2] , \CAM_MEM[2][1] ,
         \CAM_MEM[2][0] , \CAM_MEM[1][22] , \CAM_MEM[1][21] , \CAM_MEM[1][20] ,
         \CAM_MEM[1][19] , \CAM_MEM[1][18] , \CAM_MEM[1][17] ,
         \CAM_MEM[1][16] , \CAM_MEM[1][15] , \CAM_MEM[1][14] ,
         \CAM_MEM[1][13] , \CAM_MEM[1][12] , \CAM_MEM[1][11] ,
         \CAM_MEM[1][10] , \CAM_MEM[1][9] , \CAM_MEM[1][8] , \CAM_MEM[1][7] ,
         \CAM_MEM[1][6] , \CAM_MEM[1][5] , \CAM_MEM[1][4] , \CAM_MEM[1][3] ,
         \CAM_MEM[1][2] , \CAM_MEM[1][1] , \CAM_MEM[1][0] , \CAM_MEM[0][22] ,
         \CAM_MEM[0][21] , \CAM_MEM[0][20] , \CAM_MEM[0][19] ,
         \CAM_MEM[0][18] , \CAM_MEM[0][17] , \CAM_MEM[0][16] ,
         \CAM_MEM[0][15] , \CAM_MEM[0][14] , \CAM_MEM[0][13] ,
         \CAM_MEM[0][12] , \CAM_MEM[0][11] , \CAM_MEM[0][10] , \CAM_MEM[0][9] ,
         \CAM_MEM[0][8] , \CAM_MEM[0][7] , \CAM_MEM[0][6] , \CAM_MEM[0][5] ,
         \CAM_MEM[0][4] , \CAM_MEM[0][3] , \CAM_MEM[0][2] , \CAM_MEM[0][1] ,
         \CAM_MEM[0][0] , N221, N606, N607, N608, N609, N610, N611, N612, N613,
         N614, N615, N616, N617, N618, N619, N620, N621, N622, N623, N624,
         N625, N626, N627, N628, N631, N632, N633, N634, N635, N636, N637,
         N638, N639, N640, N641, N642, N643, N644, N645, N646, N671, N694,
         N717, N740, N763, N786, N809, N832, N855, N878, N901, N924, N947,
         N970, N993, N999, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n14, n15,
         n16, n17, n18, n19, n20, n21, n24, n25, n26, n27, n28, n29, n30, n31,
         n1, n12, n13, n22, n23, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399;
  wire   [15:0] VALID_BIT;

  DLL_X1 \TAG_OUT_reg[22]  ( .D(N628), .GN(n396), .Q(TAG_OUT[22]) );
  DLL_X1 \TAG_OUT_reg[21]  ( .D(N627), .GN(n398), .Q(TAG_OUT[21]) );
  DLL_X1 \TAG_OUT_reg[20]  ( .D(N626), .GN(n398), .Q(TAG_OUT[20]) );
  DLL_X1 \TAG_OUT_reg[19]  ( .D(N625), .GN(n398), .Q(TAG_OUT[19]) );
  DLL_X1 \TAG_OUT_reg[18]  ( .D(N624), .GN(n397), .Q(TAG_OUT[18]) );
  DLL_X1 \TAG_OUT_reg[17]  ( .D(N623), .GN(n397), .Q(TAG_OUT[17]) );
  DLL_X1 \TAG_OUT_reg[16]  ( .D(N622), .GN(n397), .Q(TAG_OUT[16]) );
  DLL_X1 \TAG_OUT_reg[15]  ( .D(N621), .GN(n397), .Q(TAG_OUT[15]) );
  DLL_X1 \TAG_OUT_reg[14]  ( .D(N620), .GN(n397), .Q(TAG_OUT[14]) );
  DLL_X1 \TAG_OUT_reg[13]  ( .D(N619), .GN(n397), .Q(TAG_OUT[13]) );
  DLL_X1 \TAG_OUT_reg[12]  ( .D(N618), .GN(n397), .Q(TAG_OUT[12]) );
  DLL_X1 \TAG_OUT_reg[11]  ( .D(N617), .GN(n397), .Q(TAG_OUT[11]) );
  DLL_X1 \TAG_OUT_reg[10]  ( .D(N616), .GN(n397), .Q(TAG_OUT[10]) );
  DLL_X1 \TAG_OUT_reg[9]  ( .D(N615), .GN(n397), .Q(TAG_OUT[9]) );
  DLL_X1 \TAG_OUT_reg[8]  ( .D(N614), .GN(n397), .Q(TAG_OUT[8]) );
  DLL_X1 \TAG_OUT_reg[7]  ( .D(N613), .GN(n397), .Q(TAG_OUT[7]) );
  DLL_X1 \TAG_OUT_reg[6]  ( .D(N612), .GN(n396), .Q(TAG_OUT[6]) );
  DLL_X1 \TAG_OUT_reg[5]  ( .D(N611), .GN(n396), .Q(TAG_OUT[5]) );
  DLL_X1 \TAG_OUT_reg[4]  ( .D(N610), .GN(n396), .Q(TAG_OUT[4]) );
  DLL_X1 \TAG_OUT_reg[3]  ( .D(N609), .GN(n397), .Q(TAG_OUT[3]) );
  DLL_X1 \TAG_OUT_reg[2]  ( .D(N608), .GN(n396), .Q(TAG_OUT[2]) );
  DLL_X1 \TAG_OUT_reg[1]  ( .D(N607), .GN(n396), .Q(TAG_OUT[1]) );
  DLL_X1 \TAG_OUT_reg[0]  ( .D(N606), .GN(n396), .Q(TAG_OUT[0]) );
  DLH_X1 \VALID_BIT_reg[15]  ( .G(N646), .D(n399), .Q(VALID_BIT[15]) );
  DLH_X1 \VALID_BIT_reg[14]  ( .G(N645), .D(n399), .Q(VALID_BIT[14]) );
  DLH_X1 \VALID_BIT_reg[13]  ( .G(N644), .D(n399), .Q(VALID_BIT[13]) );
  DLH_X1 \VALID_BIT_reg[12]  ( .G(N643), .D(n399), .Q(VALID_BIT[12]) );
  DLH_X1 \VALID_BIT_reg[11]  ( .G(N642), .D(n399), .Q(VALID_BIT[11]) );
  DLH_X1 \VALID_BIT_reg[10]  ( .G(N641), .D(n399), .Q(VALID_BIT[10]) );
  DLH_X1 \VALID_BIT_reg[9]  ( .G(N640), .D(n399), .Q(VALID_BIT[9]) );
  DLH_X1 \VALID_BIT_reg[8]  ( .G(N639), .D(n399), .Q(VALID_BIT[8]) );
  DLH_X1 \VALID_BIT_reg[7]  ( .G(N638), .D(n399), .Q(VALID_BIT[7]) );
  DLH_X1 \VALID_BIT_reg[6]  ( .G(N637), .D(n399), .Q(VALID_BIT[6]) );
  DLH_X1 \VALID_BIT_reg[5]  ( .G(N636), .D(n399), .Q(VALID_BIT[5]) );
  DLH_X1 \VALID_BIT_reg[4]  ( .G(N635), .D(n399), .Q(VALID_BIT[4]) );
  DLH_X1 \VALID_BIT_reg[3]  ( .G(N634), .D(n399), .Q(VALID_BIT[3]) );
  DLH_X1 \VALID_BIT_reg[2]  ( .G(N633), .D(n399), .Q(VALID_BIT[2]) );
  DLH_X1 \VALID_BIT_reg[1]  ( .G(N632), .D(n399), .Q(VALID_BIT[1]) );
  DLH_X1 \VALID_BIT_reg[0]  ( .G(N631), .D(n399), .Q(VALID_BIT[0]) );
  DLH_X1 \CAM_MEM_reg[15][22]  ( .G(N999), .D(TAG_IN[22]), .Q(
        \CAM_MEM[15][22] ) );
  DLH_X1 \CAM_MEM_reg[15][21]  ( .G(N999), .D(TAG_IN[21]), .Q(
        \CAM_MEM[15][21] ) );
  DLH_X1 \CAM_MEM_reg[15][20]  ( .G(N999), .D(TAG_IN[20]), .Q(
        \CAM_MEM[15][20] ) );
  DLH_X1 \CAM_MEM_reg[15][19]  ( .G(N999), .D(TAG_IN[19]), .Q(
        \CAM_MEM[15][19] ) );
  DLH_X1 \CAM_MEM_reg[15][18]  ( .G(N999), .D(TAG_IN[18]), .Q(
        \CAM_MEM[15][18] ) );
  DLH_X1 \CAM_MEM_reg[15][17]  ( .G(N999), .D(TAG_IN[17]), .Q(
        \CAM_MEM[15][17] ) );
  DLH_X1 \CAM_MEM_reg[15][16]  ( .G(N999), .D(TAG_IN[16]), .Q(
        \CAM_MEM[15][16] ) );
  DLH_X1 \CAM_MEM_reg[15][15]  ( .G(N999), .D(TAG_IN[15]), .Q(
        \CAM_MEM[15][15] ) );
  DLH_X1 \CAM_MEM_reg[15][14]  ( .G(N999), .D(TAG_IN[14]), .Q(
        \CAM_MEM[15][14] ) );
  DLH_X1 \CAM_MEM_reg[15][13]  ( .G(N999), .D(TAG_IN[13]), .Q(
        \CAM_MEM[15][13] ) );
  DLH_X1 \CAM_MEM_reg[15][12]  ( .G(N999), .D(TAG_IN[12]), .Q(
        \CAM_MEM[15][12] ) );
  DLH_X1 \CAM_MEM_reg[15][11]  ( .G(N999), .D(TAG_IN[11]), .Q(
        \CAM_MEM[15][11] ) );
  DLH_X1 \CAM_MEM_reg[15][10]  ( .G(N999), .D(TAG_IN[10]), .Q(
        \CAM_MEM[15][10] ) );
  DLH_X1 \CAM_MEM_reg[15][9]  ( .G(N999), .D(TAG_IN[9]), .Q(\CAM_MEM[15][9] )
         );
  DLH_X1 \CAM_MEM_reg[15][8]  ( .G(N999), .D(TAG_IN[8]), .Q(\CAM_MEM[15][8] )
         );
  DLH_X1 \CAM_MEM_reg[15][7]  ( .G(N999), .D(TAG_IN[7]), .Q(\CAM_MEM[15][7] )
         );
  DLH_X1 \CAM_MEM_reg[15][6]  ( .G(N999), .D(TAG_IN[6]), .Q(\CAM_MEM[15][6] )
         );
  DLH_X1 \CAM_MEM_reg[15][5]  ( .G(N999), .D(TAG_IN[5]), .Q(\CAM_MEM[15][5] )
         );
  DLH_X1 \CAM_MEM_reg[15][4]  ( .G(N999), .D(TAG_IN[4]), .Q(\CAM_MEM[15][4] )
         );
  DLH_X1 \CAM_MEM_reg[15][3]  ( .G(N999), .D(TAG_IN[3]), .Q(\CAM_MEM[15][3] )
         );
  DLH_X1 \CAM_MEM_reg[15][2]  ( .G(N999), .D(TAG_IN[2]), .Q(\CAM_MEM[15][2] )
         );
  DLH_X1 \CAM_MEM_reg[15][1]  ( .G(N999), .D(TAG_IN[1]), .Q(\CAM_MEM[15][1] )
         );
  DLH_X1 \CAM_MEM_reg[15][0]  ( .G(N999), .D(TAG_IN[0]), .Q(\CAM_MEM[15][0] )
         );
  DLH_X1 \CAM_MEM_reg[14][22]  ( .G(N993), .D(TAG_IN[22]), .Q(
        \CAM_MEM[14][22] ) );
  DLH_X1 \CAM_MEM_reg[14][21]  ( .G(N993), .D(TAG_IN[21]), .Q(
        \CAM_MEM[14][21] ) );
  DLH_X1 \CAM_MEM_reg[14][20]  ( .G(N993), .D(TAG_IN[20]), .Q(
        \CAM_MEM[14][20] ) );
  DLH_X1 \CAM_MEM_reg[14][19]  ( .G(N993), .D(TAG_IN[19]), .Q(
        \CAM_MEM[14][19] ) );
  DLH_X1 \CAM_MEM_reg[14][18]  ( .G(N993), .D(TAG_IN[18]), .Q(
        \CAM_MEM[14][18] ) );
  DLH_X1 \CAM_MEM_reg[14][17]  ( .G(N993), .D(TAG_IN[17]), .Q(
        \CAM_MEM[14][17] ) );
  DLH_X1 \CAM_MEM_reg[14][16]  ( .G(N993), .D(TAG_IN[16]), .Q(
        \CAM_MEM[14][16] ) );
  DLH_X1 \CAM_MEM_reg[14][15]  ( .G(N993), .D(TAG_IN[15]), .Q(
        \CAM_MEM[14][15] ) );
  DLH_X1 \CAM_MEM_reg[14][14]  ( .G(N993), .D(TAG_IN[14]), .Q(
        \CAM_MEM[14][14] ) );
  DLH_X1 \CAM_MEM_reg[14][13]  ( .G(N993), .D(TAG_IN[13]), .Q(
        \CAM_MEM[14][13] ) );
  DLH_X1 \CAM_MEM_reg[14][12]  ( .G(N993), .D(TAG_IN[12]), .Q(
        \CAM_MEM[14][12] ) );
  DLH_X1 \CAM_MEM_reg[14][11]  ( .G(N993), .D(TAG_IN[11]), .Q(
        \CAM_MEM[14][11] ) );
  DLH_X1 \CAM_MEM_reg[14][10]  ( .G(N993), .D(TAG_IN[10]), .Q(
        \CAM_MEM[14][10] ) );
  DLH_X1 \CAM_MEM_reg[14][9]  ( .G(N993), .D(TAG_IN[9]), .Q(\CAM_MEM[14][9] )
         );
  DLH_X1 \CAM_MEM_reg[14][8]  ( .G(N993), .D(TAG_IN[8]), .Q(\CAM_MEM[14][8] )
         );
  DLH_X1 \CAM_MEM_reg[14][7]  ( .G(N993), .D(TAG_IN[7]), .Q(\CAM_MEM[14][7] )
         );
  DLH_X1 \CAM_MEM_reg[14][6]  ( .G(N993), .D(TAG_IN[6]), .Q(\CAM_MEM[14][6] )
         );
  DLH_X1 \CAM_MEM_reg[14][5]  ( .G(N993), .D(TAG_IN[5]), .Q(\CAM_MEM[14][5] )
         );
  DLH_X1 \CAM_MEM_reg[14][4]  ( .G(N993), .D(TAG_IN[4]), .Q(\CAM_MEM[14][4] )
         );
  DLH_X1 \CAM_MEM_reg[14][3]  ( .G(N993), .D(TAG_IN[3]), .Q(\CAM_MEM[14][3] )
         );
  DLH_X1 \CAM_MEM_reg[14][2]  ( .G(N993), .D(TAG_IN[2]), .Q(\CAM_MEM[14][2] )
         );
  DLH_X1 \CAM_MEM_reg[14][1]  ( .G(N993), .D(TAG_IN[1]), .Q(\CAM_MEM[14][1] )
         );
  DLH_X1 \CAM_MEM_reg[14][0]  ( .G(N993), .D(TAG_IN[0]), .Q(\CAM_MEM[14][0] )
         );
  DLH_X1 \CAM_MEM_reg[13][22]  ( .G(N970), .D(TAG_IN[22]), .Q(
        \CAM_MEM[13][22] ) );
  DLH_X1 \CAM_MEM_reg[13][21]  ( .G(N970), .D(TAG_IN[21]), .Q(
        \CAM_MEM[13][21] ) );
  DLH_X1 \CAM_MEM_reg[13][20]  ( .G(N970), .D(TAG_IN[20]), .Q(
        \CAM_MEM[13][20] ) );
  DLH_X1 \CAM_MEM_reg[13][19]  ( .G(N970), .D(TAG_IN[19]), .Q(
        \CAM_MEM[13][19] ) );
  DLH_X1 \CAM_MEM_reg[13][18]  ( .G(N970), .D(TAG_IN[18]), .Q(
        \CAM_MEM[13][18] ) );
  DLH_X1 \CAM_MEM_reg[13][17]  ( .G(N970), .D(TAG_IN[17]), .Q(
        \CAM_MEM[13][17] ) );
  DLH_X1 \CAM_MEM_reg[13][16]  ( .G(N970), .D(TAG_IN[16]), .Q(
        \CAM_MEM[13][16] ) );
  DLH_X1 \CAM_MEM_reg[13][15]  ( .G(N970), .D(TAG_IN[15]), .Q(
        \CAM_MEM[13][15] ) );
  DLH_X1 \CAM_MEM_reg[13][14]  ( .G(N970), .D(TAG_IN[14]), .Q(
        \CAM_MEM[13][14] ) );
  DLH_X1 \CAM_MEM_reg[13][13]  ( .G(N970), .D(TAG_IN[13]), .Q(
        \CAM_MEM[13][13] ) );
  DLH_X1 \CAM_MEM_reg[13][12]  ( .G(N970), .D(TAG_IN[12]), .Q(
        \CAM_MEM[13][12] ) );
  DLH_X1 \CAM_MEM_reg[13][11]  ( .G(N970), .D(TAG_IN[11]), .Q(
        \CAM_MEM[13][11] ) );
  DLH_X1 \CAM_MEM_reg[13][10]  ( .G(N970), .D(TAG_IN[10]), .Q(
        \CAM_MEM[13][10] ) );
  DLH_X1 \CAM_MEM_reg[13][9]  ( .G(N970), .D(TAG_IN[9]), .Q(\CAM_MEM[13][9] )
         );
  DLH_X1 \CAM_MEM_reg[13][8]  ( .G(N970), .D(TAG_IN[8]), .Q(\CAM_MEM[13][8] )
         );
  DLH_X1 \CAM_MEM_reg[13][7]  ( .G(N970), .D(TAG_IN[7]), .Q(\CAM_MEM[13][7] )
         );
  DLH_X1 \CAM_MEM_reg[13][6]  ( .G(N970), .D(TAG_IN[6]), .Q(\CAM_MEM[13][6] )
         );
  DLH_X1 \CAM_MEM_reg[13][5]  ( .G(N970), .D(TAG_IN[5]), .Q(\CAM_MEM[13][5] )
         );
  DLH_X1 \CAM_MEM_reg[13][4]  ( .G(N970), .D(TAG_IN[4]), .Q(\CAM_MEM[13][4] )
         );
  DLH_X1 \CAM_MEM_reg[13][3]  ( .G(N970), .D(TAG_IN[3]), .Q(\CAM_MEM[13][3] )
         );
  DLH_X1 \CAM_MEM_reg[13][2]  ( .G(N970), .D(TAG_IN[2]), .Q(\CAM_MEM[13][2] )
         );
  DLH_X1 \CAM_MEM_reg[13][1]  ( .G(N970), .D(TAG_IN[1]), .Q(\CAM_MEM[13][1] )
         );
  DLH_X1 \CAM_MEM_reg[13][0]  ( .G(N970), .D(TAG_IN[0]), .Q(\CAM_MEM[13][0] )
         );
  DLH_X1 \CAM_MEM_reg[12][22]  ( .G(N947), .D(TAG_IN[22]), .Q(
        \CAM_MEM[12][22] ) );
  DLH_X1 \CAM_MEM_reg[12][21]  ( .G(N947), .D(TAG_IN[21]), .Q(
        \CAM_MEM[12][21] ) );
  DLH_X1 \CAM_MEM_reg[12][20]  ( .G(N947), .D(TAG_IN[20]), .Q(
        \CAM_MEM[12][20] ) );
  DLH_X1 \CAM_MEM_reg[12][19]  ( .G(N947), .D(TAG_IN[19]), .Q(
        \CAM_MEM[12][19] ) );
  DLH_X1 \CAM_MEM_reg[12][18]  ( .G(N947), .D(TAG_IN[18]), .Q(
        \CAM_MEM[12][18] ) );
  DLH_X1 \CAM_MEM_reg[12][17]  ( .G(N947), .D(TAG_IN[17]), .Q(
        \CAM_MEM[12][17] ) );
  DLH_X1 \CAM_MEM_reg[12][16]  ( .G(N947), .D(TAG_IN[16]), .Q(
        \CAM_MEM[12][16] ) );
  DLH_X1 \CAM_MEM_reg[12][15]  ( .G(N947), .D(TAG_IN[15]), .Q(
        \CAM_MEM[12][15] ) );
  DLH_X1 \CAM_MEM_reg[12][14]  ( .G(N947), .D(TAG_IN[14]), .Q(
        \CAM_MEM[12][14] ) );
  DLH_X1 \CAM_MEM_reg[12][13]  ( .G(N947), .D(TAG_IN[13]), .Q(
        \CAM_MEM[12][13] ) );
  DLH_X1 \CAM_MEM_reg[12][12]  ( .G(N947), .D(TAG_IN[12]), .Q(
        \CAM_MEM[12][12] ) );
  DLH_X1 \CAM_MEM_reg[12][11]  ( .G(N947), .D(TAG_IN[11]), .Q(
        \CAM_MEM[12][11] ) );
  DLH_X1 \CAM_MEM_reg[12][10]  ( .G(N947), .D(TAG_IN[10]), .Q(
        \CAM_MEM[12][10] ) );
  DLH_X1 \CAM_MEM_reg[12][9]  ( .G(N947), .D(TAG_IN[9]), .Q(\CAM_MEM[12][9] )
         );
  DLH_X1 \CAM_MEM_reg[12][8]  ( .G(N947), .D(TAG_IN[8]), .Q(\CAM_MEM[12][8] )
         );
  DLH_X1 \CAM_MEM_reg[12][7]  ( .G(N947), .D(TAG_IN[7]), .Q(\CAM_MEM[12][7] )
         );
  DLH_X1 \CAM_MEM_reg[12][6]  ( .G(N947), .D(TAG_IN[6]), .Q(\CAM_MEM[12][6] )
         );
  DLH_X1 \CAM_MEM_reg[12][5]  ( .G(N947), .D(TAG_IN[5]), .Q(\CAM_MEM[12][5] )
         );
  DLH_X1 \CAM_MEM_reg[12][4]  ( .G(N947), .D(TAG_IN[4]), .Q(\CAM_MEM[12][4] )
         );
  DLH_X1 \CAM_MEM_reg[12][3]  ( .G(N947), .D(TAG_IN[3]), .Q(\CAM_MEM[12][3] )
         );
  DLH_X1 \CAM_MEM_reg[12][2]  ( .G(N947), .D(TAG_IN[2]), .Q(\CAM_MEM[12][2] )
         );
  DLH_X1 \CAM_MEM_reg[12][1]  ( .G(N947), .D(TAG_IN[1]), .Q(\CAM_MEM[12][1] )
         );
  DLH_X1 \CAM_MEM_reg[12][0]  ( .G(N947), .D(TAG_IN[0]), .Q(\CAM_MEM[12][0] )
         );
  DLH_X1 \CAM_MEM_reg[11][22]  ( .G(N924), .D(TAG_IN[22]), .Q(
        \CAM_MEM[11][22] ) );
  DLH_X1 \CAM_MEM_reg[11][21]  ( .G(N924), .D(TAG_IN[21]), .Q(
        \CAM_MEM[11][21] ) );
  DLH_X1 \CAM_MEM_reg[11][20]  ( .G(N924), .D(TAG_IN[20]), .Q(
        \CAM_MEM[11][20] ) );
  DLH_X1 \CAM_MEM_reg[11][19]  ( .G(N924), .D(TAG_IN[19]), .Q(
        \CAM_MEM[11][19] ) );
  DLH_X1 \CAM_MEM_reg[11][18]  ( .G(N924), .D(TAG_IN[18]), .Q(
        \CAM_MEM[11][18] ) );
  DLH_X1 \CAM_MEM_reg[11][17]  ( .G(N924), .D(TAG_IN[17]), .Q(
        \CAM_MEM[11][17] ) );
  DLH_X1 \CAM_MEM_reg[11][16]  ( .G(N924), .D(TAG_IN[16]), .Q(
        \CAM_MEM[11][16] ) );
  DLH_X1 \CAM_MEM_reg[11][15]  ( .G(N924), .D(TAG_IN[15]), .Q(
        \CAM_MEM[11][15] ) );
  DLH_X1 \CAM_MEM_reg[11][14]  ( .G(N924), .D(TAG_IN[14]), .Q(
        \CAM_MEM[11][14] ) );
  DLH_X1 \CAM_MEM_reg[11][13]  ( .G(N924), .D(TAG_IN[13]), .Q(
        \CAM_MEM[11][13] ) );
  DLH_X1 \CAM_MEM_reg[11][12]  ( .G(N924), .D(TAG_IN[12]), .Q(
        \CAM_MEM[11][12] ) );
  DLH_X1 \CAM_MEM_reg[11][11]  ( .G(N924), .D(TAG_IN[11]), .Q(
        \CAM_MEM[11][11] ) );
  DLH_X1 \CAM_MEM_reg[11][10]  ( .G(N924), .D(TAG_IN[10]), .Q(
        \CAM_MEM[11][10] ) );
  DLH_X1 \CAM_MEM_reg[11][9]  ( .G(N924), .D(TAG_IN[9]), .Q(\CAM_MEM[11][9] )
         );
  DLH_X1 \CAM_MEM_reg[11][8]  ( .G(N924), .D(TAG_IN[8]), .Q(\CAM_MEM[11][8] )
         );
  DLH_X1 \CAM_MEM_reg[11][7]  ( .G(N924), .D(TAG_IN[7]), .Q(\CAM_MEM[11][7] )
         );
  DLH_X1 \CAM_MEM_reg[11][6]  ( .G(N924), .D(TAG_IN[6]), .Q(\CAM_MEM[11][6] )
         );
  DLH_X1 \CAM_MEM_reg[11][5]  ( .G(N924), .D(TAG_IN[5]), .Q(\CAM_MEM[11][5] )
         );
  DLH_X1 \CAM_MEM_reg[11][4]  ( .G(N924), .D(TAG_IN[4]), .Q(\CAM_MEM[11][4] )
         );
  DLH_X1 \CAM_MEM_reg[11][3]  ( .G(N924), .D(TAG_IN[3]), .Q(\CAM_MEM[11][3] )
         );
  DLH_X1 \CAM_MEM_reg[11][2]  ( .G(N924), .D(TAG_IN[2]), .Q(\CAM_MEM[11][2] )
         );
  DLH_X1 \CAM_MEM_reg[11][1]  ( .G(N924), .D(TAG_IN[1]), .Q(\CAM_MEM[11][1] )
         );
  DLH_X1 \CAM_MEM_reg[11][0]  ( .G(N924), .D(TAG_IN[0]), .Q(\CAM_MEM[11][0] )
         );
  DLH_X1 \CAM_MEM_reg[10][22]  ( .G(N901), .D(TAG_IN[22]), .Q(
        \CAM_MEM[10][22] ) );
  DLH_X1 \CAM_MEM_reg[10][21]  ( .G(N901), .D(TAG_IN[21]), .Q(
        \CAM_MEM[10][21] ) );
  DLH_X1 \CAM_MEM_reg[10][20]  ( .G(N901), .D(TAG_IN[20]), .Q(
        \CAM_MEM[10][20] ) );
  DLH_X1 \CAM_MEM_reg[10][19]  ( .G(N901), .D(TAG_IN[19]), .Q(
        \CAM_MEM[10][19] ) );
  DLH_X1 \CAM_MEM_reg[10][18]  ( .G(N901), .D(TAG_IN[18]), .Q(
        \CAM_MEM[10][18] ) );
  DLH_X1 \CAM_MEM_reg[10][17]  ( .G(N901), .D(TAG_IN[17]), .Q(
        \CAM_MEM[10][17] ) );
  DLH_X1 \CAM_MEM_reg[10][16]  ( .G(N901), .D(TAG_IN[16]), .Q(
        \CAM_MEM[10][16] ) );
  DLH_X1 \CAM_MEM_reg[10][15]  ( .G(N901), .D(TAG_IN[15]), .Q(
        \CAM_MEM[10][15] ) );
  DLH_X1 \CAM_MEM_reg[10][14]  ( .G(N901), .D(TAG_IN[14]), .Q(
        \CAM_MEM[10][14] ) );
  DLH_X1 \CAM_MEM_reg[10][13]  ( .G(N901), .D(TAG_IN[13]), .Q(
        \CAM_MEM[10][13] ) );
  DLH_X1 \CAM_MEM_reg[10][12]  ( .G(N901), .D(TAG_IN[12]), .Q(
        \CAM_MEM[10][12] ) );
  DLH_X1 \CAM_MEM_reg[10][11]  ( .G(N901), .D(TAG_IN[11]), .Q(
        \CAM_MEM[10][11] ) );
  DLH_X1 \CAM_MEM_reg[10][10]  ( .G(N901), .D(TAG_IN[10]), .Q(
        \CAM_MEM[10][10] ) );
  DLH_X1 \CAM_MEM_reg[10][9]  ( .G(N901), .D(TAG_IN[9]), .Q(\CAM_MEM[10][9] )
         );
  DLH_X1 \CAM_MEM_reg[10][8]  ( .G(N901), .D(TAG_IN[8]), .Q(\CAM_MEM[10][8] )
         );
  DLH_X1 \CAM_MEM_reg[10][7]  ( .G(N901), .D(TAG_IN[7]), .Q(\CAM_MEM[10][7] )
         );
  DLH_X1 \CAM_MEM_reg[10][6]  ( .G(N901), .D(TAG_IN[6]), .Q(\CAM_MEM[10][6] )
         );
  DLH_X1 \CAM_MEM_reg[10][5]  ( .G(N901), .D(TAG_IN[5]), .Q(\CAM_MEM[10][5] )
         );
  DLH_X1 \CAM_MEM_reg[10][4]  ( .G(N901), .D(TAG_IN[4]), .Q(\CAM_MEM[10][4] )
         );
  DLH_X1 \CAM_MEM_reg[10][3]  ( .G(N901), .D(TAG_IN[3]), .Q(\CAM_MEM[10][3] )
         );
  DLH_X1 \CAM_MEM_reg[10][2]  ( .G(N901), .D(TAG_IN[2]), .Q(\CAM_MEM[10][2] )
         );
  DLH_X1 \CAM_MEM_reg[10][1]  ( .G(N901), .D(TAG_IN[1]), .Q(\CAM_MEM[10][1] )
         );
  DLH_X1 \CAM_MEM_reg[10][0]  ( .G(N901), .D(TAG_IN[0]), .Q(\CAM_MEM[10][0] )
         );
  DLH_X1 \CAM_MEM_reg[9][22]  ( .G(N878), .D(TAG_IN[22]), .Q(\CAM_MEM[9][22] )
         );
  DLH_X1 \CAM_MEM_reg[9][21]  ( .G(N878), .D(TAG_IN[21]), .Q(\CAM_MEM[9][21] )
         );
  DLH_X1 \CAM_MEM_reg[9][20]  ( .G(N878), .D(TAG_IN[20]), .Q(\CAM_MEM[9][20] )
         );
  DLH_X1 \CAM_MEM_reg[9][19]  ( .G(N878), .D(TAG_IN[19]), .Q(\CAM_MEM[9][19] )
         );
  DLH_X1 \CAM_MEM_reg[9][18]  ( .G(N878), .D(TAG_IN[18]), .Q(\CAM_MEM[9][18] )
         );
  DLH_X1 \CAM_MEM_reg[9][17]  ( .G(N878), .D(TAG_IN[17]), .Q(\CAM_MEM[9][17] )
         );
  DLH_X1 \CAM_MEM_reg[9][16]  ( .G(N878), .D(TAG_IN[16]), .Q(\CAM_MEM[9][16] )
         );
  DLH_X1 \CAM_MEM_reg[9][15]  ( .G(N878), .D(TAG_IN[15]), .Q(\CAM_MEM[9][15] )
         );
  DLH_X1 \CAM_MEM_reg[9][14]  ( .G(N878), .D(TAG_IN[14]), .Q(\CAM_MEM[9][14] )
         );
  DLH_X1 \CAM_MEM_reg[9][13]  ( .G(N878), .D(TAG_IN[13]), .Q(\CAM_MEM[9][13] )
         );
  DLH_X1 \CAM_MEM_reg[9][12]  ( .G(N878), .D(TAG_IN[12]), .Q(\CAM_MEM[9][12] )
         );
  DLH_X1 \CAM_MEM_reg[9][11]  ( .G(N878), .D(TAG_IN[11]), .Q(\CAM_MEM[9][11] )
         );
  DLH_X1 \CAM_MEM_reg[9][10]  ( .G(N878), .D(TAG_IN[10]), .Q(\CAM_MEM[9][10] )
         );
  DLH_X1 \CAM_MEM_reg[9][9]  ( .G(N878), .D(TAG_IN[9]), .Q(\CAM_MEM[9][9] ) );
  DLH_X1 \CAM_MEM_reg[9][8]  ( .G(N878), .D(TAG_IN[8]), .Q(\CAM_MEM[9][8] ) );
  DLH_X1 \CAM_MEM_reg[9][7]  ( .G(N878), .D(TAG_IN[7]), .Q(\CAM_MEM[9][7] ) );
  DLH_X1 \CAM_MEM_reg[9][6]  ( .G(N878), .D(TAG_IN[6]), .Q(\CAM_MEM[9][6] ) );
  DLH_X1 \CAM_MEM_reg[9][5]  ( .G(N878), .D(TAG_IN[5]), .Q(\CAM_MEM[9][5] ) );
  DLH_X1 \CAM_MEM_reg[9][4]  ( .G(N878), .D(TAG_IN[4]), .Q(\CAM_MEM[9][4] ) );
  DLH_X1 \CAM_MEM_reg[9][3]  ( .G(N878), .D(TAG_IN[3]), .Q(\CAM_MEM[9][3] ) );
  DLH_X1 \CAM_MEM_reg[9][2]  ( .G(N878), .D(TAG_IN[2]), .Q(\CAM_MEM[9][2] ) );
  DLH_X1 \CAM_MEM_reg[9][1]  ( .G(N878), .D(TAG_IN[1]), .Q(\CAM_MEM[9][1] ) );
  DLH_X1 \CAM_MEM_reg[9][0]  ( .G(N878), .D(TAG_IN[0]), .Q(\CAM_MEM[9][0] ) );
  DLH_X1 \CAM_MEM_reg[8][22]  ( .G(N855), .D(TAG_IN[22]), .Q(\CAM_MEM[8][22] )
         );
  DLH_X1 \CAM_MEM_reg[8][21]  ( .G(N855), .D(TAG_IN[21]), .Q(\CAM_MEM[8][21] )
         );
  DLH_X1 \CAM_MEM_reg[8][20]  ( .G(N855), .D(TAG_IN[20]), .Q(\CAM_MEM[8][20] )
         );
  DLH_X1 \CAM_MEM_reg[8][19]  ( .G(N855), .D(TAG_IN[19]), .Q(\CAM_MEM[8][19] )
         );
  DLH_X1 \CAM_MEM_reg[8][18]  ( .G(N855), .D(TAG_IN[18]), .Q(\CAM_MEM[8][18] )
         );
  DLH_X1 \CAM_MEM_reg[8][17]  ( .G(N855), .D(TAG_IN[17]), .Q(\CAM_MEM[8][17] )
         );
  DLH_X1 \CAM_MEM_reg[8][16]  ( .G(N855), .D(TAG_IN[16]), .Q(\CAM_MEM[8][16] )
         );
  DLH_X1 \CAM_MEM_reg[8][15]  ( .G(N855), .D(TAG_IN[15]), .Q(\CAM_MEM[8][15] )
         );
  DLH_X1 \CAM_MEM_reg[8][14]  ( .G(N855), .D(TAG_IN[14]), .Q(\CAM_MEM[8][14] )
         );
  DLH_X1 \CAM_MEM_reg[8][13]  ( .G(N855), .D(TAG_IN[13]), .Q(\CAM_MEM[8][13] )
         );
  DLH_X1 \CAM_MEM_reg[8][12]  ( .G(N855), .D(TAG_IN[12]), .Q(\CAM_MEM[8][12] )
         );
  DLH_X1 \CAM_MEM_reg[8][11]  ( .G(N855), .D(TAG_IN[11]), .Q(\CAM_MEM[8][11] )
         );
  DLH_X1 \CAM_MEM_reg[8][10]  ( .G(N855), .D(TAG_IN[10]), .Q(\CAM_MEM[8][10] )
         );
  DLH_X1 \CAM_MEM_reg[8][9]  ( .G(N855), .D(TAG_IN[9]), .Q(\CAM_MEM[8][9] ) );
  DLH_X1 \CAM_MEM_reg[8][8]  ( .G(N855), .D(TAG_IN[8]), .Q(\CAM_MEM[8][8] ) );
  DLH_X1 \CAM_MEM_reg[8][7]  ( .G(N855), .D(TAG_IN[7]), .Q(\CAM_MEM[8][7] ) );
  DLH_X1 \CAM_MEM_reg[8][6]  ( .G(N855), .D(TAG_IN[6]), .Q(\CAM_MEM[8][6] ) );
  DLH_X1 \CAM_MEM_reg[8][5]  ( .G(N855), .D(TAG_IN[5]), .Q(\CAM_MEM[8][5] ) );
  DLH_X1 \CAM_MEM_reg[8][4]  ( .G(N855), .D(TAG_IN[4]), .Q(\CAM_MEM[8][4] ) );
  DLH_X1 \CAM_MEM_reg[8][3]  ( .G(N855), .D(TAG_IN[3]), .Q(\CAM_MEM[8][3] ) );
  DLH_X1 \CAM_MEM_reg[8][2]  ( .G(N855), .D(TAG_IN[2]), .Q(\CAM_MEM[8][2] ) );
  DLH_X1 \CAM_MEM_reg[8][1]  ( .G(N855), .D(TAG_IN[1]), .Q(\CAM_MEM[8][1] ) );
  DLH_X1 \CAM_MEM_reg[8][0]  ( .G(N855), .D(TAG_IN[0]), .Q(\CAM_MEM[8][0] ) );
  DLH_X1 \CAM_MEM_reg[7][22]  ( .G(N832), .D(TAG_IN[22]), .Q(\CAM_MEM[7][22] )
         );
  DLH_X1 \CAM_MEM_reg[7][21]  ( .G(N832), .D(TAG_IN[21]), .Q(\CAM_MEM[7][21] )
         );
  DLH_X1 \CAM_MEM_reg[7][20]  ( .G(N832), .D(TAG_IN[20]), .Q(\CAM_MEM[7][20] )
         );
  DLH_X1 \CAM_MEM_reg[7][19]  ( .G(N832), .D(TAG_IN[19]), .Q(\CAM_MEM[7][19] )
         );
  DLH_X1 \CAM_MEM_reg[7][18]  ( .G(N832), .D(TAG_IN[18]), .Q(\CAM_MEM[7][18] )
         );
  DLH_X1 \CAM_MEM_reg[7][17]  ( .G(N832), .D(TAG_IN[17]), .Q(\CAM_MEM[7][17] )
         );
  DLH_X1 \CAM_MEM_reg[7][16]  ( .G(N832), .D(TAG_IN[16]), .Q(\CAM_MEM[7][16] )
         );
  DLH_X1 \CAM_MEM_reg[7][15]  ( .G(N832), .D(TAG_IN[15]), .Q(\CAM_MEM[7][15] )
         );
  DLH_X1 \CAM_MEM_reg[7][14]  ( .G(N832), .D(TAG_IN[14]), .Q(\CAM_MEM[7][14] )
         );
  DLH_X1 \CAM_MEM_reg[7][13]  ( .G(N832), .D(TAG_IN[13]), .Q(\CAM_MEM[7][13] )
         );
  DLH_X1 \CAM_MEM_reg[7][12]  ( .G(N832), .D(TAG_IN[12]), .Q(\CAM_MEM[7][12] )
         );
  DLH_X1 \CAM_MEM_reg[7][11]  ( .G(N832), .D(TAG_IN[11]), .Q(\CAM_MEM[7][11] )
         );
  DLH_X1 \CAM_MEM_reg[7][10]  ( .G(N832), .D(TAG_IN[10]), .Q(\CAM_MEM[7][10] )
         );
  DLH_X1 \CAM_MEM_reg[7][9]  ( .G(N832), .D(TAG_IN[9]), .Q(\CAM_MEM[7][9] ) );
  DLH_X1 \CAM_MEM_reg[7][8]  ( .G(N832), .D(TAG_IN[8]), .Q(\CAM_MEM[7][8] ) );
  DLH_X1 \CAM_MEM_reg[7][7]  ( .G(N832), .D(TAG_IN[7]), .Q(\CAM_MEM[7][7] ) );
  DLH_X1 \CAM_MEM_reg[7][6]  ( .G(N832), .D(TAG_IN[6]), .Q(\CAM_MEM[7][6] ) );
  DLH_X1 \CAM_MEM_reg[7][5]  ( .G(N832), .D(TAG_IN[5]), .Q(\CAM_MEM[7][5] ) );
  DLH_X1 \CAM_MEM_reg[7][4]  ( .G(N832), .D(TAG_IN[4]), .Q(\CAM_MEM[7][4] ) );
  DLH_X1 \CAM_MEM_reg[7][3]  ( .G(N832), .D(TAG_IN[3]), .Q(\CAM_MEM[7][3] ) );
  DLH_X1 \CAM_MEM_reg[7][2]  ( .G(N832), .D(TAG_IN[2]), .Q(\CAM_MEM[7][2] ) );
  DLH_X1 \CAM_MEM_reg[7][1]  ( .G(N832), .D(TAG_IN[1]), .Q(\CAM_MEM[7][1] ) );
  DLH_X1 \CAM_MEM_reg[7][0]  ( .G(N832), .D(TAG_IN[0]), .Q(\CAM_MEM[7][0] ) );
  DLH_X1 \CAM_MEM_reg[6][22]  ( .G(N809), .D(TAG_IN[22]), .Q(\CAM_MEM[6][22] )
         );
  DLH_X1 \CAM_MEM_reg[6][21]  ( .G(N809), .D(TAG_IN[21]), .Q(\CAM_MEM[6][21] )
         );
  DLH_X1 \CAM_MEM_reg[6][20]  ( .G(N809), .D(TAG_IN[20]), .Q(\CAM_MEM[6][20] )
         );
  DLH_X1 \CAM_MEM_reg[6][19]  ( .G(N809), .D(TAG_IN[19]), .Q(\CAM_MEM[6][19] )
         );
  DLH_X1 \CAM_MEM_reg[6][18]  ( .G(N809), .D(TAG_IN[18]), .Q(\CAM_MEM[6][18] )
         );
  DLH_X1 \CAM_MEM_reg[6][17]  ( .G(N809), .D(TAG_IN[17]), .Q(\CAM_MEM[6][17] )
         );
  DLH_X1 \CAM_MEM_reg[6][16]  ( .G(N809), .D(TAG_IN[16]), .Q(\CAM_MEM[6][16] )
         );
  DLH_X1 \CAM_MEM_reg[6][15]  ( .G(N809), .D(TAG_IN[15]), .Q(\CAM_MEM[6][15] )
         );
  DLH_X1 \CAM_MEM_reg[6][14]  ( .G(N809), .D(TAG_IN[14]), .Q(\CAM_MEM[6][14] )
         );
  DLH_X1 \CAM_MEM_reg[6][13]  ( .G(N809), .D(TAG_IN[13]), .Q(\CAM_MEM[6][13] )
         );
  DLH_X1 \CAM_MEM_reg[6][12]  ( .G(N809), .D(TAG_IN[12]), .Q(\CAM_MEM[6][12] )
         );
  DLH_X1 \CAM_MEM_reg[6][11]  ( .G(N809), .D(TAG_IN[11]), .Q(\CAM_MEM[6][11] )
         );
  DLH_X1 \CAM_MEM_reg[6][10]  ( .G(N809), .D(TAG_IN[10]), .Q(\CAM_MEM[6][10] )
         );
  DLH_X1 \CAM_MEM_reg[6][9]  ( .G(N809), .D(TAG_IN[9]), .Q(\CAM_MEM[6][9] ) );
  DLH_X1 \CAM_MEM_reg[6][8]  ( .G(N809), .D(TAG_IN[8]), .Q(\CAM_MEM[6][8] ) );
  DLH_X1 \CAM_MEM_reg[6][7]  ( .G(N809), .D(TAG_IN[7]), .Q(\CAM_MEM[6][7] ) );
  DLH_X1 \CAM_MEM_reg[6][6]  ( .G(N809), .D(TAG_IN[6]), .Q(\CAM_MEM[6][6] ) );
  DLH_X1 \CAM_MEM_reg[6][5]  ( .G(N809), .D(TAG_IN[5]), .Q(\CAM_MEM[6][5] ) );
  DLH_X1 \CAM_MEM_reg[6][4]  ( .G(N809), .D(TAG_IN[4]), .Q(\CAM_MEM[6][4] ) );
  DLH_X1 \CAM_MEM_reg[6][3]  ( .G(N809), .D(TAG_IN[3]), .Q(\CAM_MEM[6][3] ) );
  DLH_X1 \CAM_MEM_reg[6][2]  ( .G(N809), .D(TAG_IN[2]), .Q(\CAM_MEM[6][2] ) );
  DLH_X1 \CAM_MEM_reg[6][1]  ( .G(N809), .D(TAG_IN[1]), .Q(\CAM_MEM[6][1] ) );
  DLH_X1 \CAM_MEM_reg[6][0]  ( .G(N809), .D(TAG_IN[0]), .Q(\CAM_MEM[6][0] ) );
  DLH_X1 \CAM_MEM_reg[5][22]  ( .G(N786), .D(TAG_IN[22]), .Q(\CAM_MEM[5][22] )
         );
  DLH_X1 \CAM_MEM_reg[5][21]  ( .G(N786), .D(TAG_IN[21]), .Q(\CAM_MEM[5][21] )
         );
  DLH_X1 \CAM_MEM_reg[5][20]  ( .G(N786), .D(TAG_IN[20]), .Q(\CAM_MEM[5][20] )
         );
  DLH_X1 \CAM_MEM_reg[5][19]  ( .G(N786), .D(TAG_IN[19]), .Q(\CAM_MEM[5][19] )
         );
  DLH_X1 \CAM_MEM_reg[5][18]  ( .G(N786), .D(TAG_IN[18]), .Q(\CAM_MEM[5][18] )
         );
  DLH_X1 \CAM_MEM_reg[5][17]  ( .G(N786), .D(TAG_IN[17]), .Q(\CAM_MEM[5][17] )
         );
  DLH_X1 \CAM_MEM_reg[5][16]  ( .G(N786), .D(TAG_IN[16]), .Q(\CAM_MEM[5][16] )
         );
  DLH_X1 \CAM_MEM_reg[5][15]  ( .G(N786), .D(TAG_IN[15]), .Q(\CAM_MEM[5][15] )
         );
  DLH_X1 \CAM_MEM_reg[5][14]  ( .G(N786), .D(TAG_IN[14]), .Q(\CAM_MEM[5][14] )
         );
  DLH_X1 \CAM_MEM_reg[5][13]  ( .G(N786), .D(TAG_IN[13]), .Q(\CAM_MEM[5][13] )
         );
  DLH_X1 \CAM_MEM_reg[5][12]  ( .G(N786), .D(TAG_IN[12]), .Q(\CAM_MEM[5][12] )
         );
  DLH_X1 \CAM_MEM_reg[5][11]  ( .G(N786), .D(TAG_IN[11]), .Q(\CAM_MEM[5][11] )
         );
  DLH_X1 \CAM_MEM_reg[5][10]  ( .G(N786), .D(TAG_IN[10]), .Q(\CAM_MEM[5][10] )
         );
  DLH_X1 \CAM_MEM_reg[5][9]  ( .G(N786), .D(TAG_IN[9]), .Q(\CAM_MEM[5][9] ) );
  DLH_X1 \CAM_MEM_reg[5][8]  ( .G(N786), .D(TAG_IN[8]), .Q(\CAM_MEM[5][8] ) );
  DLH_X1 \CAM_MEM_reg[5][7]  ( .G(N786), .D(TAG_IN[7]), .Q(\CAM_MEM[5][7] ) );
  DLH_X1 \CAM_MEM_reg[5][6]  ( .G(N786), .D(TAG_IN[6]), .Q(\CAM_MEM[5][6] ) );
  DLH_X1 \CAM_MEM_reg[5][5]  ( .G(N786), .D(TAG_IN[5]), .Q(\CAM_MEM[5][5] ) );
  DLH_X1 \CAM_MEM_reg[5][4]  ( .G(N786), .D(TAG_IN[4]), .Q(\CAM_MEM[5][4] ) );
  DLH_X1 \CAM_MEM_reg[5][3]  ( .G(N786), .D(TAG_IN[3]), .Q(\CAM_MEM[5][3] ) );
  DLH_X1 \CAM_MEM_reg[5][2]  ( .G(N786), .D(TAG_IN[2]), .Q(\CAM_MEM[5][2] ) );
  DLH_X1 \CAM_MEM_reg[5][1]  ( .G(N786), .D(TAG_IN[1]), .Q(\CAM_MEM[5][1] ) );
  DLH_X1 \CAM_MEM_reg[5][0]  ( .G(N786), .D(TAG_IN[0]), .Q(\CAM_MEM[5][0] ) );
  DLH_X1 \CAM_MEM_reg[4][22]  ( .G(N763), .D(TAG_IN[22]), .Q(\CAM_MEM[4][22] )
         );
  DLH_X1 \CAM_MEM_reg[4][21]  ( .G(N763), .D(TAG_IN[21]), .Q(\CAM_MEM[4][21] )
         );
  DLH_X1 \CAM_MEM_reg[4][20]  ( .G(N763), .D(TAG_IN[20]), .Q(\CAM_MEM[4][20] )
         );
  DLH_X1 \CAM_MEM_reg[4][19]  ( .G(N763), .D(TAG_IN[19]), .Q(\CAM_MEM[4][19] )
         );
  DLH_X1 \CAM_MEM_reg[4][18]  ( .G(N763), .D(TAG_IN[18]), .Q(\CAM_MEM[4][18] )
         );
  DLH_X1 \CAM_MEM_reg[4][17]  ( .G(N763), .D(TAG_IN[17]), .Q(\CAM_MEM[4][17] )
         );
  DLH_X1 \CAM_MEM_reg[4][16]  ( .G(N763), .D(TAG_IN[16]), .Q(\CAM_MEM[4][16] )
         );
  DLH_X1 \CAM_MEM_reg[4][15]  ( .G(N763), .D(TAG_IN[15]), .Q(\CAM_MEM[4][15] )
         );
  DLH_X1 \CAM_MEM_reg[4][14]  ( .G(N763), .D(TAG_IN[14]), .Q(\CAM_MEM[4][14] )
         );
  DLH_X1 \CAM_MEM_reg[4][13]  ( .G(N763), .D(TAG_IN[13]), .Q(\CAM_MEM[4][13] )
         );
  DLH_X1 \CAM_MEM_reg[4][12]  ( .G(N763), .D(TAG_IN[12]), .Q(\CAM_MEM[4][12] )
         );
  DLH_X1 \CAM_MEM_reg[4][11]  ( .G(N763), .D(TAG_IN[11]), .Q(\CAM_MEM[4][11] )
         );
  DLH_X1 \CAM_MEM_reg[4][10]  ( .G(N763), .D(TAG_IN[10]), .Q(\CAM_MEM[4][10] )
         );
  DLH_X1 \CAM_MEM_reg[4][9]  ( .G(N763), .D(TAG_IN[9]), .Q(\CAM_MEM[4][9] ) );
  DLH_X1 \CAM_MEM_reg[4][8]  ( .G(N763), .D(TAG_IN[8]), .Q(\CAM_MEM[4][8] ) );
  DLH_X1 \CAM_MEM_reg[4][7]  ( .G(N763), .D(TAG_IN[7]), .Q(\CAM_MEM[4][7] ) );
  DLH_X1 \CAM_MEM_reg[4][6]  ( .G(N763), .D(TAG_IN[6]), .Q(\CAM_MEM[4][6] ) );
  DLH_X1 \CAM_MEM_reg[4][5]  ( .G(N763), .D(TAG_IN[5]), .Q(\CAM_MEM[4][5] ) );
  DLH_X1 \CAM_MEM_reg[4][4]  ( .G(N763), .D(TAG_IN[4]), .Q(\CAM_MEM[4][4] ) );
  DLH_X1 \CAM_MEM_reg[4][3]  ( .G(N763), .D(TAG_IN[3]), .Q(\CAM_MEM[4][3] ) );
  DLH_X1 \CAM_MEM_reg[4][2]  ( .G(N763), .D(TAG_IN[2]), .Q(\CAM_MEM[4][2] ) );
  DLH_X1 \CAM_MEM_reg[4][1]  ( .G(N763), .D(TAG_IN[1]), .Q(\CAM_MEM[4][1] ) );
  DLH_X1 \CAM_MEM_reg[4][0]  ( .G(N763), .D(TAG_IN[0]), .Q(\CAM_MEM[4][0] ) );
  DLH_X1 \CAM_MEM_reg[3][22]  ( .G(N740), .D(TAG_IN[22]), .Q(\CAM_MEM[3][22] )
         );
  DLH_X1 \CAM_MEM_reg[3][21]  ( .G(N740), .D(TAG_IN[21]), .Q(\CAM_MEM[3][21] )
         );
  DLH_X1 \CAM_MEM_reg[3][20]  ( .G(N740), .D(TAG_IN[20]), .Q(\CAM_MEM[3][20] )
         );
  DLH_X1 \CAM_MEM_reg[3][19]  ( .G(N740), .D(TAG_IN[19]), .Q(\CAM_MEM[3][19] )
         );
  DLH_X1 \CAM_MEM_reg[3][18]  ( .G(N740), .D(TAG_IN[18]), .Q(\CAM_MEM[3][18] )
         );
  DLH_X1 \CAM_MEM_reg[3][17]  ( .G(N740), .D(TAG_IN[17]), .Q(\CAM_MEM[3][17] )
         );
  DLH_X1 \CAM_MEM_reg[3][16]  ( .G(N740), .D(TAG_IN[16]), .Q(\CAM_MEM[3][16] )
         );
  DLH_X1 \CAM_MEM_reg[3][15]  ( .G(N740), .D(TAG_IN[15]), .Q(\CAM_MEM[3][15] )
         );
  DLH_X1 \CAM_MEM_reg[3][14]  ( .G(N740), .D(TAG_IN[14]), .Q(\CAM_MEM[3][14] )
         );
  DLH_X1 \CAM_MEM_reg[3][13]  ( .G(N740), .D(TAG_IN[13]), .Q(\CAM_MEM[3][13] )
         );
  DLH_X1 \CAM_MEM_reg[3][12]  ( .G(N740), .D(TAG_IN[12]), .Q(\CAM_MEM[3][12] )
         );
  DLH_X1 \CAM_MEM_reg[3][11]  ( .G(N740), .D(TAG_IN[11]), .Q(\CAM_MEM[3][11] )
         );
  DLH_X1 \CAM_MEM_reg[3][10]  ( .G(N740), .D(TAG_IN[10]), .Q(\CAM_MEM[3][10] )
         );
  DLH_X1 \CAM_MEM_reg[3][9]  ( .G(N740), .D(TAG_IN[9]), .Q(\CAM_MEM[3][9] ) );
  DLH_X1 \CAM_MEM_reg[3][8]  ( .G(N740), .D(TAG_IN[8]), .Q(\CAM_MEM[3][8] ) );
  DLH_X1 \CAM_MEM_reg[3][7]  ( .G(N740), .D(TAG_IN[7]), .Q(\CAM_MEM[3][7] ) );
  DLH_X1 \CAM_MEM_reg[3][6]  ( .G(N740), .D(TAG_IN[6]), .Q(\CAM_MEM[3][6] ) );
  DLH_X1 \CAM_MEM_reg[3][5]  ( .G(N740), .D(TAG_IN[5]), .Q(\CAM_MEM[3][5] ) );
  DLH_X1 \CAM_MEM_reg[3][4]  ( .G(N740), .D(TAG_IN[4]), .Q(\CAM_MEM[3][4] ) );
  DLH_X1 \CAM_MEM_reg[3][3]  ( .G(N740), .D(TAG_IN[3]), .Q(\CAM_MEM[3][3] ) );
  DLH_X1 \CAM_MEM_reg[3][2]  ( .G(N740), .D(TAG_IN[2]), .Q(\CAM_MEM[3][2] ) );
  DLH_X1 \CAM_MEM_reg[3][1]  ( .G(N740), .D(TAG_IN[1]), .Q(\CAM_MEM[3][1] ) );
  DLH_X1 \CAM_MEM_reg[3][0]  ( .G(N740), .D(TAG_IN[0]), .Q(\CAM_MEM[3][0] ) );
  DLH_X1 \CAM_MEM_reg[2][22]  ( .G(N717), .D(TAG_IN[22]), .Q(\CAM_MEM[2][22] )
         );
  DLH_X1 \CAM_MEM_reg[2][21]  ( .G(N717), .D(TAG_IN[21]), .Q(\CAM_MEM[2][21] )
         );
  DLH_X1 \CAM_MEM_reg[2][20]  ( .G(N717), .D(TAG_IN[20]), .Q(\CAM_MEM[2][20] )
         );
  DLH_X1 \CAM_MEM_reg[2][19]  ( .G(N717), .D(TAG_IN[19]), .Q(\CAM_MEM[2][19] )
         );
  DLH_X1 \CAM_MEM_reg[2][18]  ( .G(N717), .D(TAG_IN[18]), .Q(\CAM_MEM[2][18] )
         );
  DLH_X1 \CAM_MEM_reg[2][17]  ( .G(N717), .D(TAG_IN[17]), .Q(\CAM_MEM[2][17] )
         );
  DLH_X1 \CAM_MEM_reg[2][16]  ( .G(N717), .D(TAG_IN[16]), .Q(\CAM_MEM[2][16] )
         );
  DLH_X1 \CAM_MEM_reg[2][15]  ( .G(N717), .D(TAG_IN[15]), .Q(\CAM_MEM[2][15] )
         );
  DLH_X1 \CAM_MEM_reg[2][14]  ( .G(N717), .D(TAG_IN[14]), .Q(\CAM_MEM[2][14] )
         );
  DLH_X1 \CAM_MEM_reg[2][13]  ( .G(N717), .D(TAG_IN[13]), .Q(\CAM_MEM[2][13] )
         );
  DLH_X1 \CAM_MEM_reg[2][12]  ( .G(N717), .D(TAG_IN[12]), .Q(\CAM_MEM[2][12] )
         );
  DLH_X1 \CAM_MEM_reg[2][11]  ( .G(N717), .D(TAG_IN[11]), .Q(\CAM_MEM[2][11] )
         );
  DLH_X1 \CAM_MEM_reg[2][10]  ( .G(N717), .D(TAG_IN[10]), .Q(\CAM_MEM[2][10] )
         );
  DLH_X1 \CAM_MEM_reg[2][9]  ( .G(N717), .D(TAG_IN[9]), .Q(\CAM_MEM[2][9] ) );
  DLH_X1 \CAM_MEM_reg[2][8]  ( .G(N717), .D(TAG_IN[8]), .Q(\CAM_MEM[2][8] ) );
  DLH_X1 \CAM_MEM_reg[2][7]  ( .G(N717), .D(TAG_IN[7]), .Q(\CAM_MEM[2][7] ) );
  DLH_X1 \CAM_MEM_reg[2][6]  ( .G(N717), .D(TAG_IN[6]), .Q(\CAM_MEM[2][6] ) );
  DLH_X1 \CAM_MEM_reg[2][5]  ( .G(N717), .D(TAG_IN[5]), .Q(\CAM_MEM[2][5] ) );
  DLH_X1 \CAM_MEM_reg[2][4]  ( .G(N717), .D(TAG_IN[4]), .Q(\CAM_MEM[2][4] ) );
  DLH_X1 \CAM_MEM_reg[2][3]  ( .G(N717), .D(TAG_IN[3]), .Q(\CAM_MEM[2][3] ) );
  DLH_X1 \CAM_MEM_reg[2][2]  ( .G(N717), .D(TAG_IN[2]), .Q(\CAM_MEM[2][2] ) );
  DLH_X1 \CAM_MEM_reg[2][1]  ( .G(N717), .D(TAG_IN[1]), .Q(\CAM_MEM[2][1] ) );
  DLH_X1 \CAM_MEM_reg[2][0]  ( .G(N717), .D(TAG_IN[0]), .Q(\CAM_MEM[2][0] ) );
  DLH_X1 \CAM_MEM_reg[1][22]  ( .G(N694), .D(TAG_IN[22]), .Q(\CAM_MEM[1][22] )
         );
  DLH_X1 \CAM_MEM_reg[1][21]  ( .G(N694), .D(TAG_IN[21]), .Q(\CAM_MEM[1][21] )
         );
  DLH_X1 \CAM_MEM_reg[1][20]  ( .G(N694), .D(TAG_IN[20]), .Q(\CAM_MEM[1][20] )
         );
  DLH_X1 \CAM_MEM_reg[1][19]  ( .G(N694), .D(TAG_IN[19]), .Q(\CAM_MEM[1][19] )
         );
  DLH_X1 \CAM_MEM_reg[1][18]  ( .G(N694), .D(TAG_IN[18]), .Q(\CAM_MEM[1][18] )
         );
  DLH_X1 \CAM_MEM_reg[1][17]  ( .G(N694), .D(TAG_IN[17]), .Q(\CAM_MEM[1][17] )
         );
  DLH_X1 \CAM_MEM_reg[1][16]  ( .G(N694), .D(TAG_IN[16]), .Q(\CAM_MEM[1][16] )
         );
  DLH_X1 \CAM_MEM_reg[1][15]  ( .G(N694), .D(TAG_IN[15]), .Q(\CAM_MEM[1][15] )
         );
  DLH_X1 \CAM_MEM_reg[1][14]  ( .G(N694), .D(TAG_IN[14]), .Q(\CAM_MEM[1][14] )
         );
  DLH_X1 \CAM_MEM_reg[1][13]  ( .G(N694), .D(TAG_IN[13]), .Q(\CAM_MEM[1][13] )
         );
  DLH_X1 \CAM_MEM_reg[1][12]  ( .G(N694), .D(TAG_IN[12]), .Q(\CAM_MEM[1][12] )
         );
  DLH_X1 \CAM_MEM_reg[1][11]  ( .G(N694), .D(TAG_IN[11]), .Q(\CAM_MEM[1][11] )
         );
  DLH_X1 \CAM_MEM_reg[1][10]  ( .G(N694), .D(TAG_IN[10]), .Q(\CAM_MEM[1][10] )
         );
  DLH_X1 \CAM_MEM_reg[1][9]  ( .G(N694), .D(TAG_IN[9]), .Q(\CAM_MEM[1][9] ) );
  DLH_X1 \CAM_MEM_reg[1][8]  ( .G(N694), .D(TAG_IN[8]), .Q(\CAM_MEM[1][8] ) );
  DLH_X1 \CAM_MEM_reg[1][7]  ( .G(N694), .D(TAG_IN[7]), .Q(\CAM_MEM[1][7] ) );
  DLH_X1 \CAM_MEM_reg[1][6]  ( .G(N694), .D(TAG_IN[6]), .Q(\CAM_MEM[1][6] ) );
  DLH_X1 \CAM_MEM_reg[1][5]  ( .G(N694), .D(TAG_IN[5]), .Q(\CAM_MEM[1][5] ) );
  DLH_X1 \CAM_MEM_reg[1][4]  ( .G(N694), .D(TAG_IN[4]), .Q(\CAM_MEM[1][4] ) );
  DLH_X1 \CAM_MEM_reg[1][3]  ( .G(N694), .D(TAG_IN[3]), .Q(\CAM_MEM[1][3] ) );
  DLH_X1 \CAM_MEM_reg[1][2]  ( .G(N694), .D(TAG_IN[2]), .Q(\CAM_MEM[1][2] ) );
  DLH_X1 \CAM_MEM_reg[1][1]  ( .G(N694), .D(TAG_IN[1]), .Q(\CAM_MEM[1][1] ) );
  DLH_X1 \CAM_MEM_reg[1][0]  ( .G(N694), .D(TAG_IN[0]), .Q(\CAM_MEM[1][0] ) );
  DLH_X1 \CAM_MEM_reg[0][22]  ( .G(N671), .D(TAG_IN[22]), .Q(\CAM_MEM[0][22] )
         );
  DLH_X1 \CAM_MEM_reg[0][21]  ( .G(N671), .D(TAG_IN[21]), .Q(\CAM_MEM[0][21] )
         );
  DLH_X1 \CAM_MEM_reg[0][20]  ( .G(N671), .D(TAG_IN[20]), .Q(\CAM_MEM[0][20] )
         );
  DLH_X1 \CAM_MEM_reg[0][19]  ( .G(N671), .D(TAG_IN[19]), .Q(\CAM_MEM[0][19] )
         );
  DLH_X1 \CAM_MEM_reg[0][18]  ( .G(N671), .D(TAG_IN[18]), .Q(\CAM_MEM[0][18] )
         );
  DLH_X1 \CAM_MEM_reg[0][17]  ( .G(N671), .D(TAG_IN[17]), .Q(\CAM_MEM[0][17] )
         );
  DLH_X1 \CAM_MEM_reg[0][16]  ( .G(N671), .D(TAG_IN[16]), .Q(\CAM_MEM[0][16] )
         );
  DLH_X1 \CAM_MEM_reg[0][15]  ( .G(N671), .D(TAG_IN[15]), .Q(\CAM_MEM[0][15] )
         );
  DLH_X1 \CAM_MEM_reg[0][14]  ( .G(N671), .D(TAG_IN[14]), .Q(\CAM_MEM[0][14] )
         );
  DLH_X1 \CAM_MEM_reg[0][13]  ( .G(N671), .D(TAG_IN[13]), .Q(\CAM_MEM[0][13] )
         );
  DLH_X1 \CAM_MEM_reg[0][12]  ( .G(N671), .D(TAG_IN[12]), .Q(\CAM_MEM[0][12] )
         );
  DLH_X1 \CAM_MEM_reg[0][11]  ( .G(N671), .D(TAG_IN[11]), .Q(\CAM_MEM[0][11] )
         );
  DLH_X1 \CAM_MEM_reg[0][10]  ( .G(N671), .D(TAG_IN[10]), .Q(\CAM_MEM[0][10] )
         );
  DLH_X1 \CAM_MEM_reg[0][9]  ( .G(N671), .D(TAG_IN[9]), .Q(\CAM_MEM[0][9] ) );
  DLH_X1 \CAM_MEM_reg[0][8]  ( .G(N671), .D(TAG_IN[8]), .Q(\CAM_MEM[0][8] ) );
  DLH_X1 \CAM_MEM_reg[0][7]  ( .G(N671), .D(TAG_IN[7]), .Q(\CAM_MEM[0][7] ) );
  DLH_X1 \CAM_MEM_reg[0][6]  ( .G(N671), .D(TAG_IN[6]), .Q(\CAM_MEM[0][6] ) );
  DLH_X1 \CAM_MEM_reg[0][5]  ( .G(N671), .D(TAG_IN[5]), .Q(\CAM_MEM[0][5] ) );
  DLH_X1 \CAM_MEM_reg[0][4]  ( .G(N671), .D(TAG_IN[4]), .Q(\CAM_MEM[0][4] ) );
  DLH_X1 \CAM_MEM_reg[0][3]  ( .G(N671), .D(TAG_IN[3]), .Q(\CAM_MEM[0][3] ) );
  DLH_X1 \CAM_MEM_reg[0][2]  ( .G(N671), .D(TAG_IN[2]), .Q(\CAM_MEM[0][2] ) );
  DLH_X1 \CAM_MEM_reg[0][1]  ( .G(N671), .D(TAG_IN[1]), .Q(\CAM_MEM[0][1] ) );
  DLH_X1 \CAM_MEM_reg[0][0]  ( .G(N671), .D(TAG_IN[0]), .Q(\CAM_MEM[0][0] ) );
  NAND3_X1 U3 ( .A1(n2), .A2(n3), .A3(N221), .ZN(n29) );
  NAND2_X1 U13 ( .A1(SET_INDEX[0]), .A2(n11), .ZN(n5) );
  NAND2_X1 U15 ( .A1(n11), .A2(n392), .ZN(n7) );
  NAND2_X1 U24 ( .A1(n16), .A2(SET_INDEX[0]), .ZN(n14) );
  NAND2_X1 U26 ( .A1(n16), .A2(n392), .ZN(n15) );
  NAND2_X1 U28 ( .A1(WE), .A2(n399), .ZN(n3) );
  NAND2_X1 U36 ( .A1(n19), .A2(SET_INDEX[0]), .ZN(n17) );
  NAND2_X1 U38 ( .A1(n19), .A2(n392), .ZN(n18) );
  NAND2_X1 U42 ( .A1(SET_INDEX[2]), .A2(SET_INDEX[1]), .ZN(n6) );
  NAND2_X1 U45 ( .A1(SET_INDEX[2]), .A2(n393), .ZN(n8) );
  NAND2_X1 U48 ( .A1(SET_INDEX[1]), .A2(n394), .ZN(n9) );
  NAND2_X1 U50 ( .A1(n24), .A2(SET_INDEX[0]), .ZN(n20) );
  NAND2_X1 U52 ( .A1(n24), .A2(n392), .ZN(n21) );
  NAND2_X1 U56 ( .A1(n393), .A2(n394), .ZN(n10) );
  NAND3_X1 U63 ( .A1(COUNT[4]), .A2(COUNT[3]), .A3(WE), .ZN(n27) );
  NAND3_X1 U64 ( .A1(COUNT[1]), .A2(COUNT[0]), .A3(COUNT[2]), .ZN(n26) );
  DFFRS_X1 VALID_reg ( .D(n30), .CK(CLK), .RN(n31), .SN(n29), .Q(VALID), .QN(
        n28) );
  INV_X1 U4 ( .A(n396), .ZN(n399) );
  BUF_X1 U5 ( .A(SET_INDEX[3]), .Z(n363) );
  BUF_X1 U6 ( .A(RST), .Z(n396) );
  NOR2_X1 U7 ( .A1(n6), .A2(n14), .ZN(N832) );
  NOR2_X1 U8 ( .A1(n5), .A2(n6), .ZN(N999) );
  NOR2_X1 U9 ( .A1(n3), .A2(SET_INDEX[3]), .ZN(n16) );
  OAI21_X1 U10 ( .B1(n6), .B2(n20), .A(n399), .ZN(N638) );
  OAI21_X1 U11 ( .B1(n6), .B2(n17), .A(n399), .ZN(N646) );
  BUF_X1 U12 ( .A(SET_INDEX[3]), .Z(n364) );
  BUF_X1 U14 ( .A(SET_INDEX[3]), .Z(n365) );
  BUF_X1 U16 ( .A(SET_INDEX[3]), .Z(n366) );
  BUF_X1 U17 ( .A(SET_INDEX[3]), .Z(n367) );
  BUF_X1 U18 ( .A(SET_INDEX[3]), .Z(n368) );
  BUF_X1 U19 ( .A(SET_INDEX[3]), .Z(n369) );
  BUF_X1 U20 ( .A(SET_INDEX[3]), .Z(n370) );
  BUF_X1 U21 ( .A(SET_INDEX[3]), .Z(n371) );
  BUF_X1 U22 ( .A(SET_INDEX[3]), .Z(n372) );
  BUF_X1 U23 ( .A(SET_INDEX[3]), .Z(n373) );
  BUF_X1 U25 ( .A(SET_INDEX[3]), .Z(n374) );
  BUF_X1 U27 ( .A(SET_INDEX[3]), .Z(n375) );
  BUF_X1 U29 ( .A(SET_INDEX[3]), .Z(n376) );
  BUF_X1 U30 ( .A(SET_INDEX[3]), .Z(n377) );
  BUF_X1 U31 ( .A(RST), .Z(n397) );
  BUF_X1 U32 ( .A(RST), .Z(n398) );
  BUF_X1 U33 ( .A(SET_INDEX[1]), .Z(n387) );
  BUF_X1 U34 ( .A(SET_INDEX[0]), .Z(n388) );
  INV_X1 U35 ( .A(N221), .ZN(n4) );
  NOR2_X1 U37 ( .A1(n8), .A2(n15), .ZN(N763) );
  NOR2_X1 U39 ( .A1(n8), .A2(n14), .ZN(N786) );
  NOR2_X1 U40 ( .A1(n6), .A2(n15), .ZN(N809) );
  NOR2_X1 U41 ( .A1(n6), .A2(n7), .ZN(N993) );
  NOR2_X1 U43 ( .A1(n9), .A2(n15), .ZN(N717) );
  NOR2_X1 U44 ( .A1(n9), .A2(n14), .ZN(N740) );
  NOR2_X1 U46 ( .A1(n10), .A2(n15), .ZN(N671) );
  NOR2_X1 U47 ( .A1(n10), .A2(n14), .ZN(N694) );
  NOR2_X1 U49 ( .A1(n7), .A2(n8), .ZN(N947) );
  NOR2_X1 U51 ( .A1(n5), .A2(n8), .ZN(N970) );
  NOR2_X1 U53 ( .A1(n7), .A2(n9), .ZN(N901) );
  NOR2_X1 U54 ( .A1(n5), .A2(n9), .ZN(N924) );
  NOR2_X1 U55 ( .A1(n7), .A2(n10), .ZN(N855) );
  NOR2_X1 U57 ( .A1(n5), .A2(n10), .ZN(N878) );
  OAI21_X1 U58 ( .B1(n8), .B2(n21), .A(n399), .ZN(N635) );
  OAI21_X1 U59 ( .B1(n8), .B2(n20), .A(n399), .ZN(N636) );
  OAI21_X1 U60 ( .B1(n8), .B2(n18), .A(n399), .ZN(N643) );
  OAI21_X1 U61 ( .B1(n8), .B2(n17), .A(n399), .ZN(N644) );
  OAI21_X1 U62 ( .B1(n6), .B2(n21), .A(n399), .ZN(N637) );
  OAI21_X1 U65 ( .B1(n6), .B2(n18), .A(n399), .ZN(N645) );
  OAI21_X1 U66 ( .B1(n9), .B2(n21), .A(n399), .ZN(N633) );
  OAI21_X1 U67 ( .B1(n9), .B2(n20), .A(n399), .ZN(N634) );
  OAI21_X1 U68 ( .B1(n9), .B2(n18), .A(n399), .ZN(N641) );
  OAI21_X1 U69 ( .B1(n9), .B2(n17), .A(n399), .ZN(N642) );
  OAI21_X1 U70 ( .B1(n10), .B2(n21), .A(n399), .ZN(N631) );
  OAI21_X1 U71 ( .B1(n10), .B2(n20), .A(n399), .ZN(N632) );
  OAI21_X1 U72 ( .B1(n10), .B2(n18), .A(n399), .ZN(N639) );
  OAI21_X1 U73 ( .B1(n10), .B2(n17), .A(n399), .ZN(N640) );
  BUF_X1 U74 ( .A(SET_INDEX[2]), .Z(n379) );
  BUF_X1 U75 ( .A(SET_INDEX[2]), .Z(n380) );
  BUF_X1 U76 ( .A(SET_INDEX[2]), .Z(n381) );
  BUF_X1 U77 ( .A(SET_INDEX[2]), .Z(n382) );
  BUF_X1 U78 ( .A(SET_INDEX[2]), .Z(n383) );
  BUF_X1 U79 ( .A(SET_INDEX[2]), .Z(n384) );
  BUF_X1 U80 ( .A(SET_INDEX[2]), .Z(n385) );
  BUF_X1 U81 ( .A(SET_INDEX[0]), .Z(n389) );
  BUF_X1 U82 ( .A(SET_INDEX[0]), .Z(n390) );
  BUF_X1 U83 ( .A(SET_INDEX[0]), .Z(n391) );
  NOR2_X1 U84 ( .A1(n395), .A2(n3), .ZN(n11) );
  BUF_X1 U85 ( .A(SET_INDEX[1]), .Z(n386) );
  AND2_X1 U86 ( .A1(SET_INDEX[3]), .A2(WE), .ZN(n19) );
  AND2_X1 U87 ( .A1(WE), .A2(n395), .ZN(n24) );
  OAI21_X1 U88 ( .B1(WE), .B2(n4), .A(n2), .ZN(n31) );
  OAI22_X1 U89 ( .A1(n28), .A2(n399), .B1(n396), .B2(n4), .ZN(n30) );
  INV_X1 U90 ( .A(SET_INDEX[0]), .ZN(n392) );
  INV_X1 U91 ( .A(n25), .ZN(n2) );
  OAI21_X1 U92 ( .B1(n26), .B2(n27), .A(n399), .ZN(n25) );
  MUX2_X1 U93 ( .A(VALID_BIT[7]), .B(VALID_BIT[15]), .S(n363), .Z(n1) );
  MUX2_X1 U94 ( .A(VALID_BIT[3]), .B(VALID_BIT[11]), .S(n363), .Z(n12) );
  MUX2_X1 U95 ( .A(n12), .B(n1), .S(n378), .Z(n13) );
  MUX2_X1 U96 ( .A(VALID_BIT[6]), .B(VALID_BIT[14]), .S(n363), .Z(n22) );
  MUX2_X1 U97 ( .A(VALID_BIT[2]), .B(VALID_BIT[10]), .S(n363), .Z(n23) );
  MUX2_X1 U98 ( .A(n23), .B(n22), .S(n378), .Z(n32) );
  MUX2_X1 U99 ( .A(n32), .B(n13), .S(n388), .Z(n33) );
  MUX2_X1 U100 ( .A(VALID_BIT[5]), .B(VALID_BIT[13]), .S(n363), .Z(n34) );
  MUX2_X1 U101 ( .A(VALID_BIT[1]), .B(VALID_BIT[9]), .S(n363), .Z(n35) );
  MUX2_X1 U102 ( .A(n35), .B(n34), .S(n378), .Z(n36) );
  MUX2_X1 U103 ( .A(VALID_BIT[4]), .B(VALID_BIT[12]), .S(n363), .Z(n37) );
  MUX2_X1 U104 ( .A(VALID_BIT[0]), .B(VALID_BIT[8]), .S(n363), .Z(n38) );
  MUX2_X1 U105 ( .A(n38), .B(n37), .S(n378), .Z(n39) );
  MUX2_X1 U106 ( .A(n39), .B(n36), .S(n388), .Z(n40) );
  MUX2_X1 U107 ( .A(n40), .B(n33), .S(n387), .Z(N221) );
  MUX2_X1 U108 ( .A(\CAM_MEM[7][0] ), .B(\CAM_MEM[15][0] ), .S(n363), .Z(n41)
         );
  MUX2_X1 U109 ( .A(\CAM_MEM[3][0] ), .B(\CAM_MEM[11][0] ), .S(n363), .Z(n42)
         );
  MUX2_X1 U110 ( .A(n42), .B(n41), .S(n378), .Z(n43) );
  MUX2_X1 U111 ( .A(\CAM_MEM[6][0] ), .B(\CAM_MEM[14][0] ), .S(n364), .Z(n44)
         );
  MUX2_X1 U112 ( .A(\CAM_MEM[2][0] ), .B(\CAM_MEM[10][0] ), .S(n364), .Z(n45)
         );
  MUX2_X1 U113 ( .A(n45), .B(n44), .S(n379), .Z(n46) );
  MUX2_X1 U114 ( .A(n46), .B(n43), .S(n388), .Z(n47) );
  MUX2_X1 U115 ( .A(\CAM_MEM[5][0] ), .B(\CAM_MEM[13][0] ), .S(n364), .Z(n48)
         );
  MUX2_X1 U116 ( .A(\CAM_MEM[1][0] ), .B(\CAM_MEM[9][0] ), .S(n364), .Z(n49)
         );
  MUX2_X1 U117 ( .A(n49), .B(n48), .S(n379), .Z(n50) );
  MUX2_X1 U118 ( .A(\CAM_MEM[4][0] ), .B(\CAM_MEM[12][0] ), .S(n364), .Z(n51)
         );
  MUX2_X1 U119 ( .A(\CAM_MEM[0][0] ), .B(\CAM_MEM[8][0] ), .S(n364), .Z(n52)
         );
  MUX2_X1 U120 ( .A(n52), .B(n51), .S(n379), .Z(n53) );
  MUX2_X1 U121 ( .A(n53), .B(n50), .S(n388), .Z(n54) );
  MUX2_X1 U122 ( .A(n54), .B(n47), .S(n387), .Z(N606) );
  MUX2_X1 U123 ( .A(\CAM_MEM[7][1] ), .B(\CAM_MEM[15][1] ), .S(n364), .Z(n55)
         );
  MUX2_X1 U124 ( .A(\CAM_MEM[3][1] ), .B(\CAM_MEM[11][1] ), .S(n364), .Z(n56)
         );
  MUX2_X1 U125 ( .A(n56), .B(n55), .S(n379), .Z(n57) );
  MUX2_X1 U126 ( .A(\CAM_MEM[6][1] ), .B(\CAM_MEM[14][1] ), .S(n364), .Z(n58)
         );
  MUX2_X1 U127 ( .A(\CAM_MEM[2][1] ), .B(\CAM_MEM[10][1] ), .S(n364), .Z(n59)
         );
  MUX2_X1 U128 ( .A(n59), .B(n58), .S(n379), .Z(n60) );
  MUX2_X1 U129 ( .A(n60), .B(n57), .S(n388), .Z(n61) );
  MUX2_X1 U130 ( .A(\CAM_MEM[5][1] ), .B(\CAM_MEM[13][1] ), .S(n364), .Z(n62)
         );
  MUX2_X1 U131 ( .A(\CAM_MEM[1][1] ), .B(\CAM_MEM[9][1] ), .S(n364), .Z(n63)
         );
  MUX2_X1 U132 ( .A(n63), .B(n62), .S(n379), .Z(n64) );
  MUX2_X1 U133 ( .A(\CAM_MEM[4][1] ), .B(\CAM_MEM[12][1] ), .S(n364), .Z(n65)
         );
  MUX2_X1 U134 ( .A(\CAM_MEM[0][1] ), .B(\CAM_MEM[8][1] ), .S(n365), .Z(n66)
         );
  MUX2_X1 U135 ( .A(n66), .B(n65), .S(n379), .Z(n67) );
  MUX2_X1 U136 ( .A(n67), .B(n64), .S(n388), .Z(n68) );
  MUX2_X1 U137 ( .A(n68), .B(n61), .S(n387), .Z(N607) );
  MUX2_X1 U138 ( .A(\CAM_MEM[7][2] ), .B(\CAM_MEM[15][2] ), .S(n365), .Z(n69)
         );
  MUX2_X1 U139 ( .A(\CAM_MEM[3][2] ), .B(\CAM_MEM[11][2] ), .S(n365), .Z(n70)
         );
  MUX2_X1 U140 ( .A(n70), .B(n69), .S(n379), .Z(n71) );
  MUX2_X1 U141 ( .A(\CAM_MEM[6][2] ), .B(\CAM_MEM[14][2] ), .S(n365), .Z(n72)
         );
  MUX2_X1 U142 ( .A(\CAM_MEM[2][2] ), .B(\CAM_MEM[10][2] ), .S(n365), .Z(n73)
         );
  MUX2_X1 U143 ( .A(n73), .B(n72), .S(n379), .Z(n74) );
  MUX2_X1 U144 ( .A(n74), .B(n71), .S(n388), .Z(n75) );
  MUX2_X1 U145 ( .A(\CAM_MEM[5][2] ), .B(\CAM_MEM[13][2] ), .S(n365), .Z(n76)
         );
  MUX2_X1 U146 ( .A(\CAM_MEM[1][2] ), .B(\CAM_MEM[9][2] ), .S(n365), .Z(n77)
         );
  MUX2_X1 U147 ( .A(n77), .B(n76), .S(n379), .Z(n78) );
  MUX2_X1 U148 ( .A(\CAM_MEM[4][2] ), .B(\CAM_MEM[12][2] ), .S(n365), .Z(n79)
         );
  MUX2_X1 U149 ( .A(\CAM_MEM[0][2] ), .B(\CAM_MEM[8][2] ), .S(n365), .Z(n80)
         );
  MUX2_X1 U150 ( .A(n80), .B(n79), .S(n379), .Z(n81) );
  MUX2_X1 U151 ( .A(n81), .B(n78), .S(n388), .Z(n82) );
  MUX2_X1 U152 ( .A(n82), .B(n75), .S(n387), .Z(N608) );
  MUX2_X1 U153 ( .A(\CAM_MEM[7][3] ), .B(\CAM_MEM[15][3] ), .S(n365), .Z(n83)
         );
  MUX2_X1 U154 ( .A(\CAM_MEM[3][3] ), .B(\CAM_MEM[11][3] ), .S(n365), .Z(n84)
         );
  MUX2_X1 U155 ( .A(n84), .B(n83), .S(n379), .Z(n85) );
  MUX2_X1 U156 ( .A(\CAM_MEM[6][3] ), .B(\CAM_MEM[14][3] ), .S(n365), .Z(n86)
         );
  MUX2_X1 U157 ( .A(\CAM_MEM[2][3] ), .B(\CAM_MEM[10][3] ), .S(n365), .Z(n87)
         );
  MUX2_X1 U158 ( .A(n87), .B(n86), .S(n379), .Z(n88) );
  MUX2_X1 U159 ( .A(n88), .B(n85), .S(n388), .Z(n89) );
  MUX2_X1 U160 ( .A(\CAM_MEM[5][3] ), .B(\CAM_MEM[13][3] ), .S(n366), .Z(n90)
         );
  MUX2_X1 U161 ( .A(\CAM_MEM[1][3] ), .B(\CAM_MEM[9][3] ), .S(n366), .Z(n91)
         );
  MUX2_X1 U162 ( .A(n91), .B(n90), .S(n380), .Z(n92) );
  MUX2_X1 U163 ( .A(\CAM_MEM[4][3] ), .B(\CAM_MEM[12][3] ), .S(n366), .Z(n93)
         );
  MUX2_X1 U164 ( .A(\CAM_MEM[0][3] ), .B(\CAM_MEM[8][3] ), .S(n366), .Z(n94)
         );
  MUX2_X1 U165 ( .A(n94), .B(n93), .S(n380), .Z(n95) );
  MUX2_X1 U166 ( .A(n95), .B(n92), .S(n389), .Z(n96) );
  MUX2_X1 U167 ( .A(n96), .B(n89), .S(n387), .Z(N609) );
  MUX2_X1 U168 ( .A(\CAM_MEM[7][4] ), .B(\CAM_MEM[15][4] ), .S(n366), .Z(n97)
         );
  MUX2_X1 U169 ( .A(\CAM_MEM[3][4] ), .B(\CAM_MEM[11][4] ), .S(n366), .Z(n98)
         );
  MUX2_X1 U170 ( .A(n98), .B(n97), .S(n380), .Z(n99) );
  MUX2_X1 U171 ( .A(\CAM_MEM[6][4] ), .B(\CAM_MEM[14][4] ), .S(n366), .Z(n100)
         );
  MUX2_X1 U172 ( .A(\CAM_MEM[2][4] ), .B(\CAM_MEM[10][4] ), .S(n366), .Z(n101)
         );
  MUX2_X1 U173 ( .A(n101), .B(n100), .S(n380), .Z(n102) );
  MUX2_X1 U174 ( .A(n102), .B(n99), .S(n389), .Z(n103) );
  MUX2_X1 U175 ( .A(\CAM_MEM[5][4] ), .B(\CAM_MEM[13][4] ), .S(n366), .Z(n104)
         );
  MUX2_X1 U176 ( .A(\CAM_MEM[1][4] ), .B(\CAM_MEM[9][4] ), .S(n366), .Z(n105)
         );
  MUX2_X1 U177 ( .A(n105), .B(n104), .S(n380), .Z(n106) );
  MUX2_X1 U178 ( .A(\CAM_MEM[4][4] ), .B(\CAM_MEM[12][4] ), .S(n366), .Z(n107)
         );
  MUX2_X1 U179 ( .A(\CAM_MEM[0][4] ), .B(\CAM_MEM[8][4] ), .S(n366), .Z(n108)
         );
  MUX2_X1 U180 ( .A(n108), .B(n107), .S(n380), .Z(n109) );
  MUX2_X1 U181 ( .A(n109), .B(n106), .S(n389), .Z(n110) );
  MUX2_X1 U182 ( .A(n110), .B(n103), .S(n387), .Z(N610) );
  MUX2_X1 U183 ( .A(\CAM_MEM[7][5] ), .B(\CAM_MEM[15][5] ), .S(n366), .Z(n111)
         );
  MUX2_X1 U184 ( .A(\CAM_MEM[3][5] ), .B(\CAM_MEM[11][5] ), .S(n367), .Z(n112)
         );
  MUX2_X1 U185 ( .A(n112), .B(n111), .S(n380), .Z(n113) );
  MUX2_X1 U186 ( .A(\CAM_MEM[6][5] ), .B(\CAM_MEM[14][5] ), .S(n367), .Z(n114)
         );
  MUX2_X1 U187 ( .A(\CAM_MEM[2][5] ), .B(\CAM_MEM[10][5] ), .S(n367), .Z(n115)
         );
  MUX2_X1 U188 ( .A(n115), .B(n114), .S(n380), .Z(n116) );
  MUX2_X1 U189 ( .A(n116), .B(n113), .S(n389), .Z(n117) );
  MUX2_X1 U190 ( .A(\CAM_MEM[5][5] ), .B(\CAM_MEM[13][5] ), .S(n367), .Z(n118)
         );
  MUX2_X1 U191 ( .A(\CAM_MEM[1][5] ), .B(\CAM_MEM[9][5] ), .S(n367), .Z(n119)
         );
  MUX2_X1 U192 ( .A(n119), .B(n118), .S(n380), .Z(n120) );
  MUX2_X1 U193 ( .A(\CAM_MEM[4][5] ), .B(\CAM_MEM[12][5] ), .S(n367), .Z(n121)
         );
  MUX2_X1 U194 ( .A(\CAM_MEM[0][5] ), .B(\CAM_MEM[8][5] ), .S(n367), .Z(n122)
         );
  MUX2_X1 U195 ( .A(n122), .B(n121), .S(n380), .Z(n123) );
  MUX2_X1 U196 ( .A(n123), .B(n120), .S(n389), .Z(n124) );
  MUX2_X1 U197 ( .A(n124), .B(n117), .S(n387), .Z(N611) );
  MUX2_X1 U198 ( .A(\CAM_MEM[7][6] ), .B(\CAM_MEM[15][6] ), .S(n367), .Z(n125)
         );
  MUX2_X1 U199 ( .A(\CAM_MEM[3][6] ), .B(\CAM_MEM[11][6] ), .S(n367), .Z(n126)
         );
  MUX2_X1 U200 ( .A(n126), .B(n125), .S(n380), .Z(n127) );
  MUX2_X1 U201 ( .A(\CAM_MEM[6][6] ), .B(\CAM_MEM[14][6] ), .S(n367), .Z(n128)
         );
  MUX2_X1 U202 ( .A(\CAM_MEM[2][6] ), .B(\CAM_MEM[10][6] ), .S(n367), .Z(n129)
         );
  MUX2_X1 U203 ( .A(n129), .B(n128), .S(n380), .Z(n130) );
  MUX2_X1 U204 ( .A(n130), .B(n127), .S(n389), .Z(n131) );
  MUX2_X1 U205 ( .A(\CAM_MEM[5][6] ), .B(\CAM_MEM[13][6] ), .S(n367), .Z(n132)
         );
  MUX2_X1 U206 ( .A(\CAM_MEM[1][6] ), .B(\CAM_MEM[9][6] ), .S(n367), .Z(n133)
         );
  MUX2_X1 U207 ( .A(n133), .B(n132), .S(n380), .Z(n134) );
  MUX2_X1 U208 ( .A(\CAM_MEM[4][6] ), .B(\CAM_MEM[12][6] ), .S(n368), .Z(n135)
         );
  MUX2_X1 U209 ( .A(\CAM_MEM[0][6] ), .B(\CAM_MEM[8][6] ), .S(n368), .Z(n136)
         );
  MUX2_X1 U210 ( .A(n136), .B(n135), .S(n381), .Z(n137) );
  MUX2_X1 U211 ( .A(n137), .B(n134), .S(n389), .Z(n138) );
  MUX2_X1 U212 ( .A(n138), .B(n131), .S(n387), .Z(N612) );
  MUX2_X1 U213 ( .A(\CAM_MEM[7][7] ), .B(\CAM_MEM[15][7] ), .S(n368), .Z(n139)
         );
  MUX2_X1 U214 ( .A(\CAM_MEM[3][7] ), .B(\CAM_MEM[11][7] ), .S(n368), .Z(n140)
         );
  MUX2_X1 U215 ( .A(n140), .B(n139), .S(n381), .Z(n141) );
  MUX2_X1 U216 ( .A(\CAM_MEM[6][7] ), .B(\CAM_MEM[14][7] ), .S(n368), .Z(n142)
         );
  MUX2_X1 U217 ( .A(\CAM_MEM[2][7] ), .B(\CAM_MEM[10][7] ), .S(n368), .Z(n143)
         );
  MUX2_X1 U218 ( .A(n143), .B(n142), .S(n381), .Z(n144) );
  MUX2_X1 U219 ( .A(n144), .B(n141), .S(n389), .Z(n145) );
  MUX2_X1 U220 ( .A(\CAM_MEM[5][7] ), .B(\CAM_MEM[13][7] ), .S(n368), .Z(n146)
         );
  MUX2_X1 U221 ( .A(\CAM_MEM[1][7] ), .B(\CAM_MEM[9][7] ), .S(n368), .Z(n147)
         );
  MUX2_X1 U222 ( .A(n147), .B(n146), .S(n381), .Z(n148) );
  MUX2_X1 U223 ( .A(\CAM_MEM[4][7] ), .B(\CAM_MEM[12][7] ), .S(n368), .Z(n149)
         );
  MUX2_X1 U224 ( .A(\CAM_MEM[0][7] ), .B(\CAM_MEM[8][7] ), .S(n368), .Z(n150)
         );
  MUX2_X1 U225 ( .A(n150), .B(n149), .S(n381), .Z(n151) );
  MUX2_X1 U226 ( .A(n151), .B(n148), .S(n389), .Z(n152) );
  MUX2_X1 U227 ( .A(n152), .B(n145), .S(n387), .Z(N613) );
  MUX2_X1 U228 ( .A(\CAM_MEM[7][8] ), .B(\CAM_MEM[15][8] ), .S(n368), .Z(n153)
         );
  MUX2_X1 U229 ( .A(\CAM_MEM[3][8] ), .B(\CAM_MEM[11][8] ), .S(n368), .Z(n154)
         );
  MUX2_X1 U230 ( .A(n154), .B(n153), .S(n381), .Z(n155) );
  MUX2_X1 U231 ( .A(\CAM_MEM[6][8] ), .B(\CAM_MEM[14][8] ), .S(n368), .Z(n156)
         );
  MUX2_X1 U232 ( .A(\CAM_MEM[2][8] ), .B(\CAM_MEM[10][8] ), .S(n369), .Z(n157)
         );
  MUX2_X1 U233 ( .A(n157), .B(n156), .S(n381), .Z(n158) );
  MUX2_X1 U234 ( .A(n158), .B(n155), .S(n389), .Z(n159) );
  MUX2_X1 U235 ( .A(\CAM_MEM[5][8] ), .B(\CAM_MEM[13][8] ), .S(n369), .Z(n160)
         );
  MUX2_X1 U236 ( .A(\CAM_MEM[1][8] ), .B(\CAM_MEM[9][8] ), .S(n369), .Z(n161)
         );
  MUX2_X1 U237 ( .A(n161), .B(n160), .S(n381), .Z(n162) );
  MUX2_X1 U238 ( .A(\CAM_MEM[4][8] ), .B(\CAM_MEM[12][8] ), .S(n369), .Z(n163)
         );
  MUX2_X1 U239 ( .A(\CAM_MEM[0][8] ), .B(\CAM_MEM[8][8] ), .S(n369), .Z(n164)
         );
  MUX2_X1 U240 ( .A(n164), .B(n163), .S(n381), .Z(n165) );
  MUX2_X1 U241 ( .A(n165), .B(n162), .S(n389), .Z(n166) );
  MUX2_X1 U242 ( .A(n166), .B(n159), .S(n387), .Z(N614) );
  MUX2_X1 U243 ( .A(\CAM_MEM[7][9] ), .B(\CAM_MEM[15][9] ), .S(n369), .Z(n167)
         );
  MUX2_X1 U244 ( .A(\CAM_MEM[3][9] ), .B(\CAM_MEM[11][9] ), .S(n369), .Z(n168)
         );
  MUX2_X1 U245 ( .A(n168), .B(n167), .S(n381), .Z(n169) );
  MUX2_X1 U246 ( .A(\CAM_MEM[6][9] ), .B(\CAM_MEM[14][9] ), .S(n369), .Z(n170)
         );
  MUX2_X1 U247 ( .A(\CAM_MEM[2][9] ), .B(\CAM_MEM[10][9] ), .S(n369), .Z(n171)
         );
  MUX2_X1 U248 ( .A(n171), .B(n170), .S(n381), .Z(n172) );
  MUX2_X1 U249 ( .A(n172), .B(n169), .S(n389), .Z(n173) );
  MUX2_X1 U250 ( .A(\CAM_MEM[5][9] ), .B(\CAM_MEM[13][9] ), .S(n369), .Z(n174)
         );
  MUX2_X1 U251 ( .A(\CAM_MEM[1][9] ), .B(\CAM_MEM[9][9] ), .S(n369), .Z(n175)
         );
  MUX2_X1 U252 ( .A(n175), .B(n174), .S(n381), .Z(n176) );
  MUX2_X1 U253 ( .A(\CAM_MEM[4][9] ), .B(\CAM_MEM[12][9] ), .S(n369), .Z(n177)
         );
  MUX2_X1 U254 ( .A(\CAM_MEM[0][9] ), .B(\CAM_MEM[8][9] ), .S(n369), .Z(n178)
         );
  MUX2_X1 U255 ( .A(n178), .B(n177), .S(n381), .Z(n179) );
  MUX2_X1 U256 ( .A(n179), .B(n176), .S(n389), .Z(n180) );
  MUX2_X1 U257 ( .A(n180), .B(n173), .S(n387), .Z(N615) );
  MUX2_X1 U258 ( .A(\CAM_MEM[7][10] ), .B(\CAM_MEM[15][10] ), .S(n370), .Z(
        n181) );
  MUX2_X1 U259 ( .A(\CAM_MEM[3][10] ), .B(\CAM_MEM[11][10] ), .S(n370), .Z(
        n182) );
  MUX2_X1 U260 ( .A(n182), .B(n181), .S(n382), .Z(n183) );
  MUX2_X1 U261 ( .A(\CAM_MEM[6][10] ), .B(\CAM_MEM[14][10] ), .S(n370), .Z(
        n184) );
  MUX2_X1 U262 ( .A(\CAM_MEM[2][10] ), .B(\CAM_MEM[10][10] ), .S(n370), .Z(
        n185) );
  MUX2_X1 U263 ( .A(n185), .B(n184), .S(n382), .Z(n186) );
  MUX2_X1 U264 ( .A(n186), .B(n183), .S(n390), .Z(n187) );
  MUX2_X1 U265 ( .A(\CAM_MEM[5][10] ), .B(\CAM_MEM[13][10] ), .S(n370), .Z(
        n188) );
  MUX2_X1 U266 ( .A(\CAM_MEM[1][10] ), .B(\CAM_MEM[9][10] ), .S(n370), .Z(n189) );
  MUX2_X1 U267 ( .A(n189), .B(n188), .S(n382), .Z(n190) );
  MUX2_X1 U268 ( .A(\CAM_MEM[4][10] ), .B(\CAM_MEM[12][10] ), .S(n370), .Z(
        n191) );
  MUX2_X1 U269 ( .A(\CAM_MEM[0][10] ), .B(\CAM_MEM[8][10] ), .S(n370), .Z(n192) );
  MUX2_X1 U270 ( .A(n192), .B(n191), .S(n382), .Z(n193) );
  MUX2_X1 U271 ( .A(n193), .B(n190), .S(n390), .Z(n194) );
  MUX2_X1 U272 ( .A(n194), .B(n187), .S(n387), .Z(N616) );
  MUX2_X1 U273 ( .A(\CAM_MEM[7][11] ), .B(\CAM_MEM[15][11] ), .S(n370), .Z(
        n195) );
  MUX2_X1 U274 ( .A(\CAM_MEM[3][11] ), .B(\CAM_MEM[11][11] ), .S(n370), .Z(
        n196) );
  MUX2_X1 U275 ( .A(n196), .B(n195), .S(n382), .Z(n197) );
  MUX2_X1 U276 ( .A(\CAM_MEM[6][11] ), .B(\CAM_MEM[14][11] ), .S(n370), .Z(
        n198) );
  MUX2_X1 U277 ( .A(\CAM_MEM[2][11] ), .B(\CAM_MEM[10][11] ), .S(n370), .Z(
        n199) );
  MUX2_X1 U278 ( .A(n199), .B(n198), .S(n382), .Z(n200) );
  MUX2_X1 U279 ( .A(n200), .B(n197), .S(n390), .Z(n201) );
  MUX2_X1 U280 ( .A(\CAM_MEM[5][11] ), .B(\CAM_MEM[13][11] ), .S(n370), .Z(
        n202) );
  MUX2_X1 U281 ( .A(\CAM_MEM[1][11] ), .B(\CAM_MEM[9][11] ), .S(n371), .Z(n203) );
  MUX2_X1 U282 ( .A(n203), .B(n202), .S(n382), .Z(n204) );
  MUX2_X1 U283 ( .A(\CAM_MEM[4][11] ), .B(\CAM_MEM[12][11] ), .S(n371), .Z(
        n205) );
  MUX2_X1 U284 ( .A(\CAM_MEM[0][11] ), .B(\CAM_MEM[8][11] ), .S(n371), .Z(n206) );
  MUX2_X1 U285 ( .A(n206), .B(n205), .S(n382), .Z(n207) );
  MUX2_X1 U286 ( .A(n207), .B(n204), .S(n390), .Z(n208) );
  MUX2_X1 U287 ( .A(n208), .B(n201), .S(n387), .Z(N617) );
  MUX2_X1 U288 ( .A(\CAM_MEM[7][12] ), .B(\CAM_MEM[15][12] ), .S(n371), .Z(
        n209) );
  MUX2_X1 U289 ( .A(\CAM_MEM[3][12] ), .B(\CAM_MEM[11][12] ), .S(n371), .Z(
        n210) );
  MUX2_X1 U290 ( .A(n210), .B(n209), .S(n382), .Z(n211) );
  MUX2_X1 U291 ( .A(\CAM_MEM[6][12] ), .B(\CAM_MEM[14][12] ), .S(n371), .Z(
        n212) );
  MUX2_X1 U292 ( .A(\CAM_MEM[2][12] ), .B(\CAM_MEM[10][12] ), .S(n371), .Z(
        n213) );
  MUX2_X1 U293 ( .A(n213), .B(n212), .S(n382), .Z(n214) );
  MUX2_X1 U294 ( .A(n214), .B(n211), .S(n390), .Z(n215) );
  MUX2_X1 U295 ( .A(\CAM_MEM[5][12] ), .B(\CAM_MEM[13][12] ), .S(n371), .Z(
        n216) );
  MUX2_X1 U296 ( .A(\CAM_MEM[1][12] ), .B(\CAM_MEM[9][12] ), .S(n371), .Z(n217) );
  MUX2_X1 U297 ( .A(n217), .B(n216), .S(n382), .Z(n218) );
  MUX2_X1 U298 ( .A(\CAM_MEM[4][12] ), .B(\CAM_MEM[12][12] ), .S(n371), .Z(
        n219) );
  MUX2_X1 U299 ( .A(\CAM_MEM[0][12] ), .B(\CAM_MEM[8][12] ), .S(n371), .Z(n220) );
  MUX2_X1 U300 ( .A(n220), .B(n219), .S(n382), .Z(n221) );
  MUX2_X1 U301 ( .A(n221), .B(n218), .S(n390), .Z(n222) );
  MUX2_X1 U302 ( .A(n222), .B(n215), .S(n386), .Z(N618) );
  MUX2_X1 U303 ( .A(\CAM_MEM[7][13] ), .B(\CAM_MEM[15][13] ), .S(n371), .Z(
        n223) );
  MUX2_X1 U304 ( .A(\CAM_MEM[3][13] ), .B(\CAM_MEM[11][13] ), .S(n371), .Z(
        n224) );
  MUX2_X1 U305 ( .A(n224), .B(n223), .S(n382), .Z(n225) );
  MUX2_X1 U306 ( .A(\CAM_MEM[6][13] ), .B(\CAM_MEM[14][13] ), .S(n372), .Z(
        n226) );
  MUX2_X1 U307 ( .A(\CAM_MEM[2][13] ), .B(\CAM_MEM[10][13] ), .S(n372), .Z(
        n227) );
  MUX2_X1 U308 ( .A(n227), .B(n226), .S(n383), .Z(n228) );
  MUX2_X1 U309 ( .A(n228), .B(n225), .S(n390), .Z(n229) );
  MUX2_X1 U310 ( .A(\CAM_MEM[5][13] ), .B(\CAM_MEM[13][13] ), .S(n372), .Z(
        n230) );
  MUX2_X1 U311 ( .A(\CAM_MEM[1][13] ), .B(\CAM_MEM[9][13] ), .S(n372), .Z(n231) );
  MUX2_X1 U312 ( .A(n231), .B(n230), .S(n383), .Z(n232) );
  MUX2_X1 U313 ( .A(\CAM_MEM[4][13] ), .B(\CAM_MEM[12][13] ), .S(n372), .Z(
        n233) );
  MUX2_X1 U314 ( .A(\CAM_MEM[0][13] ), .B(\CAM_MEM[8][13] ), .S(n372), .Z(n234) );
  MUX2_X1 U315 ( .A(n234), .B(n233), .S(n383), .Z(n235) );
  MUX2_X1 U316 ( .A(n235), .B(n232), .S(n390), .Z(n236) );
  MUX2_X1 U317 ( .A(n236), .B(n229), .S(n386), .Z(N619) );
  MUX2_X1 U318 ( .A(\CAM_MEM[7][14] ), .B(\CAM_MEM[15][14] ), .S(n372), .Z(
        n237) );
  MUX2_X1 U319 ( .A(\CAM_MEM[3][14] ), .B(\CAM_MEM[11][14] ), .S(n372), .Z(
        n238) );
  MUX2_X1 U320 ( .A(n238), .B(n237), .S(n383), .Z(n239) );
  MUX2_X1 U321 ( .A(\CAM_MEM[6][14] ), .B(\CAM_MEM[14][14] ), .S(n372), .Z(
        n240) );
  MUX2_X1 U322 ( .A(\CAM_MEM[2][14] ), .B(\CAM_MEM[10][14] ), .S(n372), .Z(
        n241) );
  MUX2_X1 U323 ( .A(n241), .B(n240), .S(n383), .Z(n242) );
  MUX2_X1 U324 ( .A(n242), .B(n239), .S(n390), .Z(n243) );
  MUX2_X1 U325 ( .A(\CAM_MEM[5][14] ), .B(\CAM_MEM[13][14] ), .S(n372), .Z(
        n244) );
  MUX2_X1 U326 ( .A(\CAM_MEM[1][14] ), .B(\CAM_MEM[9][14] ), .S(n372), .Z(n245) );
  MUX2_X1 U327 ( .A(n245), .B(n244), .S(n383), .Z(n246) );
  MUX2_X1 U328 ( .A(\CAM_MEM[4][14] ), .B(\CAM_MEM[12][14] ), .S(n372), .Z(
        n247) );
  MUX2_X1 U329 ( .A(\CAM_MEM[0][14] ), .B(\CAM_MEM[8][14] ), .S(n373), .Z(n248) );
  MUX2_X1 U330 ( .A(n248), .B(n247), .S(n383), .Z(n249) );
  MUX2_X1 U331 ( .A(n249), .B(n246), .S(n390), .Z(n250) );
  MUX2_X1 U332 ( .A(n250), .B(n243), .S(n386), .Z(N620) );
  MUX2_X1 U333 ( .A(\CAM_MEM[7][15] ), .B(\CAM_MEM[15][15] ), .S(n373), .Z(
        n251) );
  MUX2_X1 U334 ( .A(\CAM_MEM[3][15] ), .B(\CAM_MEM[11][15] ), .S(n373), .Z(
        n252) );
  MUX2_X1 U335 ( .A(n252), .B(n251), .S(n383), .Z(n253) );
  MUX2_X1 U336 ( .A(\CAM_MEM[6][15] ), .B(\CAM_MEM[14][15] ), .S(n373), .Z(
        n254) );
  MUX2_X1 U337 ( .A(\CAM_MEM[2][15] ), .B(\CAM_MEM[10][15] ), .S(n373), .Z(
        n255) );
  MUX2_X1 U338 ( .A(n255), .B(n254), .S(n383), .Z(n256) );
  MUX2_X1 U339 ( .A(n256), .B(n253), .S(n390), .Z(n257) );
  MUX2_X1 U340 ( .A(\CAM_MEM[5][15] ), .B(\CAM_MEM[13][15] ), .S(n373), .Z(
        n258) );
  MUX2_X1 U341 ( .A(\CAM_MEM[1][15] ), .B(\CAM_MEM[9][15] ), .S(n373), .Z(n259) );
  MUX2_X1 U342 ( .A(n259), .B(n258), .S(n383), .Z(n260) );
  MUX2_X1 U343 ( .A(\CAM_MEM[4][15] ), .B(\CAM_MEM[12][15] ), .S(n373), .Z(
        n261) );
  MUX2_X1 U344 ( .A(\CAM_MEM[0][15] ), .B(\CAM_MEM[8][15] ), .S(n373), .Z(n262) );
  MUX2_X1 U345 ( .A(n262), .B(n261), .S(n383), .Z(n263) );
  MUX2_X1 U346 ( .A(n263), .B(n260), .S(n390), .Z(n264) );
  MUX2_X1 U347 ( .A(n264), .B(n257), .S(n386), .Z(N621) );
  MUX2_X1 U348 ( .A(\CAM_MEM[7][16] ), .B(\CAM_MEM[15][16] ), .S(n373), .Z(
        n265) );
  MUX2_X1 U349 ( .A(\CAM_MEM[3][16] ), .B(\CAM_MEM[11][16] ), .S(n373), .Z(
        n266) );
  MUX2_X1 U350 ( .A(n266), .B(n265), .S(n383), .Z(n267) );
  MUX2_X1 U351 ( .A(\CAM_MEM[6][16] ), .B(\CAM_MEM[14][16] ), .S(n373), .Z(
        n268) );
  MUX2_X1 U352 ( .A(\CAM_MEM[2][16] ), .B(\CAM_MEM[10][16] ), .S(n373), .Z(
        n269) );
  MUX2_X1 U353 ( .A(n269), .B(n268), .S(n383), .Z(n270) );
  MUX2_X1 U354 ( .A(n270), .B(n267), .S(n390), .Z(n271) );
  MUX2_X1 U355 ( .A(\CAM_MEM[5][16] ), .B(\CAM_MEM[13][16] ), .S(n374), .Z(
        n272) );
  MUX2_X1 U356 ( .A(\CAM_MEM[1][16] ), .B(\CAM_MEM[9][16] ), .S(n374), .Z(n273) );
  MUX2_X1 U357 ( .A(n273), .B(n272), .S(n384), .Z(n274) );
  MUX2_X1 U358 ( .A(\CAM_MEM[4][16] ), .B(\CAM_MEM[12][16] ), .S(n374), .Z(
        n275) );
  MUX2_X1 U359 ( .A(\CAM_MEM[0][16] ), .B(\CAM_MEM[8][16] ), .S(n374), .Z(n276) );
  MUX2_X1 U360 ( .A(n276), .B(n275), .S(n384), .Z(n277) );
  MUX2_X1 U361 ( .A(n277), .B(n274), .S(n391), .Z(n278) );
  MUX2_X1 U362 ( .A(n278), .B(n271), .S(n386), .Z(N622) );
  MUX2_X1 U363 ( .A(\CAM_MEM[7][17] ), .B(\CAM_MEM[15][17] ), .S(n374), .Z(
        n279) );
  MUX2_X1 U364 ( .A(\CAM_MEM[3][17] ), .B(\CAM_MEM[11][17] ), .S(n374), .Z(
        n280) );
  MUX2_X1 U365 ( .A(n280), .B(n279), .S(n384), .Z(n281) );
  MUX2_X1 U366 ( .A(\CAM_MEM[6][17] ), .B(\CAM_MEM[14][17] ), .S(n374), .Z(
        n282) );
  MUX2_X1 U367 ( .A(\CAM_MEM[2][17] ), .B(\CAM_MEM[10][17] ), .S(n374), .Z(
        n283) );
  MUX2_X1 U368 ( .A(n283), .B(n282), .S(n384), .Z(n284) );
  MUX2_X1 U369 ( .A(n284), .B(n281), .S(n391), .Z(n285) );
  MUX2_X1 U370 ( .A(\CAM_MEM[5][17] ), .B(\CAM_MEM[13][17] ), .S(n374), .Z(
        n286) );
  MUX2_X1 U371 ( .A(\CAM_MEM[1][17] ), .B(\CAM_MEM[9][17] ), .S(n374), .Z(n287) );
  MUX2_X1 U372 ( .A(n287), .B(n286), .S(n384), .Z(n288) );
  MUX2_X1 U373 ( .A(\CAM_MEM[4][17] ), .B(\CAM_MEM[12][17] ), .S(n374), .Z(
        n289) );
  MUX2_X1 U374 ( .A(\CAM_MEM[0][17] ), .B(\CAM_MEM[8][17] ), .S(n374), .Z(n290) );
  MUX2_X1 U375 ( .A(n290), .B(n289), .S(n384), .Z(n291) );
  MUX2_X1 U376 ( .A(n291), .B(n288), .S(n391), .Z(n292) );
  MUX2_X1 U377 ( .A(n292), .B(n285), .S(n386), .Z(N623) );
  MUX2_X1 U378 ( .A(\CAM_MEM[7][18] ), .B(\CAM_MEM[15][18] ), .S(n374), .Z(
        n293) );
  MUX2_X1 U379 ( .A(\CAM_MEM[3][18] ), .B(\CAM_MEM[11][18] ), .S(n375), .Z(
        n294) );
  MUX2_X1 U380 ( .A(n294), .B(n293), .S(n384), .Z(n295) );
  MUX2_X1 U381 ( .A(\CAM_MEM[6][18] ), .B(\CAM_MEM[14][18] ), .S(n375), .Z(
        n296) );
  MUX2_X1 U382 ( .A(\CAM_MEM[2][18] ), .B(\CAM_MEM[10][18] ), .S(n375), .Z(
        n297) );
  MUX2_X1 U383 ( .A(n297), .B(n296), .S(n384), .Z(n298) );
  MUX2_X1 U384 ( .A(n298), .B(n295), .S(n391), .Z(n299) );
  MUX2_X1 U385 ( .A(\CAM_MEM[5][18] ), .B(\CAM_MEM[13][18] ), .S(n375), .Z(
        n300) );
  MUX2_X1 U386 ( .A(\CAM_MEM[1][18] ), .B(\CAM_MEM[9][18] ), .S(n375), .Z(n301) );
  MUX2_X1 U387 ( .A(n301), .B(n300), .S(n384), .Z(n302) );
  MUX2_X1 U388 ( .A(\CAM_MEM[4][18] ), .B(\CAM_MEM[12][18] ), .S(n375), .Z(
        n303) );
  MUX2_X1 U389 ( .A(\CAM_MEM[0][18] ), .B(\CAM_MEM[8][18] ), .S(n375), .Z(n304) );
  MUX2_X1 U390 ( .A(n304), .B(n303), .S(n384), .Z(n305) );
  MUX2_X1 U391 ( .A(n305), .B(n302), .S(n391), .Z(n306) );
  MUX2_X1 U392 ( .A(n306), .B(n299), .S(n386), .Z(N624) );
  MUX2_X1 U393 ( .A(\CAM_MEM[7][19] ), .B(\CAM_MEM[15][19] ), .S(n375), .Z(
        n307) );
  MUX2_X1 U394 ( .A(\CAM_MEM[3][19] ), .B(\CAM_MEM[11][19] ), .S(n375), .Z(
        n308) );
  MUX2_X1 U395 ( .A(n308), .B(n307), .S(n384), .Z(n309) );
  MUX2_X1 U396 ( .A(\CAM_MEM[6][19] ), .B(\CAM_MEM[14][19] ), .S(n375), .Z(
        n310) );
  MUX2_X1 U397 ( .A(\CAM_MEM[2][19] ), .B(\CAM_MEM[10][19] ), .S(n375), .Z(
        n311) );
  MUX2_X1 U398 ( .A(n311), .B(n310), .S(n384), .Z(n312) );
  MUX2_X1 U399 ( .A(n312), .B(n309), .S(n391), .Z(n313) );
  MUX2_X1 U400 ( .A(\CAM_MEM[5][19] ), .B(\CAM_MEM[13][19] ), .S(n375), .Z(
        n314) );
  MUX2_X1 U401 ( .A(\CAM_MEM[1][19] ), .B(\CAM_MEM[9][19] ), .S(n375), .Z(n315) );
  MUX2_X1 U402 ( .A(n315), .B(n314), .S(n384), .Z(n316) );
  MUX2_X1 U403 ( .A(\CAM_MEM[4][19] ), .B(\CAM_MEM[12][19] ), .S(n376), .Z(
        n317) );
  MUX2_X1 U404 ( .A(\CAM_MEM[0][19] ), .B(\CAM_MEM[8][19] ), .S(n376), .Z(n318) );
  MUX2_X1 U405 ( .A(n318), .B(n317), .S(n385), .Z(n319) );
  MUX2_X1 U406 ( .A(n319), .B(n316), .S(n391), .Z(n320) );
  MUX2_X1 U407 ( .A(n320), .B(n313), .S(n386), .Z(N625) );
  MUX2_X1 U408 ( .A(\CAM_MEM[7][20] ), .B(\CAM_MEM[15][20] ), .S(n376), .Z(
        n321) );
  MUX2_X1 U409 ( .A(\CAM_MEM[3][20] ), .B(\CAM_MEM[11][20] ), .S(n376), .Z(
        n322) );
  MUX2_X1 U410 ( .A(n322), .B(n321), .S(n385), .Z(n323) );
  MUX2_X1 U411 ( .A(\CAM_MEM[6][20] ), .B(\CAM_MEM[14][20] ), .S(n376), .Z(
        n324) );
  MUX2_X1 U412 ( .A(\CAM_MEM[2][20] ), .B(\CAM_MEM[10][20] ), .S(n376), .Z(
        n325) );
  MUX2_X1 U413 ( .A(n325), .B(n324), .S(n385), .Z(n326) );
  MUX2_X1 U414 ( .A(n326), .B(n323), .S(n391), .Z(n327) );
  MUX2_X1 U415 ( .A(\CAM_MEM[5][20] ), .B(\CAM_MEM[13][20] ), .S(n376), .Z(
        n328) );
  MUX2_X1 U416 ( .A(\CAM_MEM[1][20] ), .B(\CAM_MEM[9][20] ), .S(n376), .Z(n329) );
  MUX2_X1 U417 ( .A(n329), .B(n328), .S(n385), .Z(n330) );
  MUX2_X1 U418 ( .A(\CAM_MEM[4][20] ), .B(\CAM_MEM[12][20] ), .S(n376), .Z(
        n331) );
  MUX2_X1 U419 ( .A(\CAM_MEM[0][20] ), .B(\CAM_MEM[8][20] ), .S(n376), .Z(n332) );
  MUX2_X1 U420 ( .A(n332), .B(n331), .S(n385), .Z(n333) );
  MUX2_X1 U421 ( .A(n333), .B(n330), .S(n391), .Z(n334) );
  MUX2_X1 U422 ( .A(n334), .B(n327), .S(n386), .Z(N626) );
  MUX2_X1 U423 ( .A(\CAM_MEM[7][21] ), .B(\CAM_MEM[15][21] ), .S(n376), .Z(
        n335) );
  MUX2_X1 U424 ( .A(\CAM_MEM[3][21] ), .B(\CAM_MEM[11][21] ), .S(n376), .Z(
        n336) );
  MUX2_X1 U425 ( .A(n336), .B(n335), .S(n385), .Z(n337) );
  MUX2_X1 U426 ( .A(\CAM_MEM[6][21] ), .B(\CAM_MEM[14][21] ), .S(n376), .Z(
        n338) );
  MUX2_X1 U427 ( .A(\CAM_MEM[2][21] ), .B(\CAM_MEM[10][21] ), .S(n377), .Z(
        n339) );
  MUX2_X1 U428 ( .A(n339), .B(n338), .S(n385), .Z(n340) );
  MUX2_X1 U429 ( .A(n340), .B(n337), .S(n391), .Z(n341) );
  MUX2_X1 U430 ( .A(\CAM_MEM[5][21] ), .B(\CAM_MEM[13][21] ), .S(n377), .Z(
        n342) );
  MUX2_X1 U431 ( .A(\CAM_MEM[1][21] ), .B(\CAM_MEM[9][21] ), .S(n377), .Z(n343) );
  MUX2_X1 U432 ( .A(n343), .B(n342), .S(n385), .Z(n344) );
  MUX2_X1 U433 ( .A(\CAM_MEM[4][21] ), .B(\CAM_MEM[12][21] ), .S(n377), .Z(
        n345) );
  MUX2_X1 U434 ( .A(\CAM_MEM[0][21] ), .B(\CAM_MEM[8][21] ), .S(n377), .Z(n346) );
  MUX2_X1 U435 ( .A(n346), .B(n345), .S(n385), .Z(n347) );
  MUX2_X1 U436 ( .A(n347), .B(n344), .S(n391), .Z(n348) );
  MUX2_X1 U437 ( .A(n348), .B(n341), .S(n386), .Z(N627) );
  MUX2_X1 U438 ( .A(\CAM_MEM[7][22] ), .B(\CAM_MEM[15][22] ), .S(n377), .Z(
        n349) );
  MUX2_X1 U439 ( .A(\CAM_MEM[3][22] ), .B(\CAM_MEM[11][22] ), .S(n377), .Z(
        n350) );
  MUX2_X1 U440 ( .A(n350), .B(n349), .S(n385), .Z(n351) );
  MUX2_X1 U441 ( .A(\CAM_MEM[6][22] ), .B(\CAM_MEM[14][22] ), .S(n377), .Z(
        n352) );
  MUX2_X1 U442 ( .A(\CAM_MEM[2][22] ), .B(\CAM_MEM[10][22] ), .S(n377), .Z(
        n353) );
  MUX2_X1 U443 ( .A(n353), .B(n352), .S(n385), .Z(n354) );
  MUX2_X1 U444 ( .A(n354), .B(n351), .S(n391), .Z(n355) );
  MUX2_X1 U445 ( .A(\CAM_MEM[5][22] ), .B(\CAM_MEM[13][22] ), .S(n377), .Z(
        n356) );
  MUX2_X1 U446 ( .A(\CAM_MEM[1][22] ), .B(\CAM_MEM[9][22] ), .S(n377), .Z(n357) );
  MUX2_X1 U447 ( .A(n357), .B(n356), .S(n385), .Z(n358) );
  MUX2_X1 U448 ( .A(\CAM_MEM[4][22] ), .B(\CAM_MEM[12][22] ), .S(n377), .Z(
        n359) );
  MUX2_X1 U449 ( .A(\CAM_MEM[0][22] ), .B(\CAM_MEM[8][22] ), .S(n377), .Z(n360) );
  MUX2_X1 U450 ( .A(n360), .B(n359), .S(n385), .Z(n361) );
  MUX2_X1 U451 ( .A(n361), .B(n358), .S(n391), .Z(n362) );
  MUX2_X1 U452 ( .A(n362), .B(n355), .S(n386), .Z(N628) );
  CLKBUF_X1 U453 ( .A(SET_INDEX[2]), .Z(n378) );
  INV_X1 U454 ( .A(SET_INDEX[1]), .ZN(n393) );
  INV_X1 U455 ( .A(SET_INDEX[2]), .ZN(n394) );
  INV_X1 U456 ( .A(SET_INDEX[3]), .ZN(n395) );
endmodule


module MUX21_GEN_N5 ( A, B, SEL, Y );
  input [4:0] A;
  input [4:0] B;
  output [4:0] Y;
  input SEL;
  wire   SB;
  wire   [4:0] Y1;
  wire   [4:0] Y2;

  INV_1_122 UIV ( .A(SEL), .Y(SB) );
  NAND_GATE_1134 UND1_0 ( .A(A[0]), .B(SEL), .Y(Y1[0]) );
  NAND_GATE_1133 UND2_0 ( .A(B[0]), .B(SB), .Y(Y2[0]) );
  NAND_GATE_1132 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_1131 UND1_1 ( .A(A[1]), .B(SEL), .Y(Y1[1]) );
  NAND_GATE_1130 UND2_1 ( .A(B[1]), .B(SB), .Y(Y2[1]) );
  NAND_GATE_1129 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_1128 UND1_2 ( .A(A[2]), .B(SEL), .Y(Y1[2]) );
  NAND_GATE_1127 UND2_2 ( .A(B[2]), .B(SB), .Y(Y2[2]) );
  NAND_GATE_1126 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_1125 UND1_3 ( .A(A[3]), .B(SEL), .Y(Y1[3]) );
  NAND_GATE_1124 UND2_3 ( .A(B[3]), .B(SB), .Y(Y2[3]) );
  NAND_GATE_1123 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_1122 UND1_4 ( .A(A[4]), .B(SEL), .Y(Y1[4]) );
  NAND_GATE_1121 UND2_4 ( .A(B[4]), .B(SB), .Y(Y2[4]) );
  NAND_GATE_1120 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
endmodule


module FORW_FSM_OPCODE_SIZE6_N_ADDR5 ( CLK, RST, CMP_A_EXE, CMP_A_MEM, 
        CMP_B_EXE, CMP_B_MEM, CMP_C_EXE, CMP_C_MEM, CMP_BRANCH_ID, 
        CMP_BRANCH_EXE, CMP_BRANCH_MEM, OPCODE_IF, OPCODE_ID, OPCODE_EXE, 
        OPCODE_MEM, OPCODE_WB, MUX_A, MUX_B, MUX_C, MUX_D, RST_DIV, 
        STALL_BRANCH, STALL );
  input [5:0] OPCODE_IF;
  input [5:0] OPCODE_ID;
  input [5:0] OPCODE_EXE;
  input [5:0] OPCODE_MEM;
  input [5:0] OPCODE_WB;
  output [1:0] MUX_A;
  output [1:0] MUX_B;
  output [1:0] MUX_C;
  output [1:0] MUX_D;
  input CLK, RST, CMP_A_EXE, CMP_A_MEM, CMP_B_EXE, CMP_B_MEM, CMP_C_EXE,
         CMP_C_MEM, CMP_BRANCH_ID, CMP_BRANCH_EXE, CMP_BRANCH_MEM;
  output RST_DIV, STALL_BRANCH, STALL;
  wire   N341, N342, N380, N381, N382, N438, N439, N440, N458, N459,
         \CURRENT_STATE_D[1] , N508, N509, N510, N511, N512, N513, N514, N515,
         N516, N517, N518, N519, N520, N521, N522, N523, N524, N525, N526,
         N527, N528, N529, N530, N531, N532, N533, N534, N535, N536, N537,
         N538, N539, N578, N579, N580, N581, N582, N583, N584, N585, N586,
         N587, N588, N589, N590, N591, N592, N593, N594, N595, N596, N597,
         N598, N599, N600, N601, N602, N603, N604, N605, N606, N607, N608,
         N609, n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n106,
         n108, n110, n112, n114, n115, n116, n118, n120, n121, n122, n123,
         n124, n125, n127, n129, n131, n133, n135, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n237, n238, n239, n240, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n256, n257, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n341, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n56, n66, n97, n105, n107, n109, n111, n113, n117,
         n119, n126, n128, n130, n132, n134, n136, n210, n211, n235, n236,
         n241, n242, n243, n254, n255, n258, n259, n260, n261, n289;
  wire   [31:0] CNT_MUL;
  wire   [31:0] CNT_DIV;

  DFFR_X1 \CURRENT_STATE_C_reg[1]  ( .D(N459), .CK(CLK), .RN(n40), .QN(
        MUX_C[1]) );
  DFFR_X1 \CURRENT_STATE_C_reg[0]  ( .D(N458), .CK(CLK), .RN(n38), .QN(
        MUX_C[0]) );
  DFFR_X1 \CNT_DIV_reg[0]  ( .D(n441), .CK(CLK), .RN(n38), .Q(CNT_DIV[0]), 
        .QN(n468) );
  DFFR_X1 \CNT_DIV_reg[10]  ( .D(n440), .CK(CLK), .RN(n38), .Q(CNT_DIV[10]), 
        .QN(n448) );
  DFFR_X1 \CNT_DIV_reg[31]  ( .D(n439), .CK(CLK), .RN(n38), .Q(CNT_DIV[31]), 
        .QN(n461) );
  DFFR_X1 \CNT_MUL_reg[30]  ( .D(n438), .CK(CLK), .RN(n38), .Q(CNT_MUL[30]) );
  DFFR_X1 \CNT_MUL_reg[0]  ( .D(n437), .CK(CLK), .RN(n38), .Q(CNT_MUL[0]) );
  DFFR_X1 \CNT_MUL_reg[1]  ( .D(n436), .CK(CLK), .RN(n38), .Q(CNT_MUL[1]), 
        .QN(n451) );
  DFFR_X1 \CNT_MUL_reg[2]  ( .D(n435), .CK(CLK), .RN(n38), .Q(CNT_MUL[2]) );
  DFFR_X1 \CNT_MUL_reg[3]  ( .D(n434), .CK(CLK), .RN(n38), .Q(CNT_MUL[3]) );
  DFFR_X1 \CNT_MUL_reg[4]  ( .D(n433), .CK(CLK), .RN(n38), .Q(CNT_MUL[4]) );
  DFFR_X1 \CNT_MUL_reg[5]  ( .D(n432), .CK(CLK), .RN(n38), .Q(CNT_MUL[5]) );
  DFFR_X1 \CNT_MUL_reg[6]  ( .D(n431), .CK(CLK), .RN(n38), .Q(CNT_MUL[6]) );
  DFFR_X1 \CNT_MUL_reg[7]  ( .D(n430), .CK(CLK), .RN(n39), .Q(CNT_MUL[7]) );
  DFFR_X1 \CNT_MUL_reg[8]  ( .D(n429), .CK(CLK), .RN(n39), .Q(CNT_MUL[8]) );
  DFFR_X1 \CNT_MUL_reg[9]  ( .D(n428), .CK(CLK), .RN(n39), .Q(CNT_MUL[9]) );
  DFFR_X1 \CNT_MUL_reg[10]  ( .D(n427), .CK(CLK), .RN(n39), .Q(CNT_MUL[10]) );
  DFFR_X1 \CNT_MUL_reg[11]  ( .D(n426), .CK(CLK), .RN(n39), .Q(CNT_MUL[11]) );
  DFFR_X1 \CNT_MUL_reg[12]  ( .D(n425), .CK(CLK), .RN(n39), .Q(CNT_MUL[12]) );
  DFFR_X1 \CNT_MUL_reg[13]  ( .D(n424), .CK(CLK), .RN(n39), .Q(CNT_MUL[13]) );
  DFFR_X1 \CNT_MUL_reg[14]  ( .D(n423), .CK(CLK), .RN(n39), .Q(CNT_MUL[14]) );
  DFFR_X1 \CNT_MUL_reg[15]  ( .D(n422), .CK(CLK), .RN(n39), .Q(CNT_MUL[15]) );
  DFFR_X1 \CNT_MUL_reg[16]  ( .D(n421), .CK(CLK), .RN(n39), .Q(CNT_MUL[16]) );
  DFFR_X1 \CNT_MUL_reg[17]  ( .D(n420), .CK(CLK), .RN(n39), .Q(CNT_MUL[17]) );
  DFFR_X1 \CNT_MUL_reg[18]  ( .D(n419), .CK(CLK), .RN(n39), .Q(CNT_MUL[18]) );
  DFFR_X1 \CNT_MUL_reg[19]  ( .D(n418), .CK(CLK), .RN(n39), .Q(CNT_MUL[19]) );
  DFFR_X1 \CNT_MUL_reg[20]  ( .D(n417), .CK(CLK), .RN(n40), .Q(CNT_MUL[20]) );
  DFFR_X1 \CNT_MUL_reg[21]  ( .D(n416), .CK(CLK), .RN(n40), .Q(CNT_MUL[21]) );
  DFFR_X1 \CNT_MUL_reg[22]  ( .D(n415), .CK(CLK), .RN(n40), .Q(CNT_MUL[22]) );
  DFFR_X1 \CNT_MUL_reg[23]  ( .D(n414), .CK(CLK), .RN(n40), .Q(CNT_MUL[23]) );
  DFFR_X1 \CNT_MUL_reg[24]  ( .D(n413), .CK(CLK), .RN(n40), .Q(CNT_MUL[24]) );
  DFFR_X1 \CNT_MUL_reg[25]  ( .D(n412), .CK(CLK), .RN(n40), .Q(CNT_MUL[25]) );
  DFFR_X1 \CNT_MUL_reg[26]  ( .D(n411), .CK(CLK), .RN(n40), .Q(CNT_MUL[26]) );
  DFFR_X1 \CNT_MUL_reg[27]  ( .D(n410), .CK(CLK), .RN(n40), .Q(CNT_MUL[27]) );
  DFFR_X1 \CNT_MUL_reg[28]  ( .D(n409), .CK(CLK), .RN(n40), .Q(CNT_MUL[28]) );
  DFFR_X1 \CNT_MUL_reg[29]  ( .D(n408), .CK(CLK), .RN(n40), .Q(CNT_MUL[29]) );
  DFFR_X1 \CNT_MUL_reg[31]  ( .D(n407), .CK(CLK), .RN(n40), .Q(CNT_MUL[31]) );
  DFFS_X1 RST_DIV_reg ( .D(n406), .CK(CLK), .SN(n43), .Q(RST_DIV), .QN(n341)
         );
  DFFR_X1 \CNT_DIV_reg[29]  ( .D(n405), .CK(CLK), .RN(n40), .Q(CNT_DIV[29]), 
        .QN(n459) );
  DFFR_X1 \CNT_DIV_reg[27]  ( .D(n404), .CK(CLK), .RN(n41), .Q(CNT_DIV[27]), 
        .QN(n457) );
  DFFR_X1 \CNT_DIV_reg[25]  ( .D(n403), .CK(CLK), .RN(n41), .Q(CNT_DIV[25]), 
        .QN(n455) );
  DFFR_X1 \CNT_DIV_reg[23]  ( .D(n402), .CK(CLK), .RN(n41), .Q(CNT_DIV[23]), 
        .QN(n453) );
  DFFR_X1 \CNT_DIV_reg[21]  ( .D(n401), .CK(CLK), .RN(n41), .Q(CNT_DIV[21]), 
        .QN(n8) );
  DFFR_X1 \CNT_DIV_reg[19]  ( .D(n400), .CK(CLK), .RN(n41), .Q(CNT_DIV[19]), 
        .QN(n11) );
  DFFR_X1 \CNT_DIV_reg[17]  ( .D(n399), .CK(CLK), .RN(n41), .Q(CNT_DIV[17]), 
        .QN(n10) );
  DFFR_X1 \CNT_DIV_reg[15]  ( .D(n398), .CK(CLK), .RN(n41), .Q(CNT_DIV[15]), 
        .QN(n9) );
  DFFR_X1 \CNT_DIV_reg[13]  ( .D(n397), .CK(CLK), .RN(n41), .Q(CNT_DIV[13]), 
        .QN(n18) );
  DFFR_X1 \CNT_DIV_reg[11]  ( .D(n396), .CK(CLK), .RN(n41), .Q(CNT_DIV[11]), 
        .QN(n12) );
  DFFR_X1 \CNT_DIV_reg[9]  ( .D(n395), .CK(CLK), .RN(n41), .Q(CNT_DIV[9]), 
        .QN(n467) );
  DFFR_X1 \CNT_DIV_reg[7]  ( .D(n394), .CK(CLK), .RN(n41), .Q(CNT_DIV[7]), 
        .QN(n465) );
  DFFR_X1 \CNT_DIV_reg[5]  ( .D(n393), .CK(CLK), .RN(n41), .Q(CNT_DIV[5]), 
        .QN(n463) );
  DFFR_X1 \CNT_DIV_reg[3]  ( .D(n392), .CK(CLK), .RN(n41), .Q(CNT_DIV[3]), 
        .QN(n462) );
  DFFR_X1 \CNT_DIV_reg[1]  ( .D(n391), .CK(CLK), .RN(n42), .Q(CNT_DIV[1]), 
        .QN(n5) );
  DFFR_X1 \CNT_DIV_reg[2]  ( .D(n390), .CK(CLK), .RN(n42), .Q(CNT_DIV[2]), 
        .QN(n6) );
  DFFR_X1 \CNT_DIV_reg[4]  ( .D(n389), .CK(CLK), .RN(n42), .Q(CNT_DIV[4]), 
        .QN(n19) );
  DFFR_X1 \CNT_DIV_reg[6]  ( .D(n388), .CK(CLK), .RN(n42), .Q(CNT_DIV[6]), 
        .QN(n464) );
  DFFR_X1 \CNT_DIV_reg[8]  ( .D(n387), .CK(CLK), .RN(n42), .Q(CNT_DIV[8]), 
        .QN(n466) );
  DFFR_X1 \CNT_DIV_reg[12]  ( .D(n386), .CK(CLK), .RN(n42), .Q(CNT_DIV[12]), 
        .QN(n17) );
  DFFR_X1 \CNT_DIV_reg[14]  ( .D(n385), .CK(CLK), .RN(n42), .Q(CNT_DIV[14]), 
        .QN(n16) );
  DFFR_X1 \CNT_DIV_reg[16]  ( .D(n384), .CK(CLK), .RN(n42), .Q(CNT_DIV[16]), 
        .QN(n15) );
  DFFR_X1 \CNT_DIV_reg[18]  ( .D(n383), .CK(CLK), .RN(n42), .Q(CNT_DIV[18]), 
        .QN(n14) );
  DFFR_X1 \CNT_DIV_reg[20]  ( .D(n382), .CK(CLK), .RN(n42), .Q(CNT_DIV[20]), 
        .QN(n13) );
  DFFR_X1 \CNT_DIV_reg[22]  ( .D(n381), .CK(CLK), .RN(n42), .Q(CNT_DIV[22]), 
        .QN(n452) );
  DFFR_X1 \CNT_DIV_reg[24]  ( .D(n380), .CK(CLK), .RN(n42), .Q(CNT_DIV[24]), 
        .QN(n454) );
  DFFR_X1 \CNT_DIV_reg[26]  ( .D(n379), .CK(CLK), .RN(n42), .Q(CNT_DIV[26]), 
        .QN(n456) );
  DFFR_X1 \CNT_DIV_reg[28]  ( .D(n378), .CK(CLK), .RN(n43), .Q(CNT_DIV[28]), 
        .QN(n458) );
  DFFR_X1 \CNT_DIV_reg[30]  ( .D(n377), .CK(CLK), .RN(n43), .Q(CNT_DIV[30]), 
        .QN(n460) );
  DFFR_X1 STALL_INSTR_reg ( .D(n376), .CK(CLK), .RN(n43), .QN(n445) );
  DFFR_X1 \CURRENT_STATE_B_reg[2]  ( .D(N440), .CK(CLK), .RN(n43), .Q(n22), 
        .QN(n449) );
  DFFR_X1 \CURRENT_STATE_A_reg[2]  ( .D(N382), .CK(CLK), .RN(n43), .Q(n1), 
        .QN(n450) );
  DFFR_X1 \CURRENT_STATE_B_reg[0]  ( .D(N438), .CK(CLK), .RN(n43), .Q(n21), 
        .QN(n50) );
  DFFR_X1 \CURRENT_STATE_B_reg[1]  ( .D(N439), .CK(CLK), .RN(n43), .Q(n23), 
        .QN(n51) );
  DFFR_X1 \CURRENT_STATE_A_reg[0]  ( .D(N380), .CK(CLK), .RN(n43), .Q(n7), 
        .QN(n52) );
  DFFR_X1 \CURRENT_STATE_A_reg[1]  ( .D(N381), .CK(CLK), .RN(n43), .QN(n53) );
  DFFR_X1 \CURRENT_STATE_D_reg[2]  ( .D(n375), .CK(CLK), .RN(n43), .Q(n3), 
        .QN(n446) );
  DFFR_X1 \CURRENT_STATE_D_reg[0]  ( .D(n374), .CK(CLK), .RN(n43), .QN(n447)
         );
  DFFR_X1 \CURRENT_STATE_D_reg[1]  ( .D(n373), .CK(CLK), .RN(n38), .Q(
        \CURRENT_STATE_D[1] ), .QN(n4) );
  OAI33_X1 U5 ( .A1(n59), .A2(n447), .A3(n60), .B1(n61), .B2(n62), .B3(n63), 
        .ZN(n58) );
  NAND3_X1 U14 ( .A1(n73), .A2(n446), .A3(n74), .ZN(n72) );
  NAND3_X1 U28 ( .A1(OPCODE_IF[2]), .A2(n84), .A3(n85), .ZN(n62) );
  NAND3_X1 U32 ( .A1(n86), .A2(n88), .A3(n89), .ZN(n87) );
  NAND2_X1 U38 ( .A1(N608), .A2(n32), .ZN(n99) );
  NAND2_X1 U40 ( .A1(N606), .A2(n32), .ZN(n101) );
  NAND2_X1 U42 ( .A1(N604), .A2(n32), .ZN(n102) );
  NAND2_X1 U44 ( .A1(N602), .A2(n32), .ZN(n103) );
  NAND2_X1 U46 ( .A1(N600), .A2(n32), .ZN(n104) );
  NAND2_X1 U48 ( .A1(N598), .A2(n32), .ZN(n106) );
  NAND2_X1 U51 ( .A1(N596), .A2(n32), .ZN(n108) );
  NAND2_X1 U54 ( .A1(N594), .A2(n32), .ZN(n110) );
  NAND2_X1 U57 ( .A1(N592), .A2(n32), .ZN(n112) );
  NAND2_X1 U60 ( .A1(N590), .A2(n32), .ZN(n114) );
  NAND2_X1 U63 ( .A1(N586), .A2(n32), .ZN(n115) );
  NAND2_X1 U65 ( .A1(N584), .A2(n32), .ZN(n116) );
  NAND2_X1 U67 ( .A1(N582), .A2(n32), .ZN(n118) );
  NAND2_X1 U70 ( .A1(N580), .A2(n33), .ZN(n120) );
  NAND2_X1 U72 ( .A1(N579), .A2(n33), .ZN(n121) );
  NAND2_X1 U74 ( .A1(N581), .A2(n33), .ZN(n122) );
  NAND2_X1 U76 ( .A1(N583), .A2(n33), .ZN(n123) );
  NAND2_X1 U78 ( .A1(N585), .A2(n33), .ZN(n124) );
  NAND2_X1 U80 ( .A1(N587), .A2(n33), .ZN(n125) );
  NAND2_X1 U82 ( .A1(N589), .A2(n33), .ZN(n127) );
  NAND2_X1 U85 ( .A1(N591), .A2(n33), .ZN(n129) );
  NAND2_X1 U88 ( .A1(N593), .A2(n33), .ZN(n131) );
  NAND2_X1 U91 ( .A1(N595), .A2(n33), .ZN(n133) );
  NAND2_X1 U94 ( .A1(N597), .A2(n33), .ZN(n135) );
  NAND2_X1 U97 ( .A1(N599), .A2(n33), .ZN(n137) );
  NAND2_X1 U100 ( .A1(N601), .A2(n33), .ZN(n138) );
  NAND2_X1 U102 ( .A1(N603), .A2(n34), .ZN(n139) );
  NAND2_X1 U104 ( .A1(N605), .A2(n34), .ZN(n140) );
  NAND2_X1 U106 ( .A1(N607), .A2(n34), .ZN(n141) );
  NAND2_X1 U173 ( .A1(n179), .A2(n144), .ZN(n175) );
  NAND2_X1 U177 ( .A1(n183), .A2(n184), .ZN(n92) );
  NAND2_X1 U191 ( .A1(N609), .A2(n34), .ZN(n194) );
  NAND2_X1 U193 ( .A1(N588), .A2(n34), .ZN(n195) );
  NAND2_X1 U195 ( .A1(N578), .A2(n34), .ZN(n196) );
  OAI33_X1 U199 ( .A1(n181), .A2(N342), .A3(n180), .B1(n199), .B2(n82), .B3(n5), .ZN(n198) );
  NAND3_X1 U203 ( .A1(n466), .A2(n465), .A3(n467), .ZN(n207) );
  NAND2_X1 U212 ( .A1(N342), .A2(n468), .ZN(n199) );
  NAND2_X1 U215 ( .A1(n88), .A2(n209), .ZN(n197) );
  NAND3_X1 U216 ( .A1(OPCODE_ID[0]), .A2(n95), .A3(n182), .ZN(n209) );
  NAND3_X1 U223 ( .A1(CMP_C_EXE), .A2(n218), .A3(n219), .ZN(n217) );
  NAND2_X1 U265 ( .A1(n263), .A2(n264), .ZN(n244) );
  NAND3_X1 U266 ( .A1(n265), .A2(n266), .A3(n267), .ZN(n264) );
  OAI33_X1 U272 ( .A1(n279), .A2(OPCODE_ID[5]), .A3(OPCODE_ID[0]), .B1(n280), 
        .B2(n266), .B3(n269), .ZN(n274) );
  NAND2_X1 U274 ( .A1(OPCODE_ID[1]), .A2(n265), .ZN(n280) );
  NAND2_X1 U277 ( .A1(OPCODE_ID[0]), .A2(OPCODE_ID[5]), .ZN(n283) );
  NAND3_X1 U282 ( .A1(n285), .A2(n278), .A3(n286), .ZN(n270) );
  NAND2_X1 U291 ( .A1(OPCODE_ID[3]), .A2(n278), .ZN(n277) );
  NAND3_X1 U298 ( .A1(n88), .A2(n95), .A3(n60), .ZN(n249) );
  NAND2_X1 U311 ( .A1(n298), .A2(n299), .ZN(n293) );
  NAND2_X1 U312 ( .A1(OPCODE_MEM[0]), .A2(n298), .ZN(n294) );
  NAND3_X1 U318 ( .A1(n299), .A2(n297), .A3(OPCODE_MEM[2]), .ZN(n292) );
  NAND2_X1 U324 ( .A1(n305), .A2(n231), .ZN(n79) );
  NAND3_X1 U330 ( .A1(OPCODE_EXE[0]), .A2(n313), .A3(n312), .ZN(n307) );
  NAND3_X1 U335 ( .A1(OPCODE_EXE[1]), .A2(n316), .A3(n320), .ZN(n181) );
  NAND2_X1 U343 ( .A1(n320), .A2(OPCODE_EXE[3]), .ZN(n212) );
  FORW_FSM_OPCODE_SIZE6_N_ADDR5_DW01_inc_0 r233 ( .A(CNT_DIV), .SUM({N609, 
        N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, 
        N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, 
        N584, N583, N582, N581, N580, N579, N578}) );
  FORW_FSM_OPCODE_SIZE6_N_ADDR5_DW01_inc_1 r232 ( .A(CNT_MUL), .SUM({N539, 
        N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, 
        N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, 
        N514, N513, N512, N511, N510, N509, N508}) );
  INV_X1 U3 ( .A(n1), .ZN(n2) );
  NAND2_X1 U4 ( .A1(n52), .A2(n53), .ZN(n49) );
  AOI21_X2 U6 ( .B1(n21), .B2(n22), .A(n23), .ZN(MUX_B[1]) );
  BUF_X1 U7 ( .A(n142), .Z(n31) );
  BUF_X1 U8 ( .A(n146), .Z(n28) );
  BUF_X1 U9 ( .A(n142), .Z(n30) );
  BUF_X1 U10 ( .A(n142), .Z(n29) );
  BUF_X1 U11 ( .A(n146), .Z(n27) );
  BUF_X1 U12 ( .A(n146), .Z(n26) );
  NOR2_X1 U13 ( .A1(n77), .A2(n230), .ZN(n67) );
  INV_X1 U15 ( .A(n144), .ZN(n142) );
  AOI21_X1 U16 ( .B1(n248), .B2(n249), .A(n233), .ZN(n247) );
  INV_X1 U17 ( .A(n175), .ZN(n146) );
  BUF_X1 U18 ( .A(n98), .Z(n37) );
  BUF_X1 U19 ( .A(n98), .Z(n35) );
  BUF_X1 U20 ( .A(n100), .Z(n32) );
  BUF_X1 U21 ( .A(n100), .Z(n33) );
  BUF_X1 U22 ( .A(n98), .Z(n36) );
  INV_X1 U23 ( .A(n245), .ZN(n75) );
  BUF_X1 U24 ( .A(n100), .Z(n34) );
  INV_X1 U25 ( .A(n230), .ZN(n248) );
  INV_X1 U26 ( .A(n69), .ZN(n250) );
  INV_X1 U27 ( .A(n218), .ZN(n61) );
  INV_X1 U29 ( .A(n79), .ZN(n60) );
  INV_X1 U30 ( .A(n281), .ZN(n269) );
  NOR2_X1 U31 ( .A1(n3), .A2(n4), .ZN(MUX_D[1]) );
  INV_X1 U33 ( .A(n62), .ZN(n70) );
  INV_X1 U34 ( .A(n54), .ZN(n57) );
  OR3_X1 U35 ( .A1(CMP_BRANCH_EXE), .A2(CMP_BRANCH_ID), .A3(n3), .ZN(n63) );
  INV_X1 U36 ( .A(n76), .ZN(n73) );
  AOI21_X1 U37 ( .B1(n77), .B2(CMP_BRANCH_EXE), .A(CMP_BRANCH_ID), .ZN(n76) );
  OAI21_X1 U39 ( .B1(n305), .B2(n231), .A(n79), .ZN(n77) );
  NOR2_X1 U41 ( .A1(n231), .A2(n290), .ZN(n230) );
  OAI21_X1 U43 ( .B1(n193), .B2(N342), .A(n88), .ZN(n144) );
  NOR2_X1 U45 ( .A1(n295), .A2(n296), .ZN(n218) );
  AOI21_X1 U47 ( .B1(n294), .B2(n293), .A(n297), .ZN(n296) );
  INV_X1 U49 ( .A(n301), .ZN(n295) );
  OAI21_X1 U50 ( .B1(n302), .B2(n303), .A(n300), .ZN(n301) );
  NOR4_X1 U52 ( .A1(n230), .A2(n231), .A3(n251), .A4(n252), .ZN(N382) );
  NOR4_X1 U53 ( .A1(n230), .A2(n231), .A3(n232), .A4(n233), .ZN(N440) );
  NOR2_X1 U55 ( .A1(n61), .A2(n219), .ZN(n69) );
  NAND4_X1 U56 ( .A1(n263), .A2(n270), .A3(n271), .A4(n272), .ZN(n245) );
  AOI21_X1 U58 ( .B1(n282), .B2(n281), .A(n284), .ZN(n271) );
  NOR4_X1 U59 ( .A1(n273), .A2(n274), .A3(n275), .A4(n276), .ZN(n272) );
  NOR2_X1 U61 ( .A1(n91), .A2(n197), .ZN(n100) );
  OAI21_X1 U62 ( .B1(N342), .B2(n193), .A(n143), .ZN(n91) );
  NOR2_X1 U64 ( .A1(n285), .A2(n278), .ZN(n281) );
  OAI22_X1 U66 ( .A1(n80), .A2(n88), .B1(N341), .B2(n90), .ZN(n179) );
  AOI21_X1 U68 ( .B1(CMP_B_EXE), .B2(n77), .A(n250), .ZN(n246) );
  INV_X1 U69 ( .A(N341), .ZN(n88) );
  INV_X1 U71 ( .A(N342), .ZN(n95) );
  INV_X1 U73 ( .A(n197), .ZN(n98) );
  NOR2_X1 U75 ( .A1(n268), .A2(n277), .ZN(n284) );
  NOR2_X1 U77 ( .A1(CMP_B_EXE), .A2(CMP_A_EXE), .ZN(n180) );
  AOI21_X1 U79 ( .B1(CMP_A_EXE), .B2(n77), .A(n250), .ZN(n288) );
  NOR2_X1 U81 ( .A1(n193), .A2(n182), .ZN(n263) );
  NOR2_X1 U83 ( .A1(n232), .A2(n239), .ZN(n238) );
  INV_X1 U84 ( .A(CMP_B_MEM), .ZN(n239) );
  AND2_X1 U86 ( .A1(n284), .A2(n286), .ZN(n193) );
  INV_X1 U87 ( .A(CMP_B_EXE), .ZN(n233) );
  OAI21_X1 U89 ( .B1(n36), .B2(n6), .A(n120), .ZN(n390) );
  OAI21_X1 U90 ( .B1(n36), .B2(n5), .A(n121), .ZN(n391) );
  INV_X1 U92 ( .A(n92), .ZN(n80) );
  INV_X1 U93 ( .A(n290), .ZN(n305) );
  INV_X1 U95 ( .A(CMP_A_EXE), .ZN(n252) );
  NOR2_X1 U96 ( .A1(\CURRENT_STATE_D[1] ), .A2(n446), .ZN(STALL_BRANCH) );
  OAI21_X1 U98 ( .B1(n446), .B2(n4), .A(n83), .ZN(n54) );
  OR3_X1 U99 ( .A1(CMP_BRANCH_MEM), .A2(n62), .A3(n63), .ZN(n83) );
  INV_X1 U101 ( .A(OPCODE_IF[1]), .ZN(n84) );
  NOR3_X1 U103 ( .A1(OPCODE_IF[3]), .A2(OPCODE_IF[5]), .A3(OPCODE_IF[4]), .ZN(
        n85) );
  INV_X1 U105 ( .A(n145), .ZN(n407) );
  AOI22_X1 U107 ( .A1(n31), .A2(CNT_MUL[31]), .B1(n28), .B2(N539), .ZN(n145)
         );
  OAI22_X1 U108 ( .A1(n447), .A2(n57), .B1(n64), .B2(n54), .ZN(n374) );
  NOR2_X1 U109 ( .A1(n65), .A2(n3), .ZN(n64) );
  AOI211_X1 U110 ( .C1(CMP_BRANCH_EXE), .C2(n67), .A(n68), .B(CMP_BRANCH_ID), 
        .ZN(n65) );
  OAI21_X1 U111 ( .B1(CMP_BRANCH_EXE), .B2(n69), .A(n70), .ZN(n68) );
  OAI22_X1 U112 ( .A1(n54), .A2(n55), .B1(n4), .B2(n57), .ZN(n373) );
  INV_X1 U113 ( .A(n58), .ZN(n55) );
  INV_X1 U114 ( .A(STALL_BRANCH), .ZN(n59) );
  NOR2_X1 U115 ( .A1(n447), .A2(n3), .ZN(MUX_D[0]) );
  OAI21_X1 U116 ( .B1(n446), .B2(n71), .A(n72), .ZN(n375) );
  AOI211_X1 U117 ( .C1(n447), .C2(n77), .A(n54), .B(n78), .ZN(n71) );
  AOI21_X1 U118 ( .B1(CMP_BRANCH_ID), .B2(n75), .A(n62), .ZN(n74) );
  OAI21_X1 U119 ( .B1(n453), .B2(n36), .A(n138), .ZN(n402) );
  OAI21_X1 U120 ( .B1(n457), .B2(n36), .A(n140), .ZN(n404) );
  OAI21_X1 U121 ( .B1(n461), .B2(n36), .A(n194), .ZN(n439) );
  OAI21_X1 U122 ( .B1(n458), .B2(n35), .A(n101), .ZN(n378) );
  OAI21_X1 U123 ( .B1(n454), .B2(n35), .A(n103), .ZN(n380) );
  OAI21_X1 U124 ( .B1(n455), .B2(n36), .A(n139), .ZN(n403) );
  OAI21_X1 U125 ( .B1(n459), .B2(n36), .A(n141), .ZN(n405) );
  OAI21_X1 U126 ( .B1(n460), .B2(n35), .A(n99), .ZN(n377) );
  OAI21_X1 U127 ( .B1(n456), .B2(n35), .A(n102), .ZN(n379) );
  OAI21_X1 U128 ( .B1(n452), .B2(n35), .A(n104), .ZN(n381) );
  OR2_X1 U129 ( .A1(n49), .A2(n450), .ZN(n24) );
  INV_X1 U130 ( .A(n147), .ZN(n408) );
  AOI22_X1 U131 ( .A1(n31), .A2(CNT_MUL[29]), .B1(n28), .B2(N537), .ZN(n147)
         );
  INV_X1 U132 ( .A(n148), .ZN(n409) );
  AOI22_X1 U133 ( .A1(n31), .A2(CNT_MUL[28]), .B1(n28), .B2(N536), .ZN(n148)
         );
  INV_X1 U134 ( .A(n149), .ZN(n410) );
  AOI22_X1 U135 ( .A1(n31), .A2(CNT_MUL[27]), .B1(n28), .B2(N535), .ZN(n149)
         );
  INV_X1 U136 ( .A(n150), .ZN(n411) );
  AOI22_X1 U137 ( .A1(n31), .A2(CNT_MUL[26]), .B1(n28), .B2(N534), .ZN(n150)
         );
  INV_X1 U138 ( .A(n151), .ZN(n412) );
  AOI22_X1 U139 ( .A1(n30), .A2(CNT_MUL[25]), .B1(n27), .B2(N533), .ZN(n151)
         );
  INV_X1 U140 ( .A(n152), .ZN(n413) );
  AOI22_X1 U141 ( .A1(n30), .A2(CNT_MUL[24]), .B1(n27), .B2(N532), .ZN(n152)
         );
  INV_X1 U142 ( .A(n153), .ZN(n414) );
  AOI22_X1 U143 ( .A1(n30), .A2(CNT_MUL[23]), .B1(n27), .B2(N531), .ZN(n153)
         );
  INV_X1 U144 ( .A(n154), .ZN(n415) );
  AOI22_X1 U145 ( .A1(n30), .A2(CNT_MUL[22]), .B1(n27), .B2(N530), .ZN(n154)
         );
  INV_X1 U146 ( .A(n178), .ZN(n438) );
  AOI22_X1 U147 ( .A1(n29), .A2(CNT_MUL[30]), .B1(n26), .B2(N538), .ZN(n178)
         );
  INV_X1 U148 ( .A(n282), .ZN(n279) );
  NOR4_X1 U149 ( .A1(CMP_C_EXE), .A2(n220), .A3(n221), .A4(n222), .ZN(n215) );
  NOR3_X1 U150 ( .A1(n229), .A2(OPCODE_WB[0]), .A3(n228), .ZN(n220) );
  AOI21_X1 U151 ( .B1(n223), .B2(n224), .A(n225), .ZN(n221) );
  OAI221_X1 U152 ( .B1(OPCODE_WB[4]), .B2(n223), .C1(OPCODE_WB[1]), .C2(n224), 
        .A(CMP_C_MEM), .ZN(n222) );
  NOR4_X1 U153 ( .A1(OPCODE_ID[4]), .A2(OPCODE_ID[3]), .A3(OPCODE_ID[1]), .A4(
        n278), .ZN(n275) );
  NOR4_X1 U154 ( .A1(n283), .A2(OPCODE_ID[2]), .A3(OPCODE_ID[4]), .A4(
        OPCODE_ID[3]), .ZN(n273) );
  NOR4_X1 U155 ( .A1(n315), .A2(n313), .A3(OPCODE_EXE[2]), .A4(OPCODE_EXE[4]), 
        .ZN(n320) );
  NOR4_X1 U156 ( .A1(OPCODE_MEM[3]), .A2(OPCODE_MEM[2]), .A3(OPCODE_MEM[0]), 
        .A4(n299), .ZN(n302) );
  NOR3_X1 U157 ( .A1(OPCODE_EXE[3]), .A2(OPCODE_EXE[4]), .A3(OPCODE_EXE[1]), 
        .ZN(n312) );
  NOR3_X1 U158 ( .A1(n265), .A2(OPCODE_ID[1]), .A3(n266), .ZN(n282) );
  AOI211_X1 U159 ( .C1(n94), .C2(n468), .A(n95), .B(n96), .ZN(n93) );
  NOR2_X1 U160 ( .A1(n82), .A2(n5), .ZN(n94) );
  NAND4_X1 U161 ( .A1(n306), .A2(n212), .A3(n307), .A4(n308), .ZN(n231) );
  NOR4_X1 U162 ( .A1(n309), .A2(n96), .A3(n310), .A4(n311), .ZN(n308) );
  AND3_X1 U163 ( .A1(n312), .A2(n313), .A3(OPCODE_EXE[2]), .ZN(n310) );
  OAI211_X1 U164 ( .C1(n245), .C2(n244), .A(n445), .B(n2), .ZN(n251) );
  OAI211_X1 U165 ( .C1(n180), .C2(n181), .A(OPCODE_ID[0]), .B(n182), .ZN(n90)
         );
  AOI211_X1 U166 ( .C1(n216), .C2(n217), .A(n212), .B(n214), .ZN(N458) );
  INV_X1 U167 ( .A(n215), .ZN(n216) );
  AOI21_X1 U168 ( .B1(OPCODE_ID[1]), .B2(n268), .A(n269), .ZN(n267) );
  NOR3_X1 U169 ( .A1(n79), .A2(n80), .A3(n81), .ZN(n78) );
  NOR3_X1 U170 ( .A1(n82), .A2(n468), .A3(CNT_DIV[1]), .ZN(n81) );
  NOR3_X1 U171 ( .A1(OPCODE_MEM[2]), .A2(OPCODE_MEM[4]), .A3(n300), .ZN(n298)
         );
  NAND4_X1 U172 ( .A1(n200), .A2(n201), .A3(n202), .A4(n203), .ZN(n82) );
  NOR4_X1 U174 ( .A1(CNT_DIV[17]), .A2(CNT_DIV[16]), .A3(CNT_DIV[15]), .A4(
        CNT_DIV[14]), .ZN(n200) );
  NOR4_X1 U175 ( .A1(CNT_DIV[21]), .A2(CNT_DIV[20]), .A3(CNT_DIV[19]), .A4(
        CNT_DIV[18]), .ZN(n201) );
  NOR4_X1 U176 ( .A1(n204), .A2(n205), .A3(n206), .A4(n207), .ZN(n203) );
  NAND4_X1 U178 ( .A1(n449), .A2(n445), .A3(n244), .A4(n245), .ZN(n232) );
  NAND4_X1 U179 ( .A1(OPCODE_EXE[1]), .A2(n315), .A3(n322), .A4(n323), .ZN(
        n306) );
  INV_X1 U180 ( .A(OPCODE_EXE[2]), .ZN(n323) );
  OAI22_X1 U181 ( .A1(n31), .A2(n341), .B1(n143), .B2(n144), .ZN(n406) );
  OAI22_X1 U182 ( .A1(n451), .A2(n144), .B1(n175), .B2(n176), .ZN(n436) );
  INV_X1 U183 ( .A(N509), .ZN(n176) );
  NAND4_X1 U184 ( .A1(n306), .A2(n212), .A3(n317), .A4(n318), .ZN(n290) );
  OAI21_X1 U185 ( .B1(OPCODE_EXE[2]), .B2(OPCODE_EXE[5]), .A(n312), .ZN(n317)
         );
  NOR3_X1 U186 ( .A1(n311), .A2(n309), .A3(n319), .ZN(n318) );
  INV_X1 U187 ( .A(n181), .ZN(n319) );
  AOI21_X1 U188 ( .B1(OPCODE_ID[4]), .B2(OPCODE_ID[2]), .A(n277), .ZN(n276) );
  NAND4_X1 U189 ( .A1(OPCODE_WB[2]), .A2(n228), .A3(n227), .A4(n226), .ZN(n223) );
  AOI21_X1 U190 ( .B1(OPCODE_MEM[4]), .B2(n304), .A(n292), .ZN(n303) );
  INV_X1 U192 ( .A(OPCODE_MEM[0]), .ZN(n304) );
  AOI21_X1 U194 ( .B1(n75), .B2(n262), .A(n445), .ZN(n237) );
  INV_X1 U196 ( .A(n244), .ZN(n262) );
  NOR3_X1 U197 ( .A1(n212), .A2(n213), .A3(n214), .ZN(N459) );
  AOI21_X1 U198 ( .B1(CMP_C_EXE), .B2(n69), .A(n215), .ZN(n213) );
  NOR2_X1 U200 ( .A1(OPCODE_EXE[5]), .A2(OPCODE_EXE[3]), .ZN(n322) );
  NOR4_X1 U201 ( .A1(n185), .A2(n186), .A3(n187), .A4(n188), .ZN(n184) );
  NOR4_X1 U202 ( .A1(n189), .A2(n190), .A3(n191), .A4(n192), .ZN(n183) );
  OR4_X1 U204 ( .A1(CNT_MUL[7]), .A2(CNT_MUL[8]), .A3(CNT_MUL[9]), .A4(n451), 
        .ZN(n185) );
  AOI21_X1 U205 ( .B1(n246), .B2(CMP_B_MEM), .A(n247), .ZN(n240) );
  OR4_X1 U206 ( .A1(n226), .A2(n227), .A3(OPCODE_WB[2]), .A4(OPCODE_WB[4]), 
        .ZN(n224) );
  OAI21_X1 U207 ( .B1(n445), .B2(n86), .A(n87), .ZN(n376) );
  OAI22_X1 U208 ( .A1(n92), .A2(n88), .B1(N341), .B2(n93), .ZN(n86) );
  OAI21_X1 U209 ( .B1(N342), .B2(n90), .A(n91), .ZN(n89) );
  AND4_X1 U210 ( .A1(n266), .A2(n278), .A3(n285), .A4(n287), .ZN(n182) );
  NOR2_X1 U211 ( .A1(OPCODE_ID[2]), .A2(OPCODE_ID[1]), .ZN(n287) );
  NAND4_X1 U213 ( .A1(n464), .A2(n463), .A3(n462), .A4(n461), .ZN(n206) );
  NAND4_X1 U214 ( .A1(n460), .A2(n459), .A3(n458), .A4(n457), .ZN(n205) );
  NAND4_X1 U217 ( .A1(n456), .A2(n455), .A3(n454), .A4(n453), .ZN(n204) );
  INV_X1 U218 ( .A(n198), .ZN(n143) );
  OR4_X1 U219 ( .A1(CNT_MUL[0]), .A2(CNT_MUL[10]), .A3(CNT_MUL[11]), .A4(
        CNT_MUL[12]), .ZN(n192) );
  OR4_X1 U220 ( .A1(CNT_MUL[25]), .A2(CNT_MUL[26]), .A3(CNT_MUL[27]), .A4(
        CNT_MUL[28]), .ZN(n188) );
  OR4_X1 U221 ( .A1(CNT_MUL[13]), .A2(CNT_MUL[14]), .A3(CNT_MUL[15]), .A4(
        CNT_MUL[16]), .ZN(n191) );
  OR4_X1 U222 ( .A1(CNT_MUL[29]), .A2(CNT_MUL[2]), .A3(CNT_MUL[30]), .A4(
        CNT_MUL[31]), .ZN(n187) );
  OR4_X1 U224 ( .A1(CNT_MUL[17]), .A2(CNT_MUL[18]), .A3(CNT_MUL[19]), .A4(
        CNT_MUL[20]), .ZN(n190) );
  OR4_X1 U225 ( .A1(CNT_MUL[3]), .A2(CNT_MUL[4]), .A3(CNT_MUL[5]), .A4(
        CNT_MUL[6]), .ZN(n186) );
  INV_X1 U226 ( .A(OPCODE_ID[5]), .ZN(n278) );
  OR4_X1 U227 ( .A1(CNT_MUL[21]), .A2(CNT_MUL[22]), .A3(CNT_MUL[23]), .A4(
        CNT_MUL[24]), .ZN(n189) );
  AND4_X1 U228 ( .A1(OPCODE_EXE[2]), .A2(OPCODE_EXE[0]), .A3(n322), .A4(n214), 
        .ZN(n311) );
  AND4_X1 U229 ( .A1(OPCODE_EXE[2]), .A2(OPCODE_EXE[1]), .A3(OPCODE_EXE[4]), 
        .A4(n314), .ZN(n96) );
  NOR3_X1 U230 ( .A1(n315), .A2(OPCODE_EXE[5]), .A3(n316), .ZN(n314) );
  INV_X1 U231 ( .A(OPCODE_EXE[1]), .ZN(n214) );
  AND4_X1 U232 ( .A1(OPCODE_EXE[5]), .A2(OPCODE_EXE[3]), .A3(n321), .A4(n214), 
        .ZN(n309) );
  NOR2_X1 U233 ( .A1(OPCODE_EXE[4]), .A2(OPCODE_EXE[2]), .ZN(n321) );
  OAI211_X1 U234 ( .C1(n97), .C2(n53), .A(n24), .B(n253), .ZN(N381) );
  OAI211_X1 U235 ( .C1(n67), .C2(n252), .A(n218), .B(n256), .ZN(n253) );
  NOR2_X1 U236 ( .A1(n251), .A2(n257), .ZN(n256) );
  INV_X1 U237 ( .A(CMP_A_MEM), .ZN(n257) );
  INV_X1 U238 ( .A(OPCODE_ID[4]), .ZN(n266) );
  OAI21_X1 U239 ( .B1(n468), .B2(n35), .A(n196), .ZN(n441) );
  INV_X1 U240 ( .A(OPCODE_EXE[0]), .ZN(n315) );
  INV_X1 U241 ( .A(OPCODE_ID[2]), .ZN(n265) );
  INV_X1 U242 ( .A(OPCODE_EXE[5]), .ZN(n313) );
  OAI21_X1 U243 ( .B1(n37), .B2(n13), .A(n106), .ZN(n382) );
  OAI21_X1 U244 ( .B1(n37), .B2(n14), .A(n108), .ZN(n383) );
  OAI21_X1 U245 ( .B1(n37), .B2(n15), .A(n110), .ZN(n384) );
  OAI21_X1 U246 ( .B1(n37), .B2(n16), .A(n112), .ZN(n385) );
  OAI21_X1 U247 ( .B1(n37), .B2(n17), .A(n114), .ZN(n386) );
  OAI21_X1 U248 ( .B1(n448), .B2(n35), .A(n195), .ZN(n440) );
  OAI21_X1 U249 ( .B1(n36), .B2(n12), .A(n127), .ZN(n396) );
  OAI21_X1 U250 ( .B1(n36), .B2(n18), .A(n129), .ZN(n397) );
  OAI21_X1 U251 ( .B1(n36), .B2(n9), .A(n131), .ZN(n398) );
  OAI21_X1 U252 ( .B1(n36), .B2(n10), .A(n133), .ZN(n399) );
  OAI21_X1 U253 ( .B1(n36), .B2(n11), .A(n135), .ZN(n400) );
  OAI21_X1 U254 ( .B1(n36), .B2(n8), .A(n137), .ZN(n401) );
  INV_X1 U255 ( .A(OPCODE_ID[3]), .ZN(n285) );
  INV_X1 U256 ( .A(OPCODE_ID[0]), .ZN(n268) );
  OAI21_X1 U257 ( .B1(n466), .B2(n35), .A(n115), .ZN(n387) );
  OAI21_X1 U258 ( .B1(n464), .B2(n35), .A(n116), .ZN(n388) );
  OAI21_X1 U259 ( .B1(n37), .B2(n19), .A(n118), .ZN(n389) );
  OAI21_X1 U260 ( .B1(n462), .B2(n35), .A(n122), .ZN(n392) );
  OAI21_X1 U261 ( .B1(n463), .B2(n35), .A(n123), .ZN(n393) );
  OAI21_X1 U262 ( .B1(n465), .B2(n35), .A(n124), .ZN(n394) );
  OAI21_X1 U263 ( .B1(n467), .B2(n35), .A(n125), .ZN(n395) );
  INV_X1 U264 ( .A(OPCODE_EXE[3]), .ZN(n316) );
  AND4_X1 U267 ( .A1(n208), .A2(n452), .A3(CNT_DIV[4]), .A4(n448), .ZN(n202)
         );
  NOR4_X1 U268 ( .A1(n6), .A2(CNT_DIV[11]), .A3(CNT_DIV[12]), .A4(CNT_DIV[13]), 
        .ZN(n208) );
  OAI211_X1 U269 ( .C1(n67), .C2(n233), .A(n218), .B(n238), .ZN(n234) );
  INV_X1 U270 ( .A(OPCODE_MEM[1]), .ZN(n299) );
  OR3_X1 U271 ( .A1(OPCODE_WB[3]), .A2(OPCODE_WB[5]), .A3(OPCODE_WB[2]), .ZN(
        n229) );
  INV_X1 U273 ( .A(OPCODE_WB[1]), .ZN(n228) );
  INV_X1 U275 ( .A(OPCODE_MEM[5]), .ZN(n300) );
  AND3_X1 U276 ( .A1(OPCODE_ID[2]), .A2(OPCODE_ID[1]), .A3(OPCODE_ID[4]), .ZN(
        n286) );
  AND2_X1 U278 ( .A1(n237), .A2(n449), .ZN(n25) );
  INV_X1 U279 ( .A(n291), .ZN(n219) );
  OAI211_X1 U280 ( .C1(OPCODE_MEM[4]), .C2(n292), .A(n293), .B(n294), .ZN(n291) );
  INV_X1 U281 ( .A(OPCODE_WB[5]), .ZN(n226) );
  INV_X1 U283 ( .A(OPCODE_MEM[3]), .ZN(n297) );
  INV_X1 U284 ( .A(OPCODE_WB[3]), .ZN(n227) );
  INV_X1 U285 ( .A(OPCODE_WB[0]), .ZN(n225) );
  INV_X1 U286 ( .A(n155), .ZN(n416) );
  AOI22_X1 U287 ( .A1(n30), .A2(CNT_MUL[21]), .B1(n27), .B2(N529), .ZN(n155)
         );
  INV_X1 U288 ( .A(n156), .ZN(n417) );
  AOI22_X1 U289 ( .A1(n30), .A2(CNT_MUL[20]), .B1(n27), .B2(N528), .ZN(n156)
         );
  INV_X1 U290 ( .A(n157), .ZN(n418) );
  AOI22_X1 U292 ( .A1(n30), .A2(CNT_MUL[19]), .B1(n27), .B2(N527), .ZN(n157)
         );
  INV_X1 U293 ( .A(n158), .ZN(n419) );
  AOI22_X1 U294 ( .A1(n30), .A2(CNT_MUL[18]), .B1(n27), .B2(N526), .ZN(n158)
         );
  INV_X1 U295 ( .A(n159), .ZN(n420) );
  AOI22_X1 U296 ( .A1(n30), .A2(CNT_MUL[17]), .B1(n27), .B2(N525), .ZN(n159)
         );
  INV_X1 U297 ( .A(n160), .ZN(n421) );
  AOI22_X1 U299 ( .A1(n30), .A2(CNT_MUL[16]), .B1(n27), .B2(N524), .ZN(n160)
         );
  INV_X1 U300 ( .A(n161), .ZN(n422) );
  AOI22_X1 U301 ( .A1(n30), .A2(CNT_MUL[15]), .B1(n27), .B2(N523), .ZN(n161)
         );
  INV_X1 U302 ( .A(n162), .ZN(n423) );
  AOI22_X1 U303 ( .A1(n30), .A2(CNT_MUL[14]), .B1(n27), .B2(N522), .ZN(n162)
         );
  INV_X1 U304 ( .A(n163), .ZN(n424) );
  AOI22_X1 U305 ( .A1(n30), .A2(CNT_MUL[13]), .B1(n27), .B2(N521), .ZN(n163)
         );
  INV_X1 U306 ( .A(n164), .ZN(n425) );
  AOI22_X1 U307 ( .A1(n29), .A2(CNT_MUL[12]), .B1(n26), .B2(N520), .ZN(n164)
         );
  INV_X1 U308 ( .A(n165), .ZN(n426) );
  AOI22_X1 U309 ( .A1(n29), .A2(CNT_MUL[11]), .B1(n26), .B2(N519), .ZN(n165)
         );
  INV_X1 U310 ( .A(n166), .ZN(n427) );
  AOI22_X1 U313 ( .A1(n29), .A2(CNT_MUL[10]), .B1(n26), .B2(N518), .ZN(n166)
         );
  INV_X1 U314 ( .A(n167), .ZN(n428) );
  AOI22_X1 U315 ( .A1(n29), .A2(CNT_MUL[9]), .B1(n26), .B2(N517), .ZN(n167) );
  INV_X1 U316 ( .A(n168), .ZN(n429) );
  AOI22_X1 U317 ( .A1(n29), .A2(CNT_MUL[8]), .B1(n26), .B2(N516), .ZN(n168) );
  INV_X1 U319 ( .A(n169), .ZN(n430) );
  AOI22_X1 U320 ( .A1(n29), .A2(CNT_MUL[7]), .B1(n26), .B2(N515), .ZN(n169) );
  INV_X1 U321 ( .A(n170), .ZN(n431) );
  AOI22_X1 U322 ( .A1(n29), .A2(CNT_MUL[6]), .B1(n26), .B2(N514), .ZN(n170) );
  INV_X1 U323 ( .A(n171), .ZN(n432) );
  AOI22_X1 U325 ( .A1(n29), .A2(CNT_MUL[5]), .B1(n26), .B2(N513), .ZN(n171) );
  INV_X1 U326 ( .A(n172), .ZN(n433) );
  AOI22_X1 U327 ( .A1(n29), .A2(CNT_MUL[4]), .B1(n26), .B2(N512), .ZN(n172) );
  INV_X1 U328 ( .A(n173), .ZN(n434) );
  AOI22_X1 U329 ( .A1(n29), .A2(CNT_MUL[3]), .B1(n26), .B2(N511), .ZN(n173) );
  INV_X1 U331 ( .A(n174), .ZN(n435) );
  AOI22_X1 U332 ( .A1(n29), .A2(CNT_MUL[2]), .B1(n26), .B2(N510), .ZN(n174) );
  INV_X1 U333 ( .A(n177), .ZN(n437) );
  AOI22_X1 U334 ( .A1(n29), .A2(CNT_MUL[0]), .B1(n26), .B2(N508), .ZN(n177) );
  CLKBUF_X1 U336 ( .A(n44), .Z(n38) );
  CLKBUF_X1 U337 ( .A(n44), .Z(n39) );
  CLKBUF_X1 U338 ( .A(n44), .Z(n40) );
  CLKBUF_X1 U339 ( .A(n44), .Z(n41) );
  CLKBUF_X1 U340 ( .A(n44), .Z(n42) );
  CLKBUF_X1 U341 ( .A(n44), .Z(n43) );
  INV_X1 U342 ( .A(RST), .ZN(n44) );
  INV_X1 U344 ( .A(n449), .ZN(n45) );
  NAND3_X1 U345 ( .A1(n50), .A2(n51), .A3(n45), .ZN(n117) );
  NAND3_X1 U346 ( .A1(n445), .A2(n117), .A3(n24), .ZN(STALL) );
  OAI21_X1 U347 ( .B1(n51), .B2(n449), .A(n50), .ZN(n46) );
  INV_X1 U348 ( .A(n46), .ZN(MUX_B[0]) );
  NAND2_X1 U349 ( .A1(n450), .A2(n52), .ZN(n47) );
  NAND2_X1 U350 ( .A1(n49), .A2(n47), .ZN(MUX_A[0]) );
  NAND2_X1 U351 ( .A1(n450), .A2(n53), .ZN(n48) );
  NAND2_X1 U352 ( .A1(n49), .A2(n48), .ZN(MUX_A[1]) );
  NAND2_X1 U353 ( .A1(n237), .A2(n2), .ZN(n97) );
  INV_X1 U354 ( .A(n117), .ZN(n56) );
  OAI21_X1 U355 ( .B1(n56), .B2(n249), .A(n248), .ZN(n66) );
  AOI22_X1 U356 ( .A1(CMP_A_MEM), .A2(n288), .B1(CMP_A_EXE), .B2(n66), .ZN(
        n109) );
  INV_X1 U357 ( .A(n97), .ZN(n105) );
  NAND2_X1 U358 ( .A1(n7), .A2(n105), .ZN(n107) );
  OAI211_X1 U359 ( .C1(n109), .C2(n251), .A(n107), .B(n24), .ZN(N380) );
  INV_X1 U360 ( .A(n51), .ZN(n111) );
  NAND2_X1 U361 ( .A1(n111), .A2(n25), .ZN(n113) );
  NAND3_X1 U362 ( .A1(n234), .A2(n117), .A3(n113), .ZN(N439) );
  NAND2_X1 U363 ( .A1(n21), .A2(n25), .ZN(n119) );
  OAI211_X1 U364 ( .C1(n240), .C2(n232), .A(n119), .B(n117), .ZN(N438) );
  NOR3_X1 U365 ( .A1(CNT_MUL[0]), .A2(CNT_MUL[11]), .A3(CNT_MUL[10]), .ZN(n132) );
  NOR4_X1 U366 ( .A1(CNT_MUL[15]), .A2(CNT_MUL[14]), .A3(CNT_MUL[13]), .A4(
        CNT_MUL[12]), .ZN(n130) );
  NOR4_X1 U367 ( .A1(CNT_MUL[19]), .A2(CNT_MUL[18]), .A3(CNT_MUL[17]), .A4(
        CNT_MUL[16]), .ZN(n128) );
  NOR4_X1 U368 ( .A1(CNT_MUL[22]), .A2(CNT_MUL[21]), .A3(CNT_MUL[20]), .A4(
        CNT_MUL[1]), .ZN(n126) );
  AND4_X1 U369 ( .A1(n132), .A2(n130), .A3(n128), .A4(n126), .ZN(n236) );
  NOR4_X1 U370 ( .A1(CNT_MUL[26]), .A2(CNT_MUL[25]), .A3(CNT_MUL[24]), .A4(
        CNT_MUL[23]), .ZN(n211) );
  NOR4_X1 U371 ( .A1(CNT_MUL[2]), .A2(CNT_MUL[29]), .A3(CNT_MUL[28]), .A4(
        CNT_MUL[27]), .ZN(n210) );
  NOR4_X1 U372 ( .A1(CNT_MUL[5]), .A2(CNT_MUL[4]), .A3(CNT_MUL[3]), .A4(
        CNT_MUL[30]), .ZN(n136) );
  NOR4_X1 U373 ( .A1(CNT_MUL[9]), .A2(CNT_MUL[8]), .A3(CNT_MUL[7]), .A4(
        CNT_MUL[6]), .ZN(n134) );
  AND4_X1 U374 ( .A1(n211), .A2(n210), .A3(n136), .A4(n134), .ZN(n235) );
  AOI21_X1 U375 ( .B1(n236), .B2(n235), .A(CNT_MUL[31]), .ZN(N341) );
  NOR3_X1 U376 ( .A1(CNT_DIV[0]), .A2(CNT_DIV[11]), .A3(CNT_DIV[10]), .ZN(n254) );
  NOR4_X1 U377 ( .A1(CNT_DIV[15]), .A2(CNT_DIV[14]), .A3(CNT_DIV[13]), .A4(
        CNT_DIV[12]), .ZN(n243) );
  NOR4_X1 U378 ( .A1(CNT_DIV[19]), .A2(CNT_DIV[18]), .A3(CNT_DIV[17]), .A4(
        CNT_DIV[16]), .ZN(n242) );
  NOR4_X1 U379 ( .A1(CNT_DIV[22]), .A2(CNT_DIV[21]), .A3(CNT_DIV[20]), .A4(
        CNT_DIV[1]), .ZN(n241) );
  AND4_X1 U380 ( .A1(n254), .A2(n243), .A3(n242), .A4(n241), .ZN(n289) );
  NOR4_X1 U381 ( .A1(CNT_DIV[26]), .A2(CNT_DIV[25]), .A3(CNT_DIV[24]), .A4(
        CNT_DIV[23]), .ZN(n260) );
  NOR4_X1 U382 ( .A1(CNT_DIV[2]), .A2(CNT_DIV[29]), .A3(CNT_DIV[28]), .A4(
        CNT_DIV[27]), .ZN(n259) );
  NOR4_X1 U383 ( .A1(CNT_DIV[5]), .A2(CNT_DIV[4]), .A3(CNT_DIV[3]), .A4(
        CNT_DIV[30]), .ZN(n258) );
  NOR4_X1 U384 ( .A1(CNT_DIV[9]), .A2(CNT_DIV[8]), .A3(CNT_DIV[7]), .A4(
        CNT_DIV[6]), .ZN(n255) );
  AND4_X1 U385 ( .A1(n260), .A2(n259), .A3(n258), .A4(n255), .ZN(n261) );
  AOI21_X1 U386 ( .B1(n289), .B2(n261), .A(CNT_DIV[31]), .ZN(N342) );
endmodule


module REG_N6_0 ( D, Q, EN, RST, CLK );
  input [5:0] D;
  output [5:0] Q;
  input EN, RST, CLK;
  wire   n1;

  FD_1_115 FF_0 ( .D(D[0]), .CLK(CLK), .EN(n1), .RST(RST), .Q(Q[0]) );
  FD_1_114 FF_1 ( .D(D[1]), .CLK(CLK), .EN(n1), .RST(RST), .Q(Q[1]) );
  FD_1_113 FF_2 ( .D(D[2]), .CLK(CLK), .EN(n1), .RST(RST), .Q(Q[2]) );
  FD_1_112 FF_3 ( .D(D[3]), .CLK(CLK), .EN(n1), .RST(RST), .Q(Q[3]) );
  FD_1_111 FF_4 ( .D(D[4]), .CLK(CLK), .EN(n1), .RST(RST), .Q(Q[4]) );
  FD_1_110 FF_5 ( .D(D[5]), .CLK(CLK), .EN(n1), .RST(RST), .Q(Q[5]) );
  BUF_X1 U1 ( .A(EN), .Z(n1) );
endmodule


module EQU_COMPARATOR_N5_0 ( A, B, Y );
  input [4:0] A;
  input [4:0] B;
  output Y;

  wire   [4:0] L;

  XNOR_GATE_0 XNORING_0 ( .A(A[0]), .B(B[0]), .Y(L[0]) );
  XNOR_GATE_217 XNORING_1 ( .A(A[1]), .B(B[1]), .Y(L[1]) );
  XNOR_GATE_216 XNORING_2 ( .A(A[2]), .B(B[2]), .Y(L[2]) );
  XNOR_GATE_215 XNORING_3 ( .A(A[3]), .B(B[3]), .Y(L[3]) );
  XNOR_GATE_214 XNORING_4 ( .A(A[4]), .B(B[4]), .Y(L[4]) );
  N_AND_N5_0 ANDING ( .A(L), .Y(Y) );
endmodule


module ALU_N32_ALU_SIZE5 ( IN_A, IN_B, ALU_OP_CODE, CLK, RST, RST_DIV, OUT_ALU
 );
  input [31:0] IN_A;
  input [31:0] IN_B;
  input [4:0] ALU_OP_CODE;
  output [31:0] OUT_ALU;
  input CLK, RST, RST_DIV;
  wire   UNSIGN, SUB_ADD, MUX_SEL_ADD_S, RIGHT_LEFT, ARITH_LOG, EN_GUARD_CMP,
         EN_GUARD_LOG, EN_GUARD_P4, SIGN_SIG, Ci_P4, Co_ADDER, Co_CMP,
         UNSIGN_CMP, MSB_A_CMP, MSB_B_CMP, OUT_DIV_SIGN, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n42, n43, n44, n46, n47, n48,
         n49, n50, n51, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n41, n45, n52, n53;
  wire   [2:0] LOG_OP;
  wire   [2:0] CMP_OP;
  wire   [2:0] MUX_SEL;
  wire   [15:0] OUT_DIV_D;
  wire   [15:0] OUT_DIV_R;
  wire   [31:0] IN_A_P4;
  wire   [31:0] A_SIG;
  wire   [31:0] IN_B_P4;
  wire   [31:0] B_SIG;
  wire   [31:0] B_SIG2;
  wire   [31:0] OUT_P4;
  wire   [31:0] S_CMP;
  wire   [31:0] OUT_CMP;
  wire   [31:0] A_LOG;
  wire   [31:0] B_LOG;
  wire   [3:0] LOG_OP_SIG;
  wire   [31:0] OUT_LOG;
  wire   [31:0] OUT_SHIFT;
  wire   [31:0] OUT_MUL;
  wire   [31:0] OUT_DIV;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  NAND3_X1 U40 ( .A1(n21), .A2(n16), .A3(n17), .ZN(RIGHT_LEFT) );
  NAND2_X1 U41 ( .A1(n38), .A2(n22), .ZN(n26) );
  NAND2_X1 U42 ( .A1(n34), .A2(n38), .ZN(n20) );
  NAND2_X1 U43 ( .A1(n39), .A2(LOG_OP[2]), .ZN(LOG_OP[0]) );
  NAND2_X1 U44 ( .A1(n29), .A2(n22), .ZN(LOG_OP[2]) );
  NAND2_X1 U45 ( .A1(n40), .A2(n52), .ZN(EN_GUARD_P4) );
  NAND3_X1 U46 ( .A1(n42), .A2(n43), .A3(n44), .ZN(n40) );
  XOR2_X1 U47 ( .A(ALU_OP_CODE[0]), .B(n36), .Z(n44) );
  NAND3_X1 U48 ( .A1(n39), .A2(n53), .A3(n46), .ZN(EN_GUARD_LOG) );
  NAND3_X1 U49 ( .A1(n36), .A2(n43), .A3(n22), .ZN(n46) );
  NAND2_X1 U50 ( .A1(n30), .A2(n34), .ZN(n39) );
  NAND3_X1 U51 ( .A1(n47), .A2(n18), .A3(n48), .ZN(CMP_OP[2]) );
  NAND2_X1 U52 ( .A1(ALU_OP_CODE[0]), .A2(ALU_OP_CODE[2]), .ZN(n16) );
  NAND3_X1 U53 ( .A1(n36), .A2(n37), .A3(ALU_OP_CODE[3]), .ZN(n18) );
  NAND2_X1 U54 ( .A1(n30), .A2(n22), .ZN(n47) );
  NAND2_X1 U55 ( .A1(n37), .A2(n43), .ZN(n15) );
  D_LATCH_0 LATCH_P4_A_0 ( .D(A_SIG[0]), .EN(n9), .Q(IN_A_P4[0]) );
  D_LATCH_168 LATCH_P4_B_0 ( .D(B_SIG[0]), .EN(n5), .Q(IN_B_P4[0]) );
  D_LATCH_167 LATCH_P4_A_1 ( .D(A_SIG[1]), .EN(n5), .Q(IN_A_P4[1]) );
  D_LATCH_166 LATCH_P4_B_1 ( .D(B_SIG[1]), .EN(n5), .Q(IN_B_P4[1]) );
  D_LATCH_165 LATCH_P4_A_2 ( .D(A_SIG[2]), .EN(n5), .Q(IN_A_P4[2]) );
  D_LATCH_164 LATCH_P4_B_2 ( .D(B_SIG[2]), .EN(n5), .Q(IN_B_P4[2]) );
  D_LATCH_163 LATCH_P4_A_3 ( .D(A_SIG[3]), .EN(n5), .Q(IN_A_P4[3]) );
  D_LATCH_162 LATCH_P4_B_3 ( .D(B_SIG[3]), .EN(n5), .Q(IN_B_P4[3]) );
  D_LATCH_161 LATCH_P4_A_4 ( .D(A_SIG[4]), .EN(n5), .Q(IN_A_P4[4]) );
  D_LATCH_160 LATCH_P4_B_4 ( .D(B_SIG[4]), .EN(n5), .Q(IN_B_P4[4]) );
  D_LATCH_159 LATCH_P4_A_5 ( .D(A_SIG[5]), .EN(n5), .Q(IN_A_P4[5]) );
  D_LATCH_158 LATCH_P4_B_5 ( .D(B_SIG[5]), .EN(n5), .Q(IN_B_P4[5]) );
  D_LATCH_157 LATCH_P4_A_6 ( .D(A_SIG[6]), .EN(n5), .Q(IN_A_P4[6]) );
  D_LATCH_156 LATCH_P4_B_6 ( .D(B_SIG[6]), .EN(n5), .Q(IN_B_P4[6]) );
  D_LATCH_155 LATCH_P4_A_7 ( .D(A_SIG[7]), .EN(n6), .Q(IN_A_P4[7]) );
  D_LATCH_154 LATCH_P4_B_7 ( .D(B_SIG[7]), .EN(n6), .Q(IN_B_P4[7]) );
  D_LATCH_153 LATCH_P4_A_8 ( .D(A_SIG[8]), .EN(n6), .Q(IN_A_P4[8]) );
  D_LATCH_152 LATCH_P4_B_8 ( .D(B_SIG[8]), .EN(n6), .Q(IN_B_P4[8]) );
  D_LATCH_151 LATCH_P4_A_9 ( .D(A_SIG[9]), .EN(n6), .Q(IN_A_P4[9]) );
  D_LATCH_150 LATCH_P4_B_9 ( .D(B_SIG[9]), .EN(n6), .Q(IN_B_P4[9]) );
  D_LATCH_149 LATCH_P4_A_10 ( .D(A_SIG[10]), .EN(n6), .Q(IN_A_P4[10]) );
  D_LATCH_148 LATCH_P4_B_10 ( .D(B_SIG[10]), .EN(n6), .Q(IN_B_P4[10]) );
  D_LATCH_147 LATCH_P4_A_11 ( .D(A_SIG[11]), .EN(n6), .Q(IN_A_P4[11]) );
  D_LATCH_146 LATCH_P4_B_11 ( .D(B_SIG[11]), .EN(n6), .Q(IN_B_P4[11]) );
  D_LATCH_145 LATCH_P4_A_12 ( .D(A_SIG[12]), .EN(n6), .Q(IN_A_P4[12]) );
  D_LATCH_144 LATCH_P4_B_12 ( .D(B_SIG[12]), .EN(n6), .Q(IN_B_P4[12]) );
  D_LATCH_143 LATCH_P4_A_13 ( .D(A_SIG[13]), .EN(n6), .Q(IN_A_P4[13]) );
  D_LATCH_142 LATCH_P4_B_13 ( .D(B_SIG[13]), .EN(n7), .Q(IN_B_P4[13]) );
  D_LATCH_141 LATCH_P4_A_14 ( .D(A_SIG[14]), .EN(n7), .Q(IN_A_P4[14]) );
  D_LATCH_140 LATCH_P4_B_14 ( .D(B_SIG[14]), .EN(n7), .Q(IN_B_P4[14]) );
  D_LATCH_139 LATCH_P4_A_15 ( .D(A_SIG[15]), .EN(n7), .Q(IN_A_P4[15]) );
  D_LATCH_138 LATCH_P4_B_15 ( .D(B_SIG[15]), .EN(n7), .Q(IN_B_P4[15]) );
  D_LATCH_137 LATCH_P4_A_16 ( .D(A_SIG[16]), .EN(n7), .Q(IN_A_P4[16]) );
  D_LATCH_136 LATCH_P4_B_16 ( .D(B_SIG[16]), .EN(n7), .Q(IN_B_P4[16]) );
  D_LATCH_135 LATCH_P4_A_17 ( .D(A_SIG[17]), .EN(n7), .Q(IN_A_P4[17]) );
  D_LATCH_134 LATCH_P4_B_17 ( .D(B_SIG[17]), .EN(n7), .Q(IN_B_P4[17]) );
  D_LATCH_133 LATCH_P4_A_18 ( .D(A_SIG[18]), .EN(n7), .Q(IN_A_P4[18]) );
  D_LATCH_132 LATCH_P4_B_18 ( .D(B_SIG[18]), .EN(n7), .Q(IN_B_P4[18]) );
  D_LATCH_131 LATCH_P4_A_19 ( .D(A_SIG[19]), .EN(n7), .Q(IN_A_P4[19]) );
  D_LATCH_130 LATCH_P4_B_19 ( .D(B_SIG[19]), .EN(n7), .Q(IN_B_P4[19]) );
  D_LATCH_129 LATCH_P4_A_20 ( .D(A_SIG[20]), .EN(n8), .Q(IN_A_P4[20]) );
  D_LATCH_128 LATCH_P4_B_20 ( .D(B_SIG[20]), .EN(n8), .Q(IN_B_P4[20]) );
  D_LATCH_127 LATCH_P4_A_21 ( .D(A_SIG[21]), .EN(n8), .Q(IN_A_P4[21]) );
  D_LATCH_126 LATCH_P4_B_21 ( .D(B_SIG[21]), .EN(n8), .Q(IN_B_P4[21]) );
  D_LATCH_125 LATCH_P4_A_22 ( .D(A_SIG[22]), .EN(n8), .Q(IN_A_P4[22]) );
  D_LATCH_124 LATCH_P4_B_22 ( .D(B_SIG[22]), .EN(n8), .Q(IN_B_P4[22]) );
  D_LATCH_123 LATCH_P4_A_23 ( .D(A_SIG[23]), .EN(n8), .Q(IN_A_P4[23]) );
  D_LATCH_122 LATCH_P4_B_23 ( .D(B_SIG[23]), .EN(n8), .Q(IN_B_P4[23]) );
  D_LATCH_121 LATCH_P4_A_24 ( .D(A_SIG[24]), .EN(n8), .Q(IN_A_P4[24]) );
  D_LATCH_120 LATCH_P4_B_24 ( .D(B_SIG[24]), .EN(n8), .Q(IN_B_P4[24]) );
  D_LATCH_119 LATCH_P4_A_25 ( .D(A_SIG[25]), .EN(n8), .Q(IN_A_P4[25]) );
  D_LATCH_118 LATCH_P4_B_25 ( .D(B_SIG[25]), .EN(n8), .Q(IN_B_P4[25]) );
  D_LATCH_117 LATCH_P4_A_26 ( .D(A_SIG[26]), .EN(n8), .Q(IN_A_P4[26]) );
  D_LATCH_116 LATCH_P4_B_26 ( .D(B_SIG[26]), .EN(n9), .Q(IN_B_P4[26]) );
  D_LATCH_115 LATCH_P4_A_27 ( .D(A_SIG[27]), .EN(n9), .Q(IN_A_P4[27]) );
  D_LATCH_114 LATCH_P4_B_27 ( .D(B_SIG[27]), .EN(n9), .Q(IN_B_P4[27]) );
  D_LATCH_113 LATCH_P4_A_28 ( .D(A_SIG[28]), .EN(n9), .Q(IN_A_P4[28]) );
  D_LATCH_112 LATCH_P4_B_28 ( .D(B_SIG[28]), .EN(n9), .Q(IN_B_P4[28]) );
  D_LATCH_111 LATCH_P4_A_29 ( .D(A_SIG[29]), .EN(n9), .Q(IN_A_P4[29]) );
  D_LATCH_110 LATCH_P4_B_29 ( .D(B_SIG[29]), .EN(n9), .Q(IN_B_P4[29]) );
  D_LATCH_109 LATCH_P4_A_30 ( .D(A_SIG[30]), .EN(n9), .Q(IN_A_P4[30]) );
  D_LATCH_108 LATCH_P4_B_30 ( .D(B_SIG[30]), .EN(n9), .Q(IN_B_P4[30]) );
  D_LATCH_107 LATCH_P4_A_31 ( .D(A_SIG[31]), .EN(n9), .Q(IN_A_P4[31]) );
  D_LATCH_106 LATCH_P4_B_31 ( .D(B_SIG[31]), .EN(n9), .Q(IN_B_P4[31]) );
  D_LATCH_105 EVAL_P4_Ci ( .D(n3), .EN(n9), .Q(Ci_P4) );
  XOR_GATE_1_0 XORS_0 ( .A(IN_B_P4[0]), .B(n3), .Y(B_SIG2[0]) );
  XOR_GATE_1_669 XORS_1 ( .A(IN_B_P4[1]), .B(n3), .Y(B_SIG2[1]) );
  XOR_GATE_1_668 XORS_2 ( .A(IN_B_P4[2]), .B(n4), .Y(B_SIG2[2]) );
  XOR_GATE_1_667 XORS_3 ( .A(IN_B_P4[3]), .B(n4), .Y(B_SIG2[3]) );
  XOR_GATE_1_666 XORS_4 ( .A(IN_B_P4[4]), .B(n4), .Y(B_SIG2[4]) );
  XOR_GATE_1_665 XORS_5 ( .A(IN_B_P4[5]), .B(n4), .Y(B_SIG2[5]) );
  XOR_GATE_1_664 XORS_6 ( .A(IN_B_P4[6]), .B(n4), .Y(B_SIG2[6]) );
  XOR_GATE_1_663 XORS_7 ( .A(IN_B_P4[7]), .B(n4), .Y(B_SIG2[7]) );
  XOR_GATE_1_662 XORS_8 ( .A(IN_B_P4[8]), .B(n4), .Y(B_SIG2[8]) );
  XOR_GATE_1_661 XORS_9 ( .A(IN_B_P4[9]), .B(n4), .Y(B_SIG2[9]) );
  XOR_GATE_1_660 XORS_10 ( .A(IN_B_P4[10]), .B(n4), .Y(B_SIG2[10]) );
  XOR_GATE_1_659 XORS_11 ( .A(IN_B_P4[11]), .B(n4), .Y(B_SIG2[11]) );
  XOR_GATE_1_658 XORS_12 ( .A(IN_B_P4[12]), .B(n4), .Y(B_SIG2[12]) );
  XOR_GATE_1_657 XORS_13 ( .A(IN_B_P4[13]), .B(n4), .Y(B_SIG2[13]) );
  XOR_GATE_1_656 XORS_14 ( .A(IN_B_P4[14]), .B(n4), .Y(B_SIG2[14]) );
  XOR_GATE_1_655 XORS_15 ( .A(IN_B_P4[15]), .B(n4), .Y(B_SIG2[15]) );
  XOR_GATE_1_654 XORS_16 ( .A(IN_B_P4[16]), .B(n4), .Y(B_SIG2[16]) );
  XOR_GATE_1_653 XORS_17 ( .A(IN_B_P4[17]), .B(n3), .Y(B_SIG2[17]) );
  XOR_GATE_1_652 XORS_18 ( .A(IN_B_P4[18]), .B(n3), .Y(B_SIG2[18]) );
  XOR_GATE_1_651 XORS_19 ( .A(IN_B_P4[19]), .B(n3), .Y(B_SIG2[19]) );
  XOR_GATE_1_650 XORS_20 ( .A(IN_B_P4[20]), .B(n3), .Y(B_SIG2[20]) );
  XOR_GATE_1_649 XORS_21 ( .A(IN_B_P4[21]), .B(n3), .Y(B_SIG2[21]) );
  XOR_GATE_1_648 XORS_22 ( .A(IN_B_P4[22]), .B(n3), .Y(B_SIG2[22]) );
  XOR_GATE_1_647 XORS_23 ( .A(IN_B_P4[23]), .B(n3), .Y(B_SIG2[23]) );
  XOR_GATE_1_646 XORS_24 ( .A(IN_B_P4[24]), .B(n3), .Y(B_SIG2[24]) );
  XOR_GATE_1_645 XORS_25 ( .A(IN_B_P4[25]), .B(n3), .Y(B_SIG2[25]) );
  XOR_GATE_1_644 XORS_26 ( .A(IN_B_P4[26]), .B(n3), .Y(B_SIG2[26]) );
  XOR_GATE_1_643 XORS_27 ( .A(IN_B_P4[27]), .B(n3), .Y(B_SIG2[27]) );
  XOR_GATE_1_642 XORS_28 ( .A(IN_B_P4[28]), .B(n3), .Y(B_SIG2[28]) );
  XOR_GATE_1_641 XORS_29 ( .A(IN_B_P4[29]), .B(n3), .Y(B_SIG2[29]) );
  XOR_GATE_1_640 XORS_30 ( .A(IN_B_P4[30]), .B(n3), .Y(B_SIG2[30]) );
  XOR_GATE_1_639 XORS_31 ( .A(IN_B_P4[31]), .B(n3), .Y(B_SIG2[31]) );
  P4_ADDER_N32 ADDER_INST ( .A(IN_A_P4), .B(B_SIG2), .Ci(Ci_P4), .Co(Co_ADDER), 
        .S(OUT_P4) );
  D_LATCH_104 LATCH_CMP_0 ( .D(OUT_P4[0]), .EN(n45), .Q(S_CMP[0]) );
  D_LATCH_103 LATCH_CMP_1 ( .D(OUT_P4[1]), .EN(n45), .Q(S_CMP[1]) );
  D_LATCH_102 LATCH_CMP_2 ( .D(OUT_P4[2]), .EN(n45), .Q(S_CMP[2]) );
  D_LATCH_101 LATCH_CMP_3 ( .D(OUT_P4[3]), .EN(n45), .Q(S_CMP[3]) );
  D_LATCH_100 LATCH_CMP_4 ( .D(OUT_P4[4]), .EN(n45), .Q(S_CMP[4]) );
  D_LATCH_99 LATCH_CMP_5 ( .D(OUT_P4[5]), .EN(n45), .Q(S_CMP[5]) );
  D_LATCH_98 LATCH_CMP_6 ( .D(OUT_P4[6]), .EN(n45), .Q(S_CMP[6]) );
  D_LATCH_97 LATCH_CMP_7 ( .D(OUT_P4[7]), .EN(n45), .Q(S_CMP[7]) );
  D_LATCH_96 LATCH_CMP_8 ( .D(OUT_P4[8]), .EN(n45), .Q(S_CMP[8]) );
  D_LATCH_95 LATCH_CMP_9 ( .D(OUT_P4[9]), .EN(n45), .Q(S_CMP[9]) );
  D_LATCH_94 LATCH_CMP_10 ( .D(OUT_P4[10]), .EN(n45), .Q(S_CMP[10]) );
  D_LATCH_93 LATCH_CMP_11 ( .D(OUT_P4[11]), .EN(n45), .Q(S_CMP[11]) );
  D_LATCH_92 LATCH_CMP_12 ( .D(OUT_P4[12]), .EN(n45), .Q(S_CMP[12]) );
  D_LATCH_91 LATCH_CMP_13 ( .D(OUT_P4[13]), .EN(n45), .Q(S_CMP[13]) );
  D_LATCH_90 LATCH_CMP_14 ( .D(OUT_P4[14]), .EN(n45), .Q(S_CMP[14]) );
  D_LATCH_89 LATCH_CMP_15 ( .D(OUT_P4[15]), .EN(n45), .Q(S_CMP[15]) );
  D_LATCH_88 LATCH_CMP_16 ( .D(OUT_P4[16]), .EN(n45), .Q(S_CMP[16]) );
  D_LATCH_87 LATCH_CMP_17 ( .D(OUT_P4[17]), .EN(n45), .Q(S_CMP[17]) );
  D_LATCH_86 LATCH_CMP_18 ( .D(OUT_P4[18]), .EN(n45), .Q(S_CMP[18]) );
  D_LATCH_85 LATCH_CMP_19 ( .D(OUT_P4[19]), .EN(n45), .Q(S_CMP[19]) );
  D_LATCH_84 LATCH_CMP_20 ( .D(OUT_P4[20]), .EN(n45), .Q(S_CMP[20]) );
  D_LATCH_83 LATCH_CMP_21 ( .D(OUT_P4[21]), .EN(n45), .Q(S_CMP[21]) );
  D_LATCH_82 LATCH_CMP_22 ( .D(OUT_P4[22]), .EN(n45), .Q(S_CMP[22]) );
  D_LATCH_81 LATCH_CMP_23 ( .D(OUT_P4[23]), .EN(n45), .Q(S_CMP[23]) );
  D_LATCH_80 LATCH_CMP_24 ( .D(OUT_P4[24]), .EN(n45), .Q(S_CMP[24]) );
  D_LATCH_79 LATCH_CMP_25 ( .D(OUT_P4[25]), .EN(n45), .Q(S_CMP[25]) );
  D_LATCH_78 LATCH_CMP_26 ( .D(OUT_P4[26]), .EN(n45), .Q(S_CMP[26]) );
  D_LATCH_77 LATCH_CMP_27 ( .D(OUT_P4[27]), .EN(n45), .Q(S_CMP[27]) );
  D_LATCH_76 LATCH_CMP_28 ( .D(OUT_P4[28]), .EN(n45), .Q(S_CMP[28]) );
  D_LATCH_75 LATCH_CMP_29 ( .D(OUT_P4[29]), .EN(n45), .Q(S_CMP[29]) );
  D_LATCH_74 LATCH_CMP_30 ( .D(OUT_P4[30]), .EN(EN_GUARD_CMP), .Q(S_CMP[30])
         );
  D_LATCH_73 LATCH_CMP_31 ( .D(OUT_P4[31]), .EN(n45), .Q(S_CMP[31]) );
  D_LATCH_72 EVAL_CMP_Co ( .D(Co_ADDER), .EN(EN_GUARD_CMP), .Q(Co_CMP) );
  D_LATCH_71 EVAL_CMP_UNSIGN ( .D(UNSIGN), .EN(n45), .Q(UNSIGN_CMP) );
  D_LATCH_70 EVAL_CMP_MSB_A ( .D(IN_A[31]), .EN(EN_GUARD_CMP), .Q(MSB_A_CMP)
         );
  D_LATCH_69 EVAL_CMP_MSB_B ( .D(IN_B[31]), .EN(n45), .Q(MSB_B_CMP) );
  CMP_N32 CMP_INST ( .C(Co_CMP), .S(S_CMP), .OP_SEL(CMP_OP), .UNSIGN(
        UNSIGN_CMP), .MSB_A(MSB_A_CMP), .MSB_B(MSB_B_CMP), .Y({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, OUT_CMP[0]}) );
  D_LATCH_68 LATCH_LOG_1_0 ( .D(IN_A[0]), .EN(n10), .Q(A_LOG[0]) );
  D_LATCH_67 LATCH_LOG_2_0 ( .D(IN_B[0]), .EN(n10), .Q(B_LOG[0]) );
  D_LATCH_66 LATCH_LOG_1_1 ( .D(n1), .EN(n10), .Q(A_LOG[1]) );
  D_LATCH_65 LATCH_LOG_2_1 ( .D(n2), .EN(n10), .Q(B_LOG[1]) );
  D_LATCH_64 LATCH_LOG_1_2 ( .D(IN_A[2]), .EN(n10), .Q(A_LOG[2]) );
  D_LATCH_63 LATCH_LOG_2_2 ( .D(IN_B[2]), .EN(n10), .Q(B_LOG[2]) );
  D_LATCH_62 LATCH_LOG_1_3 ( .D(IN_A[3]), .EN(n10), .Q(A_LOG[3]) );
  D_LATCH_61 LATCH_LOG_2_3 ( .D(IN_B[3]), .EN(n10), .Q(B_LOG[3]) );
  D_LATCH_60 LATCH_LOG_1_4 ( .D(IN_A[4]), .EN(n10), .Q(A_LOG[4]) );
  D_LATCH_59 LATCH_LOG_2_4 ( .D(IN_B[4]), .EN(n10), .Q(B_LOG[4]) );
  D_LATCH_58 LATCH_LOG_1_5 ( .D(IN_A[5]), .EN(n10), .Q(A_LOG[5]) );
  D_LATCH_57 LATCH_LOG_2_5 ( .D(IN_B[5]), .EN(n10), .Q(B_LOG[5]) );
  D_LATCH_56 LATCH_LOG_1_6 ( .D(IN_A[6]), .EN(n10), .Q(A_LOG[6]) );
  D_LATCH_55 LATCH_LOG_2_6 ( .D(IN_B[6]), .EN(n11), .Q(B_LOG[6]) );
  D_LATCH_54 LATCH_LOG_1_7 ( .D(IN_A[7]), .EN(n11), .Q(A_LOG[7]) );
  D_LATCH_53 LATCH_LOG_2_7 ( .D(IN_B[7]), .EN(n11), .Q(B_LOG[7]) );
  D_LATCH_52 LATCH_LOG_1_8 ( .D(IN_A[8]), .EN(n11), .Q(A_LOG[8]) );
  D_LATCH_51 LATCH_LOG_2_8 ( .D(IN_B[8]), .EN(n11), .Q(B_LOG[8]) );
  D_LATCH_50 LATCH_LOG_1_9 ( .D(IN_A[9]), .EN(n11), .Q(A_LOG[9]) );
  D_LATCH_49 LATCH_LOG_2_9 ( .D(IN_B[9]), .EN(n11), .Q(B_LOG[9]) );
  D_LATCH_48 LATCH_LOG_1_10 ( .D(IN_A[10]), .EN(n11), .Q(A_LOG[10]) );
  D_LATCH_47 LATCH_LOG_2_10 ( .D(IN_B[10]), .EN(n11), .Q(B_LOG[10]) );
  D_LATCH_46 LATCH_LOG_1_11 ( .D(IN_A[11]), .EN(n11), .Q(A_LOG[11]) );
  D_LATCH_45 LATCH_LOG_2_11 ( .D(IN_B[11]), .EN(n11), .Q(B_LOG[11]) );
  D_LATCH_44 LATCH_LOG_1_12 ( .D(IN_A[12]), .EN(n11), .Q(A_LOG[12]) );
  D_LATCH_43 LATCH_LOG_2_12 ( .D(IN_B[12]), .EN(n11), .Q(B_LOG[12]) );
  D_LATCH_42 LATCH_LOG_1_13 ( .D(IN_A[13]), .EN(n12), .Q(A_LOG[13]) );
  D_LATCH_41 LATCH_LOG_2_13 ( .D(IN_B[13]), .EN(n12), .Q(B_LOG[13]) );
  D_LATCH_40 LATCH_LOG_1_14 ( .D(IN_A[14]), .EN(n12), .Q(A_LOG[14]) );
  D_LATCH_39 LATCH_LOG_2_14 ( .D(IN_B[14]), .EN(n12), .Q(B_LOG[14]) );
  D_LATCH_38 LATCH_LOG_1_15 ( .D(IN_A[15]), .EN(n12), .Q(A_LOG[15]) );
  D_LATCH_37 LATCH_LOG_2_15 ( .D(IN_B[15]), .EN(n12), .Q(B_LOG[15]) );
  D_LATCH_36 LATCH_LOG_1_16 ( .D(IN_A[16]), .EN(n12), .Q(A_LOG[16]) );
  D_LATCH_35 LATCH_LOG_2_16 ( .D(IN_B[16]), .EN(n12), .Q(B_LOG[16]) );
  D_LATCH_34 LATCH_LOG_1_17 ( .D(IN_A[17]), .EN(n12), .Q(A_LOG[17]) );
  D_LATCH_33 LATCH_LOG_2_17 ( .D(IN_B[17]), .EN(n12), .Q(B_LOG[17]) );
  D_LATCH_32 LATCH_LOG_1_18 ( .D(IN_A[18]), .EN(n12), .Q(A_LOG[18]) );
  D_LATCH_31 LATCH_LOG_2_18 ( .D(IN_B[18]), .EN(n12), .Q(B_LOG[18]) );
  D_LATCH_30 LATCH_LOG_1_19 ( .D(IN_A[19]), .EN(n12), .Q(A_LOG[19]) );
  D_LATCH_29 LATCH_LOG_2_19 ( .D(IN_B[19]), .EN(n13), .Q(B_LOG[19]) );
  D_LATCH_28 LATCH_LOG_1_20 ( .D(IN_A[20]), .EN(n13), .Q(A_LOG[20]) );
  D_LATCH_27 LATCH_LOG_2_20 ( .D(IN_B[20]), .EN(n13), .Q(B_LOG[20]) );
  D_LATCH_26 LATCH_LOG_1_21 ( .D(IN_A[21]), .EN(n13), .Q(A_LOG[21]) );
  D_LATCH_25 LATCH_LOG_2_21 ( .D(IN_B[21]), .EN(n13), .Q(B_LOG[21]) );
  D_LATCH_24 LATCH_LOG_1_22 ( .D(IN_A[22]), .EN(n13), .Q(A_LOG[22]) );
  D_LATCH_23 LATCH_LOG_2_22 ( .D(IN_B[22]), .EN(n13), .Q(B_LOG[22]) );
  D_LATCH_22 LATCH_LOG_1_23 ( .D(IN_A[23]), .EN(n13), .Q(A_LOG[23]) );
  D_LATCH_21 LATCH_LOG_2_23 ( .D(IN_B[23]), .EN(n13), .Q(B_LOG[23]) );
  D_LATCH_20 LATCH_LOG_1_24 ( .D(IN_A[24]), .EN(n13), .Q(A_LOG[24]) );
  D_LATCH_19 LATCH_LOG_2_24 ( .D(IN_B[24]), .EN(n13), .Q(B_LOG[24]) );
  D_LATCH_18 LATCH_LOG_1_25 ( .D(IN_A[25]), .EN(n13), .Q(A_LOG[25]) );
  D_LATCH_17 LATCH_LOG_2_25 ( .D(IN_B[25]), .EN(n13), .Q(B_LOG[25]) );
  D_LATCH_16 LATCH_LOG_1_26 ( .D(IN_A[26]), .EN(n14), .Q(A_LOG[26]) );
  D_LATCH_15 LATCH_LOG_2_26 ( .D(IN_B[26]), .EN(n14), .Q(B_LOG[26]) );
  D_LATCH_14 LATCH_LOG_1_27 ( .D(IN_A[27]), .EN(n14), .Q(A_LOG[27]) );
  D_LATCH_13 LATCH_LOG_2_27 ( .D(IN_B[27]), .EN(n14), .Q(B_LOG[27]) );
  D_LATCH_12 LATCH_LOG_1_28 ( .D(IN_A[28]), .EN(n14), .Q(A_LOG[28]) );
  D_LATCH_11 LATCH_LOG_2_28 ( .D(IN_B[28]), .EN(n14), .Q(B_LOG[28]) );
  D_LATCH_10 LATCH_LOG_1_29 ( .D(IN_A[29]), .EN(n14), .Q(A_LOG[29]) );
  D_LATCH_9 LATCH_LOG_2_29 ( .D(IN_B[29]), .EN(n14), .Q(B_LOG[29]) );
  D_LATCH_8 LATCH_LOG_1_30 ( .D(IN_A[30]), .EN(n14), .Q(A_LOG[30]) );
  D_LATCH_7 LATCH_LOG_2_30 ( .D(IN_B[30]), .EN(n14), .Q(B_LOG[30]) );
  D_LATCH_6 LATCH_LOG_1_31 ( .D(IN_A[31]), .EN(n14), .Q(A_LOG[31]) );
  D_LATCH_5 LATCH_LOG_2_31 ( .D(IN_B[31]), .EN(n14), .Q(B_LOG[31]) );
  D_LATCH_4 LATCH_LOG_3_0 ( .D(LOG_OP[0]), .EN(n14), .Q(LOG_OP_SIG[0]) );
  D_LATCH_3 LATCH_LOG_3_1 ( .D(LOG_OP[2]), .EN(n41), .Q(LOG_OP_SIG[1]) );
  D_LATCH_2 LATCH_LOG_3_2 ( .D(LOG_OP[2]), .EN(n41), .Q(LOG_OP_SIG[2]) );
  D_LATCH_1 LATCH_LOG_3_3 ( .D(1'b0), .EN(n41), .Q(LOG_OP_SIG[3]) );
  T2_LOGICALS_N32 LOG_INST ( .OP(LOG_OP_SIG), .A(A_LOG), .B(B_LOG), .Y(OUT_LOG) );
  T2_SHIFTER_N32 SHIFT_INST ( .A({IN_A[31:2], n1, IN_A[0]}), .B({IN_B[4:2], n2, 
        IN_B[0]}), .ARITH_LOG(ARITH_LOG), .RIGHT_LEFT(RIGHT_LEFT), .Y(
        OUT_SHIFT) );
  BOOTHMUL MULT_INST ( .A(IN_A[15:0]), .B(IN_B[15:0]), .CLK(CLK), .EN(1'b1), 
        .RST(RST), .P(OUT_MUL) );
  NR_DIVISOR DIVISOR_INST ( .CLK(CLK), .RST(RST_DIV), .EN(1'b1), .Z({
        IN_A[15:2], n1, IN_A[0]}), .D({IN_B[15:2], n2, IN_B[0]}), .Q(
        OUT_DIV[15:0]), .R(OUT_DIV[31:16]), .ADD_IN_D(OUT_DIV_D), .ADD_IN_R(
        OUT_DIV_R), .SIGN(OUT_DIV_SIGN), .ADD_OUT(OUT_P4[15:0]) );
  MUX21_GEN_N32_2 MUX_IN_A ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, OUT_DIV_R}), .B(
        {IN_A[31:2], n1, IN_A[0]}), .SEL(MUX_SEL_ADD_S), .Y(A_SIG) );
  MUX21_GEN_N32_1 MUXING_IN_B ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, OUT_DIV_D}), .B(
        {IN_B[31:2], n2, IN_B[0]}), .SEL(MUX_SEL_ADD_S), .Y(B_SIG) );
  MUX21_6 MUXING_IN_S ( .A(OUT_DIV_SIGN), .B(SUB_ADD), .S(MUX_SEL_ADD_S), .Y(
        SIGN_SIG) );
  MUX61_GEN_N32 MUXING ( .A(OUT_P4), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, OUT_CMP[0]}), .C(OUT_LOG), .D(OUT_SHIFT), .E(OUT_MUL), .F(
        OUT_DIV), .SEL(MUX_SEL), .Y(OUT_ALU) );
  CLKBUF_X1 U3 ( .A(IN_A[1]), .Z(n1) );
  CLKBUF_X1 U4 ( .A(IN_B[1]), .Z(n2) );
  INV_X1 U5 ( .A(LOG_OP[0]), .ZN(n32) );
  BUF_X1 U6 ( .A(SIGN_SIG), .Z(n3) );
  BUF_X1 U7 ( .A(SIGN_SIG), .Z(n4) );
  BUF_X1 U8 ( .A(EN_GUARD_LOG), .Z(n10) );
  BUF_X1 U9 ( .A(EN_GUARD_LOG), .Z(n11) );
  BUF_X1 U10 ( .A(EN_GUARD_LOG), .Z(n12) );
  BUF_X1 U11 ( .A(EN_GUARD_LOG), .Z(n13) );
  BUF_X1 U12 ( .A(EN_GUARD_LOG), .Z(n14) );
  AOI21_X1 U13 ( .B1(n33), .B2(n49), .A(n50), .ZN(CMP_OP[1]) );
  INV_X1 U14 ( .A(n47), .ZN(n50) );
  AND3_X1 U15 ( .A1(n31), .A2(n32), .A3(n26), .ZN(MUX_SEL[1]) );
  AND2_X1 U16 ( .A1(n24), .A2(n22), .ZN(MUX_SEL_ADD_S) );
  NOR2_X1 U17 ( .A1(n22), .A2(n23), .ZN(n17) );
  BUF_X1 U18 ( .A(EN_GUARD_P4), .Z(n5) );
  BUF_X1 U19 ( .A(EN_GUARD_P4), .Z(n6) );
  BUF_X1 U20 ( .A(EN_GUARD_P4), .Z(n7) );
  BUF_X1 U21 ( .A(EN_GUARD_P4), .Z(n8) );
  BUF_X1 U22 ( .A(EN_GUARD_P4), .Z(n9) );
  AOI221_X1 U23 ( .B1(n33), .B2(n21), .C1(n34), .C2(n21), .A(ARITH_LOG), .ZN(
        n31) );
  OAI22_X1 U24 ( .A1(n15), .A2(n16), .B1(n17), .B2(n18), .ZN(UNSIGN) );
  NAND4_X1 U25 ( .A1(n20), .A2(n32), .A3(n26), .A4(n35), .ZN(MUX_SEL[0]) );
  AOI22_X1 U26 ( .A1(n29), .A2(n34), .B1(n24), .B2(n34), .ZN(n35) );
  AOI22_X1 U27 ( .A1(n22), .A2(n21), .B1(n49), .B2(n23), .ZN(n48) );
  INV_X1 U28 ( .A(n52), .ZN(n45) );
  OAI211_X1 U29 ( .C1(n42), .C2(n51), .A(n47), .B(n48), .ZN(CMP_OP[0]) );
  INV_X1 U30 ( .A(n29), .ZN(n51) );
  NOR2_X1 U31 ( .A1(n36), .A2(n15), .ZN(n30) );
  AND2_X1 U32 ( .A1(n23), .A2(n21), .ZN(ARITH_LOG) );
  NAND4_X1 U33 ( .A1(n20), .A2(n25), .A3(n26), .A4(n27), .ZN(MUX_SEL[2]) );
  NOR3_X1 U34 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n27) );
  INV_X1 U35 ( .A(CMP_OP[2]), .ZN(n25) );
  INV_X1 U36 ( .A(n31), .ZN(n28) );
  INV_X1 U37 ( .A(n18), .ZN(n49) );
  INV_X1 U38 ( .A(n16), .ZN(n33) );
  NOR3_X1 U39 ( .A1(n43), .A2(ALU_OP_CODE[4]), .A3(n36), .ZN(n21) );
  AOI222_X1 U56 ( .A1(n36), .A2(ALU_OP_CODE[3]), .B1(n22), .B2(ALU_OP_CODE[1]), 
        .C1(n43), .C2(ALU_OP_CODE[2]), .ZN(n19) );
  NOR2_X1 U57 ( .A1(ALU_OP_CODE[2]), .A2(ALU_OP_CODE[0]), .ZN(n34) );
  NOR3_X1 U58 ( .A1(n36), .A2(ALU_OP_CODE[3]), .A3(n37), .ZN(n24) );
  NOR3_X1 U59 ( .A1(ALU_OP_CODE[1]), .A2(ALU_OP_CODE[3]), .A3(n37), .ZN(n38)
         );
  INV_X1 U60 ( .A(EN_GUARD_CMP), .ZN(n52) );
  OAI21_X1 U61 ( .B1(ALU_OP_CODE[4]), .B2(n19), .A(n53), .ZN(EN_GUARD_CMP) );
  INV_X1 U62 ( .A(ALU_OP_CODE[1]), .ZN(n36) );
  AND2_X1 U63 ( .A1(ALU_OP_CODE[0]), .A2(n42), .ZN(n22) );
  OAI21_X1 U64 ( .B1(ALU_OP_CODE[4]), .B2(n19), .A(n20), .ZN(SUB_ADD) );
  INV_X1 U65 ( .A(ALU_OP_CODE[3]), .ZN(n43) );
  INV_X1 U66 ( .A(ALU_OP_CODE[4]), .ZN(n37) );
  INV_X1 U67 ( .A(ALU_OP_CODE[2]), .ZN(n42) );
  NOR2_X1 U68 ( .A1(n15), .A2(ALU_OP_CODE[1]), .ZN(n29) );
  NOR2_X1 U69 ( .A1(n42), .A2(ALU_OP_CODE[0]), .ZN(n23) );
  CLKBUF_X1 U70 ( .A(EN_GUARD_LOG), .Z(n41) );
  INV_X1 U71 ( .A(RST), .ZN(n53) );
endmodule


module MUX51_GEN_N32_0 ( A, B, C, D, E, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [2:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162;

  NAND2_X4 U1 ( .A1(n38), .A2(n2), .ZN(Y[2]) );
  NAND2_X2 U2 ( .A1(n34), .A2(n4), .ZN(Y[1]) );
  AOI22_X1 U3 ( .A1(C[1]), .A2(n21), .B1(A[1]), .B2(n18), .ZN(n34) );
  AND3_X2 U4 ( .A1(n45), .A2(n44), .A3(n43), .ZN(n1) );
  AND3_X2 U5 ( .A1(n41), .A2(n40), .A3(n39), .ZN(n2) );
  AND2_X2 U6 ( .A1(n32), .A2(n31), .ZN(n3) );
  AND3_X2 U7 ( .A1(n37), .A2(n36), .A3(n35), .ZN(n4) );
  AND2_X1 U8 ( .A1(C[2]), .A2(n21), .ZN(n5) );
  AND2_X2 U9 ( .A1(A[2]), .A2(n18), .ZN(n6) );
  NOR2_X2 U10 ( .A1(n5), .A2(n6), .ZN(n38) );
  NAND2_X2 U11 ( .A1(n26), .A2(n27), .ZN(n24) );
  BUF_X4 U12 ( .A(n155), .Z(n12) );
  CLKBUF_X1 U13 ( .A(n154), .Z(n8) );
  CLKBUF_X1 U14 ( .A(n154), .Z(n9) );
  NAND3_X4 U15 ( .A1(n30), .A2(n33), .A3(n3), .ZN(Y[0]) );
  AOI22_X2 U16 ( .A1(C[0]), .A2(n21), .B1(A[0]), .B2(n18), .ZN(n30) );
  NOR2_X4 U17 ( .A1(n25), .A2(n24), .ZN(n154) );
  AOI22_X2 U18 ( .A1(C[3]), .A2(n21), .B1(A[3]), .B2(n18), .ZN(n42) );
  BUF_X4 U19 ( .A(n158), .Z(n21) );
  NAND2_X4 U20 ( .A1(n42), .A2(n1), .ZN(Y[3]) );
  BUF_X4 U21 ( .A(n157), .Z(n18) );
  AND2_X2 U22 ( .A1(SEL[2]), .A2(SEL[1]), .ZN(n7) );
  CLKBUF_X1 U23 ( .A(n157), .Z(n17) );
  CLKBUF_X1 U24 ( .A(n157), .Z(n16) );
  CLKBUF_X1 U25 ( .A(n158), .Z(n20) );
  CLKBUF_X1 U26 ( .A(n158), .Z(n19) );
  BUF_X2 U27 ( .A(n156), .Z(n15) );
  BUF_X1 U28 ( .A(n155), .Z(n11) );
  BUF_X1 U29 ( .A(n155), .Z(n10) );
  BUF_X1 U30 ( .A(n156), .Z(n14) );
  BUF_X1 U31 ( .A(n156), .Z(n13) );
  NAND2_X1 U32 ( .A1(SEL[0]), .A2(n7), .ZN(n29) );
  INV_X1 U33 ( .A(SEL[1]), .ZN(n22) );
  NAND3_X1 U34 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n22), .ZN(n28) );
  NAND2_X1 U35 ( .A1(n29), .A2(n28), .ZN(n25) );
  INV_X1 U36 ( .A(SEL[0]), .ZN(n23) );
  NAND2_X1 U37 ( .A1(n23), .A2(n7), .ZN(n26) );
  NAND3_X1 U38 ( .A1(n23), .A2(SEL[2]), .A3(n22), .ZN(n27) );
  NAND2_X1 U39 ( .A1(E[0]), .A2(n154), .ZN(n33) );
  INV_X1 U40 ( .A(n26), .ZN(n155) );
  NAND2_X1 U41 ( .A1(B[0]), .A2(n12), .ZN(n32) );
  INV_X1 U42 ( .A(n27), .ZN(n156) );
  NAND2_X1 U43 ( .A1(D[0]), .A2(n15), .ZN(n31) );
  INV_X1 U44 ( .A(n28), .ZN(n158) );
  INV_X1 U45 ( .A(n29), .ZN(n157) );
  NAND2_X1 U46 ( .A1(E[1]), .A2(n154), .ZN(n37) );
  NAND2_X1 U47 ( .A1(B[1]), .A2(n12), .ZN(n36) );
  NAND2_X1 U48 ( .A1(D[1]), .A2(n15), .ZN(n35) );
  NAND2_X1 U49 ( .A1(E[2]), .A2(n154), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B[2]), .A2(n12), .ZN(n40) );
  NAND2_X1 U51 ( .A1(D[2]), .A2(n15), .ZN(n39) );
  NAND2_X1 U52 ( .A1(E[3]), .A2(n154), .ZN(n45) );
  NAND2_X1 U53 ( .A1(B[3]), .A2(n12), .ZN(n44) );
  NAND2_X1 U54 ( .A1(D[3]), .A2(n15), .ZN(n43) );
  NAND2_X1 U55 ( .A1(E[4]), .A2(n154), .ZN(n49) );
  NAND2_X1 U56 ( .A1(B[4]), .A2(n12), .ZN(n48) );
  NAND2_X1 U57 ( .A1(D[4]), .A2(n15), .ZN(n47) );
  AOI22_X1 U58 ( .A1(C[4]), .A2(n21), .B1(A[4]), .B2(n18), .ZN(n46) );
  NAND4_X1 U59 ( .A1(n49), .A2(n48), .A3(n47), .A4(n46), .ZN(Y[4]) );
  NAND2_X1 U60 ( .A1(E[5]), .A2(n154), .ZN(n53) );
  NAND2_X1 U61 ( .A1(B[5]), .A2(n12), .ZN(n52) );
  NAND2_X1 U62 ( .A1(D[5]), .A2(n15), .ZN(n51) );
  AOI22_X1 U63 ( .A1(C[5]), .A2(n21), .B1(A[5]), .B2(n18), .ZN(n50) );
  NAND4_X1 U64 ( .A1(n53), .A2(n52), .A3(n51), .A4(n50), .ZN(Y[5]) );
  NAND2_X1 U65 ( .A1(E[6]), .A2(n9), .ZN(n57) );
  NAND2_X1 U66 ( .A1(B[6]), .A2(n11), .ZN(n56) );
  NAND2_X1 U67 ( .A1(D[6]), .A2(n14), .ZN(n55) );
  AOI22_X1 U68 ( .A1(C[6]), .A2(n20), .B1(A[6]), .B2(n17), .ZN(n54) );
  NAND4_X1 U69 ( .A1(n57), .A2(n56), .A3(n55), .A4(n54), .ZN(Y[6]) );
  NAND2_X1 U70 ( .A1(E[7]), .A2(n9), .ZN(n61) );
  NAND2_X1 U71 ( .A1(B[7]), .A2(n11), .ZN(n60) );
  NAND2_X1 U72 ( .A1(D[7]), .A2(n14), .ZN(n59) );
  AOI22_X1 U73 ( .A1(C[7]), .A2(n20), .B1(A[7]), .B2(n17), .ZN(n58) );
  NAND4_X1 U74 ( .A1(n61), .A2(n60), .A3(n59), .A4(n58), .ZN(Y[7]) );
  NAND2_X1 U75 ( .A1(E[8]), .A2(n9), .ZN(n65) );
  NAND2_X1 U76 ( .A1(B[8]), .A2(n11), .ZN(n64) );
  NAND2_X1 U77 ( .A1(D[8]), .A2(n14), .ZN(n63) );
  AOI22_X1 U78 ( .A1(C[8]), .A2(n20), .B1(A[8]), .B2(n17), .ZN(n62) );
  NAND4_X1 U79 ( .A1(n65), .A2(n64), .A3(n63), .A4(n62), .ZN(Y[8]) );
  NAND2_X1 U80 ( .A1(E[9]), .A2(n9), .ZN(n69) );
  NAND2_X1 U81 ( .A1(B[9]), .A2(n11), .ZN(n68) );
  NAND2_X1 U82 ( .A1(D[9]), .A2(n14), .ZN(n67) );
  AOI22_X1 U83 ( .A1(C[9]), .A2(n20), .B1(A[9]), .B2(n17), .ZN(n66) );
  NAND4_X1 U84 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(Y[9]) );
  NAND2_X1 U85 ( .A1(E[10]), .A2(n9), .ZN(n73) );
  NAND2_X1 U86 ( .A1(B[10]), .A2(n11), .ZN(n72) );
  NAND2_X1 U87 ( .A1(D[10]), .A2(n14), .ZN(n71) );
  AOI22_X1 U88 ( .A1(C[10]), .A2(n20), .B1(A[10]), .B2(n17), .ZN(n70) );
  NAND4_X1 U89 ( .A1(n73), .A2(n72), .A3(n71), .A4(n70), .ZN(Y[10]) );
  NAND2_X1 U90 ( .A1(E[11]), .A2(n9), .ZN(n77) );
  NAND2_X1 U91 ( .A1(B[11]), .A2(n11), .ZN(n76) );
  NAND2_X1 U92 ( .A1(D[11]), .A2(n14), .ZN(n75) );
  AOI22_X1 U93 ( .A1(C[11]), .A2(n20), .B1(A[11]), .B2(n17), .ZN(n74) );
  NAND4_X1 U94 ( .A1(n77), .A2(n76), .A3(n75), .A4(n74), .ZN(Y[11]) );
  NAND2_X1 U95 ( .A1(E[12]), .A2(n9), .ZN(n81) );
  NAND2_X1 U96 ( .A1(B[12]), .A2(n11), .ZN(n80) );
  NAND2_X1 U97 ( .A1(D[12]), .A2(n14), .ZN(n79) );
  AOI22_X1 U98 ( .A1(C[12]), .A2(n20), .B1(A[12]), .B2(n17), .ZN(n78) );
  NAND4_X1 U99 ( .A1(n81), .A2(n80), .A3(n79), .A4(n78), .ZN(Y[12]) );
  NAND2_X1 U100 ( .A1(E[13]), .A2(n9), .ZN(n85) );
  NAND2_X1 U101 ( .A1(B[13]), .A2(n11), .ZN(n84) );
  NAND2_X1 U102 ( .A1(D[13]), .A2(n14), .ZN(n83) );
  AOI22_X1 U103 ( .A1(C[13]), .A2(n20), .B1(A[13]), .B2(n17), .ZN(n82) );
  NAND4_X1 U104 ( .A1(n85), .A2(n84), .A3(n83), .A4(n82), .ZN(Y[13]) );
  NAND2_X1 U105 ( .A1(E[14]), .A2(n9), .ZN(n89) );
  NAND2_X1 U106 ( .A1(B[14]), .A2(n11), .ZN(n88) );
  NAND2_X1 U107 ( .A1(D[14]), .A2(n14), .ZN(n87) );
  AOI22_X1 U108 ( .A1(C[14]), .A2(n20), .B1(A[14]), .B2(n17), .ZN(n86) );
  NAND4_X1 U109 ( .A1(n89), .A2(n88), .A3(n87), .A4(n86), .ZN(Y[14]) );
  NAND2_X1 U110 ( .A1(E[15]), .A2(n9), .ZN(n93) );
  NAND2_X1 U111 ( .A1(B[15]), .A2(n11), .ZN(n92) );
  NAND2_X1 U112 ( .A1(D[15]), .A2(n14), .ZN(n91) );
  AOI22_X1 U113 ( .A1(C[15]), .A2(n20), .B1(A[15]), .B2(n17), .ZN(n90) );
  NAND4_X1 U114 ( .A1(n93), .A2(n92), .A3(n91), .A4(n90), .ZN(Y[15]) );
  NAND2_X1 U115 ( .A1(E[16]), .A2(n9), .ZN(n97) );
  NAND2_X1 U116 ( .A1(B[16]), .A2(n11), .ZN(n96) );
  NAND2_X1 U117 ( .A1(D[16]), .A2(n14), .ZN(n95) );
  AOI22_X1 U118 ( .A1(C[16]), .A2(n20), .B1(A[16]), .B2(n17), .ZN(n94) );
  NAND4_X1 U119 ( .A1(n97), .A2(n96), .A3(n95), .A4(n94), .ZN(Y[16]) );
  NAND2_X1 U120 ( .A1(E[17]), .A2(n9), .ZN(n101) );
  NAND2_X1 U121 ( .A1(B[17]), .A2(n11), .ZN(n100) );
  NAND2_X1 U122 ( .A1(D[17]), .A2(n14), .ZN(n99) );
  AOI22_X1 U123 ( .A1(C[17]), .A2(n20), .B1(A[17]), .B2(n17), .ZN(n98) );
  NAND4_X1 U124 ( .A1(n101), .A2(n100), .A3(n99), .A4(n98), .ZN(Y[17]) );
  NAND2_X1 U125 ( .A1(E[18]), .A2(n9), .ZN(n105) );
  NAND2_X1 U126 ( .A1(B[18]), .A2(n11), .ZN(n104) );
  NAND2_X1 U127 ( .A1(D[18]), .A2(n14), .ZN(n103) );
  AOI22_X1 U128 ( .A1(C[18]), .A2(n20), .B1(A[18]), .B2(n17), .ZN(n102) );
  NAND4_X1 U129 ( .A1(n105), .A2(n104), .A3(n103), .A4(n102), .ZN(Y[18]) );
  NAND2_X1 U130 ( .A1(E[19]), .A2(n8), .ZN(n109) );
  NAND2_X1 U131 ( .A1(B[19]), .A2(n10), .ZN(n108) );
  NAND2_X1 U132 ( .A1(D[19]), .A2(n13), .ZN(n107) );
  AOI22_X1 U133 ( .A1(C[19]), .A2(n19), .B1(A[19]), .B2(n16), .ZN(n106) );
  NAND4_X1 U134 ( .A1(n109), .A2(n108), .A3(n107), .A4(n106), .ZN(Y[19]) );
  NAND2_X1 U135 ( .A1(E[20]), .A2(n8), .ZN(n113) );
  NAND2_X1 U136 ( .A1(B[20]), .A2(n10), .ZN(n112) );
  NAND2_X1 U137 ( .A1(D[20]), .A2(n13), .ZN(n111) );
  AOI22_X1 U138 ( .A1(C[20]), .A2(n19), .B1(A[20]), .B2(n16), .ZN(n110) );
  NAND4_X1 U139 ( .A1(n113), .A2(n112), .A3(n111), .A4(n110), .ZN(Y[20]) );
  NAND2_X1 U140 ( .A1(E[21]), .A2(n8), .ZN(n117) );
  NAND2_X1 U141 ( .A1(B[21]), .A2(n10), .ZN(n116) );
  NAND2_X1 U142 ( .A1(D[21]), .A2(n13), .ZN(n115) );
  AOI22_X1 U143 ( .A1(C[21]), .A2(n19), .B1(A[21]), .B2(n16), .ZN(n114) );
  NAND4_X1 U144 ( .A1(n117), .A2(n116), .A3(n115), .A4(n114), .ZN(Y[21]) );
  NAND2_X1 U145 ( .A1(E[22]), .A2(n8), .ZN(n121) );
  NAND2_X1 U146 ( .A1(B[22]), .A2(n10), .ZN(n120) );
  NAND2_X1 U147 ( .A1(D[22]), .A2(n13), .ZN(n119) );
  AOI22_X1 U148 ( .A1(C[22]), .A2(n19), .B1(A[22]), .B2(n16), .ZN(n118) );
  NAND4_X1 U149 ( .A1(n121), .A2(n120), .A3(n119), .A4(n118), .ZN(Y[22]) );
  NAND2_X1 U150 ( .A1(E[23]), .A2(n8), .ZN(n125) );
  NAND2_X1 U151 ( .A1(B[23]), .A2(n10), .ZN(n124) );
  NAND2_X1 U152 ( .A1(D[23]), .A2(n13), .ZN(n123) );
  AOI22_X1 U153 ( .A1(C[23]), .A2(n19), .B1(A[23]), .B2(n16), .ZN(n122) );
  NAND4_X1 U154 ( .A1(n125), .A2(n124), .A3(n123), .A4(n122), .ZN(Y[23]) );
  NAND2_X1 U155 ( .A1(E[24]), .A2(n8), .ZN(n129) );
  NAND2_X1 U156 ( .A1(B[24]), .A2(n10), .ZN(n128) );
  NAND2_X1 U157 ( .A1(D[24]), .A2(n13), .ZN(n127) );
  AOI22_X1 U158 ( .A1(C[24]), .A2(n19), .B1(A[24]), .B2(n16), .ZN(n126) );
  NAND4_X1 U159 ( .A1(n129), .A2(n128), .A3(n127), .A4(n126), .ZN(Y[24]) );
  NAND2_X1 U160 ( .A1(E[25]), .A2(n8), .ZN(n133) );
  NAND2_X1 U161 ( .A1(B[25]), .A2(n10), .ZN(n132) );
  NAND2_X1 U162 ( .A1(D[25]), .A2(n13), .ZN(n131) );
  AOI22_X1 U163 ( .A1(C[25]), .A2(n19), .B1(A[25]), .B2(n16), .ZN(n130) );
  NAND4_X1 U164 ( .A1(n133), .A2(n132), .A3(n131), .A4(n130), .ZN(Y[25]) );
  NAND2_X1 U165 ( .A1(E[26]), .A2(n8), .ZN(n137) );
  NAND2_X1 U166 ( .A1(B[26]), .A2(n10), .ZN(n136) );
  NAND2_X1 U167 ( .A1(D[26]), .A2(n13), .ZN(n135) );
  AOI22_X1 U168 ( .A1(C[26]), .A2(n19), .B1(A[26]), .B2(n16), .ZN(n134) );
  NAND4_X1 U169 ( .A1(n137), .A2(n136), .A3(n135), .A4(n134), .ZN(Y[26]) );
  NAND2_X1 U170 ( .A1(E[27]), .A2(n8), .ZN(n141) );
  NAND2_X1 U171 ( .A1(B[27]), .A2(n10), .ZN(n140) );
  NAND2_X1 U172 ( .A1(D[27]), .A2(n13), .ZN(n139) );
  AOI22_X1 U173 ( .A1(C[27]), .A2(n19), .B1(A[27]), .B2(n16), .ZN(n138) );
  NAND4_X1 U174 ( .A1(n141), .A2(n140), .A3(n139), .A4(n138), .ZN(Y[27]) );
  NAND2_X1 U175 ( .A1(E[28]), .A2(n8), .ZN(n145) );
  NAND2_X1 U176 ( .A1(B[28]), .A2(n10), .ZN(n144) );
  NAND2_X1 U177 ( .A1(D[28]), .A2(n13), .ZN(n143) );
  AOI22_X1 U178 ( .A1(C[28]), .A2(n19), .B1(A[28]), .B2(n16), .ZN(n142) );
  NAND4_X1 U179 ( .A1(n145), .A2(n144), .A3(n143), .A4(n142), .ZN(Y[28]) );
  NAND2_X1 U180 ( .A1(E[29]), .A2(n8), .ZN(n149) );
  NAND2_X1 U181 ( .A1(B[29]), .A2(n10), .ZN(n148) );
  NAND2_X1 U182 ( .A1(D[29]), .A2(n13), .ZN(n147) );
  AOI22_X1 U183 ( .A1(C[29]), .A2(n19), .B1(A[29]), .B2(n16), .ZN(n146) );
  NAND4_X1 U184 ( .A1(n149), .A2(n148), .A3(n147), .A4(n146), .ZN(Y[29]) );
  NAND2_X1 U185 ( .A1(E[30]), .A2(n8), .ZN(n153) );
  NAND2_X1 U186 ( .A1(B[30]), .A2(n10), .ZN(n152) );
  NAND2_X1 U187 ( .A1(D[30]), .A2(n13), .ZN(n151) );
  AOI22_X1 U188 ( .A1(C[30]), .A2(n19), .B1(A[30]), .B2(n16), .ZN(n150) );
  NAND4_X1 U189 ( .A1(n153), .A2(n152), .A3(n151), .A4(n150), .ZN(Y[30]) );
  NAND2_X1 U190 ( .A1(E[31]), .A2(n8), .ZN(n162) );
  NAND2_X1 U191 ( .A1(B[31]), .A2(n10), .ZN(n161) );
  NAND2_X1 U192 ( .A1(D[31]), .A2(n13), .ZN(n160) );
  AOI22_X1 U193 ( .A1(C[31]), .A2(n19), .B1(A[31]), .B2(n16), .ZN(n159) );
  NAND4_X1 U194 ( .A1(n162), .A2(n161), .A3(n160), .A4(n159), .ZN(Y[31]) );
endmodule


module BRANCH_N32 ( REG_A, BNEZ_SEL, CONFIRM_BRANCH, CONFIRM_JMP, BRANCH_SEL
 );
  input [31:0] REG_A;
  input BNEZ_SEL, CONFIRM_BRANCH, CONFIRM_JMP;
  output BRANCH_SEL;
  wire   OUT_COMP, OUT_INV, OUT_MUX, OUT_AND;

  EQU_COMPARATOR_N32_1 COMPARATOR_INST ( .A(REG_A), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .Y(OUT_COMP) );
  INV_1_123 INV_INST ( .A(OUT_COMP), .Y(OUT_INV) );
  MUX21_0 MUX_INST ( .A(OUT_INV), .B(OUT_COMP), .S(BNEZ_SEL), .Y(OUT_MUX) );
  AND_GATE_1_707 AND_INST ( .A(OUT_MUX), .B(CONFIRM_BRANCH), .Y(OUT_AND) );
  OR_GATE_0 OR_INST ( .A(OUT_AND), .B(CONFIRM_JMP), .Y(BRANCH_SEL) );
endmodule


module MUX41_GEN_N32_0 ( A, B, C, D, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] SEL;
  output [31:0] Y;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n1, n2,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  NAND2_X1 U70 ( .A1(n3), .A2(n4), .ZN(Y[9]) );
  NAND2_X1 U71 ( .A1(n9), .A2(n10), .ZN(Y[8]) );
  NAND2_X1 U72 ( .A1(n11), .A2(n12), .ZN(Y[7]) );
  NAND2_X1 U73 ( .A1(n13), .A2(n14), .ZN(Y[6]) );
  NAND2_X1 U74 ( .A1(n15), .A2(n16), .ZN(Y[5]) );
  NAND2_X1 U75 ( .A1(n17), .A2(n18), .ZN(Y[4]) );
  NAND2_X1 U76 ( .A1(n19), .A2(n20), .ZN(Y[3]) );
  NAND2_X1 U77 ( .A1(n21), .A2(n22), .ZN(Y[31]) );
  NAND2_X1 U78 ( .A1(n23), .A2(n24), .ZN(Y[30]) );
  NAND2_X1 U79 ( .A1(n25), .A2(n26), .ZN(Y[2]) );
  NAND2_X1 U80 ( .A1(n27), .A2(n28), .ZN(Y[29]) );
  NAND2_X1 U81 ( .A1(n29), .A2(n30), .ZN(Y[28]) );
  NAND2_X1 U82 ( .A1(n31), .A2(n32), .ZN(Y[27]) );
  NAND2_X1 U83 ( .A1(n33), .A2(n34), .ZN(Y[26]) );
  NAND2_X1 U84 ( .A1(n35), .A2(n36), .ZN(Y[25]) );
  NAND2_X1 U85 ( .A1(n37), .A2(n38), .ZN(Y[24]) );
  NAND2_X1 U86 ( .A1(n39), .A2(n40), .ZN(Y[23]) );
  NAND2_X1 U87 ( .A1(n41), .A2(n42), .ZN(Y[22]) );
  NAND2_X1 U88 ( .A1(n43), .A2(n44), .ZN(Y[21]) );
  NAND2_X1 U89 ( .A1(n45), .A2(n46), .ZN(Y[20]) );
  NAND2_X1 U90 ( .A1(n47), .A2(n48), .ZN(Y[1]) );
  NAND2_X1 U91 ( .A1(n49), .A2(n50), .ZN(Y[19]) );
  NAND2_X1 U92 ( .A1(n51), .A2(n52), .ZN(Y[18]) );
  NAND2_X1 U93 ( .A1(n53), .A2(n54), .ZN(Y[17]) );
  NAND2_X1 U94 ( .A1(n55), .A2(n56), .ZN(Y[16]) );
  NAND2_X1 U95 ( .A1(n57), .A2(n58), .ZN(Y[15]) );
  NAND2_X1 U96 ( .A1(n59), .A2(n60), .ZN(Y[14]) );
  NAND2_X1 U97 ( .A1(n61), .A2(n62), .ZN(Y[13]) );
  NAND2_X1 U98 ( .A1(n63), .A2(n64), .ZN(Y[12]) );
  NAND2_X1 U99 ( .A1(n65), .A2(n66), .ZN(Y[11]) );
  NAND2_X1 U100 ( .A1(n67), .A2(n68), .ZN(Y[10]) );
  NAND2_X1 U101 ( .A1(n69), .A2(n70), .ZN(Y[0]) );
  BUF_X1 U1 ( .A(n7), .Z(n74) );
  BUF_X1 U2 ( .A(n7), .Z(n73) );
  BUF_X1 U3 ( .A(n7), .Z(n75) );
  NOR3_X1 U4 ( .A1(n78), .A2(n72), .A3(n81), .ZN(n7) );
  BUF_X1 U5 ( .A(n6), .Z(n78) );
  BUF_X1 U6 ( .A(n5), .Z(n81) );
  BUF_X1 U7 ( .A(n6), .Z(n76) );
  BUF_X1 U8 ( .A(n6), .Z(n77) );
  BUF_X1 U9 ( .A(n5), .Z(n79) );
  BUF_X1 U10 ( .A(n5), .Z(n80) );
  NOR2_X1 U11 ( .A1(n71), .A2(SEL[1]), .ZN(n6) );
  BUF_X1 U12 ( .A(n8), .Z(n72) );
  AND2_X1 U13 ( .A1(SEL[1]), .A2(n71), .ZN(n5) );
  BUF_X1 U14 ( .A(n8), .Z(n1) );
  BUF_X1 U15 ( .A(n8), .Z(n2) );
  AND2_X1 U16 ( .A1(SEL[0]), .A2(SEL[1]), .ZN(n8) );
  INV_X1 U17 ( .A(SEL[0]), .ZN(n71) );
  AOI22_X1 U18 ( .A1(B[31]), .A2(n79), .B1(C[31]), .B2(n76), .ZN(n22) );
  AOI22_X1 U19 ( .A1(D[31]), .A2(n74), .B1(A[31]), .B2(n1), .ZN(n21) );
  AOI22_X1 U20 ( .A1(B[11]), .A2(n81), .B1(C[11]), .B2(n78), .ZN(n66) );
  AOI22_X1 U21 ( .A1(D[11]), .A2(n73), .B1(A[11]), .B2(n72), .ZN(n65) );
  AOI22_X1 U22 ( .A1(B[12]), .A2(n81), .B1(C[12]), .B2(n78), .ZN(n64) );
  AOI22_X1 U23 ( .A1(D[12]), .A2(n73), .B1(A[12]), .B2(n72), .ZN(n63) );
  AOI22_X1 U24 ( .A1(B[14]), .A2(n81), .B1(C[14]), .B2(n78), .ZN(n60) );
  AOI22_X1 U25 ( .A1(D[14]), .A2(n73), .B1(A[14]), .B2(n72), .ZN(n59) );
  AOI22_X1 U26 ( .A1(B[10]), .A2(n81), .B1(C[10]), .B2(n78), .ZN(n68) );
  AOI22_X1 U27 ( .A1(D[10]), .A2(n73), .B1(A[10]), .B2(n72), .ZN(n67) );
  AOI22_X1 U28 ( .A1(B[9]), .A2(n79), .B1(C[9]), .B2(n76), .ZN(n4) );
  AOI22_X1 U29 ( .A1(D[9]), .A2(n75), .B1(A[9]), .B2(n1), .ZN(n3) );
  AOI22_X1 U30 ( .A1(B[25]), .A2(n80), .B1(C[25]), .B2(n77), .ZN(n36) );
  AOI22_X1 U31 ( .A1(D[25]), .A2(n74), .B1(A[25]), .B2(n2), .ZN(n35) );
  AOI22_X1 U32 ( .A1(B[23]), .A2(n80), .B1(C[23]), .B2(n77), .ZN(n40) );
  AOI22_X1 U33 ( .A1(D[23]), .A2(n74), .B1(A[23]), .B2(n2), .ZN(n39) );
  AOI22_X1 U34 ( .A1(B[18]), .A2(n80), .B1(C[18]), .B2(n77), .ZN(n52) );
  AOI22_X1 U35 ( .A1(D[18]), .A2(n73), .B1(A[18]), .B2(n2), .ZN(n51) );
  AOI22_X1 U36 ( .A1(B[19]), .A2(n80), .B1(C[19]), .B2(n77), .ZN(n50) );
  AOI22_X1 U37 ( .A1(D[19]), .A2(n73), .B1(A[19]), .B2(n2), .ZN(n49) );
  AOI22_X1 U38 ( .A1(B[1]), .A2(n80), .B1(C[1]), .B2(n77), .ZN(n48) );
  AOI22_X1 U39 ( .A1(D[1]), .A2(n73), .B1(A[1]), .B2(n2), .ZN(n47) );
  AOI22_X1 U40 ( .A1(B[15]), .A2(n80), .B1(C[15]), .B2(n77), .ZN(n58) );
  AOI22_X1 U41 ( .A1(D[15]), .A2(n73), .B1(A[15]), .B2(n2), .ZN(n57) );
  AOI22_X1 U42 ( .A1(B[28]), .A2(n79), .B1(C[28]), .B2(n76), .ZN(n30) );
  AOI22_X1 U43 ( .A1(D[28]), .A2(n74), .B1(A[28]), .B2(n1), .ZN(n29) );
  AOI22_X1 U44 ( .A1(B[24]), .A2(n80), .B1(C[24]), .B2(n77), .ZN(n38) );
  AOI22_X1 U45 ( .A1(D[24]), .A2(n74), .B1(A[24]), .B2(n2), .ZN(n37) );
  AOI22_X1 U46 ( .A1(B[17]), .A2(n80), .B1(C[17]), .B2(n77), .ZN(n54) );
  AOI22_X1 U47 ( .A1(D[17]), .A2(n73), .B1(A[17]), .B2(n2), .ZN(n53) );
  AOI22_X1 U48 ( .A1(B[20]), .A2(n80), .B1(C[20]), .B2(n77), .ZN(n46) );
  AOI22_X1 U49 ( .A1(D[20]), .A2(n73), .B1(A[20]), .B2(n2), .ZN(n45) );
  AOI22_X1 U50 ( .A1(B[7]), .A2(n79), .B1(C[7]), .B2(n76), .ZN(n12) );
  AOI22_X1 U51 ( .A1(D[7]), .A2(n75), .B1(A[7]), .B2(n1), .ZN(n11) );
  AOI22_X1 U52 ( .A1(B[6]), .A2(n79), .B1(C[6]), .B2(n76), .ZN(n14) );
  AOI22_X1 U53 ( .A1(D[6]), .A2(n75), .B1(A[6]), .B2(n1), .ZN(n13) );
  AOI22_X1 U54 ( .A1(B[8]), .A2(n79), .B1(C[8]), .B2(n76), .ZN(n10) );
  AOI22_X1 U55 ( .A1(D[8]), .A2(n75), .B1(A[8]), .B2(n1), .ZN(n9) );
  AOI22_X1 U56 ( .A1(B[3]), .A2(n79), .B1(C[3]), .B2(n76), .ZN(n20) );
  AOI22_X1 U57 ( .A1(D[3]), .A2(n74), .B1(A[3]), .B2(n1), .ZN(n19) );
  AOI22_X1 U58 ( .A1(B[4]), .A2(n79), .B1(C[4]), .B2(n76), .ZN(n18) );
  AOI22_X1 U59 ( .A1(D[4]), .A2(n75), .B1(A[4]), .B2(n1), .ZN(n17) );
  AOI22_X1 U60 ( .A1(B[5]), .A2(n79), .B1(C[5]), .B2(n76), .ZN(n16) );
  AOI22_X1 U61 ( .A1(D[5]), .A2(n75), .B1(A[5]), .B2(n1), .ZN(n15) );
  AOI22_X1 U62 ( .A1(B[29]), .A2(n79), .B1(C[29]), .B2(n76), .ZN(n28) );
  AOI22_X1 U63 ( .A1(D[29]), .A2(n74), .B1(A[29]), .B2(n1), .ZN(n27) );
  AOI22_X1 U64 ( .A1(B[2]), .A2(n79), .B1(C[2]), .B2(n76), .ZN(n26) );
  AOI22_X1 U65 ( .A1(D[2]), .A2(n74), .B1(A[2]), .B2(n1), .ZN(n25) );
  AOI22_X1 U66 ( .A1(B[26]), .A2(n80), .B1(C[26]), .B2(n77), .ZN(n34) );
  AOI22_X1 U67 ( .A1(D[26]), .A2(n74), .B1(A[26]), .B2(n2), .ZN(n33) );
  AOI22_X1 U68 ( .A1(B[27]), .A2(n79), .B1(C[27]), .B2(n76), .ZN(n32) );
  AOI22_X1 U69 ( .A1(D[27]), .A2(n74), .B1(A[27]), .B2(n1), .ZN(n31) );
  AOI22_X1 U102 ( .A1(B[21]), .A2(n80), .B1(C[21]), .B2(n77), .ZN(n44) );
  AOI22_X1 U103 ( .A1(D[21]), .A2(n74), .B1(A[21]), .B2(n2), .ZN(n43) );
  AOI22_X1 U104 ( .A1(B[22]), .A2(n80), .B1(C[22]), .B2(n77), .ZN(n42) );
  AOI22_X1 U105 ( .A1(D[22]), .A2(n74), .B1(A[22]), .B2(n2), .ZN(n41) );
  AOI22_X1 U106 ( .A1(B[16]), .A2(n80), .B1(C[16]), .B2(n77), .ZN(n56) );
  AOI22_X1 U107 ( .A1(D[16]), .A2(n73), .B1(A[16]), .B2(n2), .ZN(n55) );
  AOI22_X1 U108 ( .A1(B[13]), .A2(n81), .B1(C[13]), .B2(n78), .ZN(n62) );
  AOI22_X1 U109 ( .A1(D[13]), .A2(n73), .B1(A[13]), .B2(n72), .ZN(n61) );
  AOI22_X1 U110 ( .A1(B[0]), .A2(n81), .B1(C[0]), .B2(n78), .ZN(n70) );
  AOI22_X1 U111 ( .A1(D[0]), .A2(n73), .B1(A[0]), .B2(n72), .ZN(n69) );
  AOI22_X1 U112 ( .A1(B[30]), .A2(n79), .B1(C[30]), .B2(n76), .ZN(n24) );
  AOI22_X1 U113 ( .A1(D[30]), .A2(n74), .B1(A[30]), .B2(n1), .ZN(n23) );
endmodule


module CSA_N4_0 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_RCA_1;
  wire   [3:0] S_RCA_2;

  RCA_GEN_N4_0 RCA_1 ( .A(A), .B(B), .Ci(1'b0), .S(S_RCA_1) );
  RCA_GEN_N4_31 RCA_2 ( .A(A), .B(B), .Ci(1'b1), .S(S_RCA_2) );
  MUX21_GEN_N4_0 MUX_SUM ( .A(S_RCA_2), .B(S_RCA_1), .SEL(Ci), .Y(S) );
endmodule


module MUX31_GEN_N5 ( A, B, C, SEL, Y );
  input [4:0] A;
  input [4:0] B;
  input [4:0] C;
  input [1:0] SEL;
  output [4:0] Y;
  wire   n8, n9, n10, n11, n12, n13, n14, n15, n16;

  NOR2_X1 U1 ( .A1(n10), .A2(n9), .ZN(n11) );
  NOR2_X1 U2 ( .A1(n16), .A2(SEL[0]), .ZN(n10) );
  INV_X1 U3 ( .A(SEL[1]), .ZN(n16) );
  AND2_X1 U4 ( .A1(SEL[0]), .A2(SEL[1]), .ZN(n9) );
  INV_X1 U5 ( .A(n13), .ZN(Y[2]) );
  AOI222_X1 U6 ( .A1(A[2]), .A2(n9), .B1(B[2]), .B2(n10), .C1(C[2]), .C2(n11), 
        .ZN(n13) );
  INV_X1 U7 ( .A(n12), .ZN(Y[3]) );
  AOI222_X1 U8 ( .A1(A[3]), .A2(n9), .B1(B[3]), .B2(n10), .C1(C[3]), .C2(n11), 
        .ZN(n12) );
  INV_X1 U9 ( .A(n15), .ZN(Y[0]) );
  AOI222_X1 U10 ( .A1(A[0]), .A2(n9), .B1(B[0]), .B2(n10), .C1(C[0]), .C2(n11), 
        .ZN(n15) );
  INV_X1 U11 ( .A(n14), .ZN(Y[1]) );
  AOI222_X1 U12 ( .A1(A[1]), .A2(n9), .B1(B[1]), .B2(n10), .C1(C[1]), .C2(n11), 
        .ZN(n14) );
  INV_X1 U13 ( .A(n8), .ZN(Y[4]) );
  AOI222_X1 U14 ( .A1(A[4]), .A2(n9), .B1(B[4]), .B2(n10), .C1(C[4]), .C2(n11), 
        .ZN(n8) );
endmodule


module REG_FILE_N32_N_ADDR5 ( CLK, RST, EN, RD1, RD2, WR, ADDR_WR, ADDR_RD1, 
        ADDR_RD2, DATA_IN, DATA_OUT_1, DATA_OUT_2 );
  input [4:0] ADDR_WR;
  input [4:0] ADDR_RD1;
  input [4:0] ADDR_RD2;
  input [31:0] DATA_IN;
  output [31:0] DATA_OUT_1;
  output [31:0] DATA_OUT_2;
  input CLK, RST, EN, RD1, RD2, WR;
  wire   \REGISTERS[31][31] , \REGISTERS[31][30] , \REGISTERS[31][29] ,
         \REGISTERS[31][28] , \REGISTERS[31][27] , \REGISTERS[31][26] ,
         \REGISTERS[31][25] , \REGISTERS[31][24] , \REGISTERS[31][23] ,
         \REGISTERS[31][22] , \REGISTERS[31][21] , \REGISTERS[31][20] ,
         \REGISTERS[31][19] , \REGISTERS[31][18] , \REGISTERS[31][17] ,
         \REGISTERS[31][16] , \REGISTERS[31][15] , \REGISTERS[31][14] ,
         \REGISTERS[31][13] , \REGISTERS[31][12] , \REGISTERS[31][11] ,
         \REGISTERS[31][10] , \REGISTERS[31][9] , \REGISTERS[31][8] ,
         \REGISTERS[31][7] , \REGISTERS[31][6] , \REGISTERS[31][5] ,
         \REGISTERS[31][4] , \REGISTERS[31][3] , \REGISTERS[31][2] ,
         \REGISTERS[31][1] , \REGISTERS[31][0] , \REGISTERS[30][31] ,
         \REGISTERS[30][30] , \REGISTERS[30][29] , \REGISTERS[30][28] ,
         \REGISTERS[30][27] , \REGISTERS[30][26] , \REGISTERS[30][25] ,
         \REGISTERS[30][24] , \REGISTERS[30][23] , \REGISTERS[30][22] ,
         \REGISTERS[30][21] , \REGISTERS[30][20] , \REGISTERS[30][19] ,
         \REGISTERS[30][18] , \REGISTERS[30][17] , \REGISTERS[30][16] ,
         \REGISTERS[30][15] , \REGISTERS[30][14] , \REGISTERS[30][13] ,
         \REGISTERS[30][12] , \REGISTERS[30][11] , \REGISTERS[30][10] ,
         \REGISTERS[30][9] , \REGISTERS[30][8] , \REGISTERS[30][7] ,
         \REGISTERS[30][6] , \REGISTERS[30][5] , \REGISTERS[30][4] ,
         \REGISTERS[30][3] , \REGISTERS[30][2] , \REGISTERS[30][1] ,
         \REGISTERS[30][0] , \REGISTERS[29][31] , \REGISTERS[29][30] ,
         \REGISTERS[29][29] , \REGISTERS[29][28] , \REGISTERS[29][27] ,
         \REGISTERS[29][26] , \REGISTERS[29][25] , \REGISTERS[29][24] ,
         \REGISTERS[29][23] , \REGISTERS[29][22] , \REGISTERS[29][21] ,
         \REGISTERS[29][20] , \REGISTERS[29][19] , \REGISTERS[29][18] ,
         \REGISTERS[29][17] , \REGISTERS[29][16] , \REGISTERS[29][15] ,
         \REGISTERS[29][14] , \REGISTERS[29][13] , \REGISTERS[29][12] ,
         \REGISTERS[29][11] , \REGISTERS[29][10] , \REGISTERS[29][9] ,
         \REGISTERS[29][8] , \REGISTERS[29][7] , \REGISTERS[29][6] ,
         \REGISTERS[29][5] , \REGISTERS[29][4] , \REGISTERS[29][3] ,
         \REGISTERS[29][2] , \REGISTERS[29][1] , \REGISTERS[29][0] ,
         \REGISTERS[28][31] , \REGISTERS[28][30] , \REGISTERS[28][29] ,
         \REGISTERS[28][28] , \REGISTERS[28][27] , \REGISTERS[28][26] ,
         \REGISTERS[28][25] , \REGISTERS[28][24] , \REGISTERS[28][23] ,
         \REGISTERS[28][22] , \REGISTERS[28][21] , \REGISTERS[28][20] ,
         \REGISTERS[28][19] , \REGISTERS[28][18] , \REGISTERS[28][17] ,
         \REGISTERS[28][16] , \REGISTERS[28][15] , \REGISTERS[28][14] ,
         \REGISTERS[28][13] , \REGISTERS[28][12] , \REGISTERS[28][11] ,
         \REGISTERS[28][10] , \REGISTERS[28][9] , \REGISTERS[28][8] ,
         \REGISTERS[28][7] , \REGISTERS[28][6] , \REGISTERS[28][5] ,
         \REGISTERS[28][4] , \REGISTERS[28][3] , \REGISTERS[28][2] ,
         \REGISTERS[28][1] , \REGISTERS[28][0] , \REGISTERS[27][31] ,
         \REGISTERS[27][30] , \REGISTERS[27][29] , \REGISTERS[27][28] ,
         \REGISTERS[27][27] , \REGISTERS[27][26] , \REGISTERS[27][25] ,
         \REGISTERS[27][24] , \REGISTERS[27][23] , \REGISTERS[27][22] ,
         \REGISTERS[27][21] , \REGISTERS[27][20] , \REGISTERS[27][19] ,
         \REGISTERS[27][18] , \REGISTERS[27][17] , \REGISTERS[27][16] ,
         \REGISTERS[27][15] , \REGISTERS[27][14] , \REGISTERS[27][13] ,
         \REGISTERS[27][12] , \REGISTERS[27][11] , \REGISTERS[27][10] ,
         \REGISTERS[27][9] , \REGISTERS[27][8] , \REGISTERS[27][7] ,
         \REGISTERS[27][6] , \REGISTERS[27][5] , \REGISTERS[27][4] ,
         \REGISTERS[27][3] , \REGISTERS[27][2] , \REGISTERS[27][1] ,
         \REGISTERS[27][0] , \REGISTERS[26][31] , \REGISTERS[26][30] ,
         \REGISTERS[26][29] , \REGISTERS[26][28] , \REGISTERS[26][27] ,
         \REGISTERS[26][26] , \REGISTERS[26][25] , \REGISTERS[26][24] ,
         \REGISTERS[26][23] , \REGISTERS[26][22] , \REGISTERS[26][21] ,
         \REGISTERS[26][20] , \REGISTERS[26][19] , \REGISTERS[26][18] ,
         \REGISTERS[26][17] , \REGISTERS[26][16] , \REGISTERS[26][15] ,
         \REGISTERS[26][14] , \REGISTERS[26][13] , \REGISTERS[26][12] ,
         \REGISTERS[26][11] , \REGISTERS[26][10] , \REGISTERS[26][9] ,
         \REGISTERS[26][8] , \REGISTERS[26][7] , \REGISTERS[26][6] ,
         \REGISTERS[26][5] , \REGISTERS[26][4] , \REGISTERS[26][3] ,
         \REGISTERS[26][2] , \REGISTERS[26][1] , \REGISTERS[26][0] ,
         \REGISTERS[25][31] , \REGISTERS[25][30] , \REGISTERS[25][29] ,
         \REGISTERS[25][28] , \REGISTERS[25][27] , \REGISTERS[25][26] ,
         \REGISTERS[25][25] , \REGISTERS[25][24] , \REGISTERS[25][23] ,
         \REGISTERS[25][22] , \REGISTERS[25][21] , \REGISTERS[25][20] ,
         \REGISTERS[25][19] , \REGISTERS[25][18] , \REGISTERS[25][17] ,
         \REGISTERS[25][16] , \REGISTERS[25][15] , \REGISTERS[25][14] ,
         \REGISTERS[25][13] , \REGISTERS[25][12] , \REGISTERS[25][11] ,
         \REGISTERS[25][10] , \REGISTERS[25][9] , \REGISTERS[25][8] ,
         \REGISTERS[25][7] , \REGISTERS[25][6] , \REGISTERS[25][5] ,
         \REGISTERS[25][4] , \REGISTERS[25][3] , \REGISTERS[25][2] ,
         \REGISTERS[25][1] , \REGISTERS[25][0] , \REGISTERS[24][31] ,
         \REGISTERS[24][30] , \REGISTERS[24][29] , \REGISTERS[24][28] ,
         \REGISTERS[24][27] , \REGISTERS[24][26] , \REGISTERS[24][25] ,
         \REGISTERS[24][24] , \REGISTERS[24][23] , \REGISTERS[24][22] ,
         \REGISTERS[24][21] , \REGISTERS[24][20] , \REGISTERS[24][19] ,
         \REGISTERS[24][18] , \REGISTERS[24][17] , \REGISTERS[24][16] ,
         \REGISTERS[24][15] , \REGISTERS[24][14] , \REGISTERS[24][13] ,
         \REGISTERS[24][12] , \REGISTERS[24][11] , \REGISTERS[24][10] ,
         \REGISTERS[24][9] , \REGISTERS[24][8] , \REGISTERS[24][7] ,
         \REGISTERS[24][6] , \REGISTERS[24][5] , \REGISTERS[24][4] ,
         \REGISTERS[24][3] , \REGISTERS[24][2] , \REGISTERS[24][1] ,
         \REGISTERS[24][0] , \REGISTERS[23][31] , \REGISTERS[23][30] ,
         \REGISTERS[23][29] , \REGISTERS[23][28] , \REGISTERS[23][27] ,
         \REGISTERS[23][26] , \REGISTERS[23][25] , \REGISTERS[23][24] ,
         \REGISTERS[23][23] , \REGISTERS[23][22] , \REGISTERS[23][21] ,
         \REGISTERS[23][20] , \REGISTERS[23][19] , \REGISTERS[23][18] ,
         \REGISTERS[23][17] , \REGISTERS[23][16] , \REGISTERS[23][15] ,
         \REGISTERS[23][14] , \REGISTERS[23][13] , \REGISTERS[23][12] ,
         \REGISTERS[23][11] , \REGISTERS[23][10] , \REGISTERS[23][9] ,
         \REGISTERS[23][8] , \REGISTERS[23][7] , \REGISTERS[23][6] ,
         \REGISTERS[23][5] , \REGISTERS[23][4] , \REGISTERS[23][3] ,
         \REGISTERS[23][2] , \REGISTERS[23][1] , \REGISTERS[23][0] ,
         \REGISTERS[22][31] , \REGISTERS[22][30] , \REGISTERS[22][29] ,
         \REGISTERS[22][28] , \REGISTERS[22][27] , \REGISTERS[22][26] ,
         \REGISTERS[22][25] , \REGISTERS[22][24] , \REGISTERS[22][23] ,
         \REGISTERS[22][22] , \REGISTERS[22][21] , \REGISTERS[22][20] ,
         \REGISTERS[22][19] , \REGISTERS[22][18] , \REGISTERS[22][17] ,
         \REGISTERS[22][16] , \REGISTERS[22][15] , \REGISTERS[22][14] ,
         \REGISTERS[22][13] , \REGISTERS[22][12] , \REGISTERS[22][11] ,
         \REGISTERS[22][10] , \REGISTERS[22][9] , \REGISTERS[22][8] ,
         \REGISTERS[22][7] , \REGISTERS[22][6] , \REGISTERS[22][5] ,
         \REGISTERS[22][4] , \REGISTERS[22][3] , \REGISTERS[22][2] ,
         \REGISTERS[22][1] , \REGISTERS[22][0] , \REGISTERS[21][31] ,
         \REGISTERS[21][30] , \REGISTERS[21][29] , \REGISTERS[21][28] ,
         \REGISTERS[21][27] , \REGISTERS[21][26] , \REGISTERS[21][25] ,
         \REGISTERS[21][24] , \REGISTERS[21][23] , \REGISTERS[21][22] ,
         \REGISTERS[21][21] , \REGISTERS[21][20] , \REGISTERS[21][19] ,
         \REGISTERS[21][18] , \REGISTERS[21][17] , \REGISTERS[21][16] ,
         \REGISTERS[21][15] , \REGISTERS[21][14] , \REGISTERS[21][13] ,
         \REGISTERS[21][12] , \REGISTERS[21][11] , \REGISTERS[21][10] ,
         \REGISTERS[21][9] , \REGISTERS[21][8] , \REGISTERS[21][7] ,
         \REGISTERS[21][6] , \REGISTERS[21][5] , \REGISTERS[21][4] ,
         \REGISTERS[21][3] , \REGISTERS[21][2] , \REGISTERS[21][1] ,
         \REGISTERS[21][0] , \REGISTERS[20][31] , \REGISTERS[20][30] ,
         \REGISTERS[20][29] , \REGISTERS[20][28] , \REGISTERS[20][27] ,
         \REGISTERS[20][26] , \REGISTERS[20][25] , \REGISTERS[20][24] ,
         \REGISTERS[20][23] , \REGISTERS[20][22] , \REGISTERS[20][21] ,
         \REGISTERS[20][20] , \REGISTERS[20][19] , \REGISTERS[20][18] ,
         \REGISTERS[20][17] , \REGISTERS[20][16] , \REGISTERS[20][15] ,
         \REGISTERS[20][14] , \REGISTERS[20][13] , \REGISTERS[20][12] ,
         \REGISTERS[20][11] , \REGISTERS[20][10] , \REGISTERS[20][9] ,
         \REGISTERS[20][8] , \REGISTERS[20][7] , \REGISTERS[20][6] ,
         \REGISTERS[20][5] , \REGISTERS[20][4] , \REGISTERS[20][3] ,
         \REGISTERS[20][2] , \REGISTERS[20][1] , \REGISTERS[20][0] ,
         \REGISTERS[19][31] , \REGISTERS[19][30] , \REGISTERS[19][29] ,
         \REGISTERS[19][28] , \REGISTERS[19][27] , \REGISTERS[19][26] ,
         \REGISTERS[19][25] , \REGISTERS[19][24] , \REGISTERS[19][23] ,
         \REGISTERS[19][22] , \REGISTERS[19][21] , \REGISTERS[19][20] ,
         \REGISTERS[19][19] , \REGISTERS[19][18] , \REGISTERS[19][17] ,
         \REGISTERS[19][16] , \REGISTERS[19][15] , \REGISTERS[19][14] ,
         \REGISTERS[19][13] , \REGISTERS[19][12] , \REGISTERS[19][11] ,
         \REGISTERS[19][10] , \REGISTERS[19][9] , \REGISTERS[19][8] ,
         \REGISTERS[19][7] , \REGISTERS[19][6] , \REGISTERS[19][5] ,
         \REGISTERS[19][4] , \REGISTERS[19][3] , \REGISTERS[19][2] ,
         \REGISTERS[19][1] , \REGISTERS[19][0] , \REGISTERS[18][31] ,
         \REGISTERS[18][30] , \REGISTERS[18][29] , \REGISTERS[18][28] ,
         \REGISTERS[18][27] , \REGISTERS[18][26] , \REGISTERS[18][25] ,
         \REGISTERS[18][24] , \REGISTERS[18][23] , \REGISTERS[18][22] ,
         \REGISTERS[18][21] , \REGISTERS[18][20] , \REGISTERS[18][19] ,
         \REGISTERS[18][18] , \REGISTERS[18][17] , \REGISTERS[18][16] ,
         \REGISTERS[18][15] , \REGISTERS[18][14] , \REGISTERS[18][13] ,
         \REGISTERS[18][12] , \REGISTERS[18][11] , \REGISTERS[18][10] ,
         \REGISTERS[18][9] , \REGISTERS[18][8] , \REGISTERS[18][7] ,
         \REGISTERS[18][6] , \REGISTERS[18][5] , \REGISTERS[18][4] ,
         \REGISTERS[18][3] , \REGISTERS[18][2] , \REGISTERS[18][1] ,
         \REGISTERS[18][0] , \REGISTERS[17][31] , \REGISTERS[17][30] ,
         \REGISTERS[17][29] , \REGISTERS[17][28] , \REGISTERS[17][27] ,
         \REGISTERS[17][26] , \REGISTERS[17][25] , \REGISTERS[17][24] ,
         \REGISTERS[17][23] , \REGISTERS[17][22] , \REGISTERS[17][21] ,
         \REGISTERS[17][20] , \REGISTERS[17][19] , \REGISTERS[17][18] ,
         \REGISTERS[17][17] , \REGISTERS[17][16] , \REGISTERS[17][15] ,
         \REGISTERS[17][14] , \REGISTERS[17][13] , \REGISTERS[17][12] ,
         \REGISTERS[17][11] , \REGISTERS[17][10] , \REGISTERS[17][9] ,
         \REGISTERS[17][8] , \REGISTERS[17][7] , \REGISTERS[17][6] ,
         \REGISTERS[17][5] , \REGISTERS[17][4] , \REGISTERS[17][3] ,
         \REGISTERS[17][2] , \REGISTERS[17][1] , \REGISTERS[17][0] ,
         \REGISTERS[16][31] , \REGISTERS[16][30] , \REGISTERS[16][29] ,
         \REGISTERS[16][28] , \REGISTERS[16][27] , \REGISTERS[16][26] ,
         \REGISTERS[16][25] , \REGISTERS[16][24] , \REGISTERS[16][23] ,
         \REGISTERS[16][22] , \REGISTERS[16][21] , \REGISTERS[16][20] ,
         \REGISTERS[16][19] , \REGISTERS[16][18] , \REGISTERS[16][17] ,
         \REGISTERS[16][16] , \REGISTERS[16][15] , \REGISTERS[16][14] ,
         \REGISTERS[16][13] , \REGISTERS[16][12] , \REGISTERS[16][11] ,
         \REGISTERS[16][10] , \REGISTERS[16][9] , \REGISTERS[16][8] ,
         \REGISTERS[16][7] , \REGISTERS[16][6] , \REGISTERS[16][5] ,
         \REGISTERS[16][4] , \REGISTERS[16][3] , \REGISTERS[16][2] ,
         \REGISTERS[16][1] , \REGISTERS[16][0] , \REGISTERS[15][31] ,
         \REGISTERS[15][30] , \REGISTERS[15][29] , \REGISTERS[15][28] ,
         \REGISTERS[15][27] , \REGISTERS[15][26] , \REGISTERS[15][25] ,
         \REGISTERS[15][24] , \REGISTERS[15][23] , \REGISTERS[15][22] ,
         \REGISTERS[15][21] , \REGISTERS[15][20] , \REGISTERS[15][19] ,
         \REGISTERS[15][18] , \REGISTERS[15][17] , \REGISTERS[15][16] ,
         \REGISTERS[15][15] , \REGISTERS[15][14] , \REGISTERS[15][13] ,
         \REGISTERS[15][12] , \REGISTERS[15][11] , \REGISTERS[15][10] ,
         \REGISTERS[15][9] , \REGISTERS[15][8] , \REGISTERS[15][7] ,
         \REGISTERS[15][6] , \REGISTERS[15][5] , \REGISTERS[15][4] ,
         \REGISTERS[15][3] , \REGISTERS[15][2] , \REGISTERS[15][1] ,
         \REGISTERS[15][0] , \REGISTERS[14][31] , \REGISTERS[14][30] ,
         \REGISTERS[14][29] , \REGISTERS[14][28] , \REGISTERS[14][27] ,
         \REGISTERS[14][26] , \REGISTERS[14][25] , \REGISTERS[14][24] ,
         \REGISTERS[14][23] , \REGISTERS[14][22] , \REGISTERS[14][21] ,
         \REGISTERS[14][20] , \REGISTERS[14][19] , \REGISTERS[14][18] ,
         \REGISTERS[14][17] , \REGISTERS[14][16] , \REGISTERS[14][15] ,
         \REGISTERS[14][14] , \REGISTERS[14][13] , \REGISTERS[14][12] ,
         \REGISTERS[14][11] , \REGISTERS[14][10] , \REGISTERS[14][9] ,
         \REGISTERS[14][8] , \REGISTERS[14][7] , \REGISTERS[14][6] ,
         \REGISTERS[14][5] , \REGISTERS[14][4] , \REGISTERS[14][3] ,
         \REGISTERS[14][2] , \REGISTERS[14][1] , \REGISTERS[14][0] ,
         \REGISTERS[13][31] , \REGISTERS[13][30] , \REGISTERS[13][29] ,
         \REGISTERS[13][28] , \REGISTERS[13][27] , \REGISTERS[13][26] ,
         \REGISTERS[13][25] , \REGISTERS[13][24] , \REGISTERS[13][23] ,
         \REGISTERS[13][22] , \REGISTERS[13][21] , \REGISTERS[13][20] ,
         \REGISTERS[13][19] , \REGISTERS[13][18] , \REGISTERS[13][17] ,
         \REGISTERS[13][16] , \REGISTERS[13][15] , \REGISTERS[13][14] ,
         \REGISTERS[13][13] , \REGISTERS[13][12] , \REGISTERS[13][11] ,
         \REGISTERS[13][10] , \REGISTERS[13][9] , \REGISTERS[13][8] ,
         \REGISTERS[13][7] , \REGISTERS[13][6] , \REGISTERS[13][5] ,
         \REGISTERS[13][4] , \REGISTERS[13][3] , \REGISTERS[13][2] ,
         \REGISTERS[13][1] , \REGISTERS[13][0] , \REGISTERS[12][31] ,
         \REGISTERS[12][30] , \REGISTERS[12][29] , \REGISTERS[12][28] ,
         \REGISTERS[12][27] , \REGISTERS[12][26] , \REGISTERS[12][25] ,
         \REGISTERS[12][24] , \REGISTERS[12][23] , \REGISTERS[12][22] ,
         \REGISTERS[12][21] , \REGISTERS[12][20] , \REGISTERS[12][19] ,
         \REGISTERS[12][18] , \REGISTERS[12][17] , \REGISTERS[12][16] ,
         \REGISTERS[12][15] , \REGISTERS[12][14] , \REGISTERS[12][13] ,
         \REGISTERS[12][12] , \REGISTERS[12][11] , \REGISTERS[12][10] ,
         \REGISTERS[12][9] , \REGISTERS[12][8] , \REGISTERS[12][7] ,
         \REGISTERS[12][6] , \REGISTERS[12][5] , \REGISTERS[12][4] ,
         \REGISTERS[12][3] , \REGISTERS[12][2] , \REGISTERS[12][1] ,
         \REGISTERS[12][0] , \REGISTERS[11][31] , \REGISTERS[11][30] ,
         \REGISTERS[11][29] , \REGISTERS[11][28] , \REGISTERS[11][27] ,
         \REGISTERS[11][26] , \REGISTERS[11][25] , \REGISTERS[11][24] ,
         \REGISTERS[11][23] , \REGISTERS[11][22] , \REGISTERS[11][21] ,
         \REGISTERS[11][20] , \REGISTERS[11][19] , \REGISTERS[11][18] ,
         \REGISTERS[11][17] , \REGISTERS[11][16] , \REGISTERS[11][15] ,
         \REGISTERS[11][14] , \REGISTERS[11][13] , \REGISTERS[11][12] ,
         \REGISTERS[11][11] , \REGISTERS[11][10] , \REGISTERS[11][9] ,
         \REGISTERS[11][8] , \REGISTERS[11][7] , \REGISTERS[11][6] ,
         \REGISTERS[11][5] , \REGISTERS[11][4] , \REGISTERS[11][3] ,
         \REGISTERS[11][2] , \REGISTERS[11][1] , \REGISTERS[11][0] ,
         \REGISTERS[10][31] , \REGISTERS[10][30] , \REGISTERS[10][29] ,
         \REGISTERS[10][28] , \REGISTERS[10][27] , \REGISTERS[10][26] ,
         \REGISTERS[10][25] , \REGISTERS[10][24] , \REGISTERS[10][23] ,
         \REGISTERS[10][22] , \REGISTERS[10][21] , \REGISTERS[10][20] ,
         \REGISTERS[10][19] , \REGISTERS[10][18] , \REGISTERS[10][17] ,
         \REGISTERS[10][16] , \REGISTERS[10][15] , \REGISTERS[10][14] ,
         \REGISTERS[10][13] , \REGISTERS[10][12] , \REGISTERS[10][11] ,
         \REGISTERS[10][10] , \REGISTERS[10][9] , \REGISTERS[10][8] ,
         \REGISTERS[10][7] , \REGISTERS[10][6] , \REGISTERS[10][5] ,
         \REGISTERS[10][4] , \REGISTERS[10][3] , \REGISTERS[10][2] ,
         \REGISTERS[10][1] , \REGISTERS[10][0] , \REGISTERS[9][31] ,
         \REGISTERS[9][30] , \REGISTERS[9][29] , \REGISTERS[9][28] ,
         \REGISTERS[9][27] , \REGISTERS[9][26] , \REGISTERS[9][25] ,
         \REGISTERS[9][24] , \REGISTERS[9][23] , \REGISTERS[9][22] ,
         \REGISTERS[9][21] , \REGISTERS[9][20] , \REGISTERS[9][19] ,
         \REGISTERS[9][18] , \REGISTERS[9][17] , \REGISTERS[9][16] ,
         \REGISTERS[9][15] , \REGISTERS[9][14] , \REGISTERS[9][13] ,
         \REGISTERS[9][12] , \REGISTERS[9][11] , \REGISTERS[9][10] ,
         \REGISTERS[9][9] , \REGISTERS[9][8] , \REGISTERS[9][7] ,
         \REGISTERS[9][6] , \REGISTERS[9][5] , \REGISTERS[9][4] ,
         \REGISTERS[9][3] , \REGISTERS[9][2] , \REGISTERS[9][1] ,
         \REGISTERS[9][0] , \REGISTERS[8][31] , \REGISTERS[8][30] ,
         \REGISTERS[8][29] , \REGISTERS[8][28] , \REGISTERS[8][27] ,
         \REGISTERS[8][26] , \REGISTERS[8][25] , \REGISTERS[8][24] ,
         \REGISTERS[8][23] , \REGISTERS[8][22] , \REGISTERS[8][21] ,
         \REGISTERS[8][20] , \REGISTERS[8][19] , \REGISTERS[8][18] ,
         \REGISTERS[8][17] , \REGISTERS[8][16] , \REGISTERS[8][15] ,
         \REGISTERS[8][14] , \REGISTERS[8][13] , \REGISTERS[8][12] ,
         \REGISTERS[8][11] , \REGISTERS[8][10] , \REGISTERS[8][9] ,
         \REGISTERS[8][8] , \REGISTERS[8][7] , \REGISTERS[8][6] ,
         \REGISTERS[8][5] , \REGISTERS[8][4] , \REGISTERS[8][3] ,
         \REGISTERS[8][2] , \REGISTERS[8][1] , \REGISTERS[8][0] ,
         \REGISTERS[7][31] , \REGISTERS[7][30] , \REGISTERS[7][29] ,
         \REGISTERS[7][28] , \REGISTERS[7][27] , \REGISTERS[7][26] ,
         \REGISTERS[7][25] , \REGISTERS[7][24] , \REGISTERS[7][23] ,
         \REGISTERS[7][22] , \REGISTERS[7][21] , \REGISTERS[7][20] ,
         \REGISTERS[7][19] , \REGISTERS[7][18] , \REGISTERS[7][17] ,
         \REGISTERS[7][16] , \REGISTERS[7][15] , \REGISTERS[7][14] ,
         \REGISTERS[7][13] , \REGISTERS[7][12] , \REGISTERS[7][11] ,
         \REGISTERS[7][10] , \REGISTERS[7][9] , \REGISTERS[7][8] ,
         \REGISTERS[7][7] , \REGISTERS[7][6] , \REGISTERS[7][5] ,
         \REGISTERS[7][4] , \REGISTERS[7][3] , \REGISTERS[7][2] ,
         \REGISTERS[7][1] , \REGISTERS[7][0] , \REGISTERS[6][31] ,
         \REGISTERS[6][30] , \REGISTERS[6][29] , \REGISTERS[6][28] ,
         \REGISTERS[6][27] , \REGISTERS[6][26] , \REGISTERS[6][25] ,
         \REGISTERS[6][24] , \REGISTERS[6][23] , \REGISTERS[6][22] ,
         \REGISTERS[6][21] , \REGISTERS[6][20] , \REGISTERS[6][19] ,
         \REGISTERS[6][18] , \REGISTERS[6][17] , \REGISTERS[6][16] ,
         \REGISTERS[6][15] , \REGISTERS[6][14] , \REGISTERS[6][13] ,
         \REGISTERS[6][12] , \REGISTERS[6][11] , \REGISTERS[6][10] ,
         \REGISTERS[6][9] , \REGISTERS[6][8] , \REGISTERS[6][7] ,
         \REGISTERS[6][6] , \REGISTERS[6][5] , \REGISTERS[6][4] ,
         \REGISTERS[6][3] , \REGISTERS[6][2] , \REGISTERS[6][1] ,
         \REGISTERS[6][0] , \REGISTERS[5][31] , \REGISTERS[5][30] ,
         \REGISTERS[5][29] , \REGISTERS[5][28] , \REGISTERS[5][27] ,
         \REGISTERS[5][26] , \REGISTERS[5][25] , \REGISTERS[5][24] ,
         \REGISTERS[5][23] , \REGISTERS[5][22] , \REGISTERS[5][21] ,
         \REGISTERS[5][20] , \REGISTERS[5][19] , \REGISTERS[5][18] ,
         \REGISTERS[5][17] , \REGISTERS[5][16] , \REGISTERS[5][15] ,
         \REGISTERS[5][14] , \REGISTERS[5][13] , \REGISTERS[5][12] ,
         \REGISTERS[5][11] , \REGISTERS[5][10] , \REGISTERS[5][9] ,
         \REGISTERS[5][8] , \REGISTERS[5][7] , \REGISTERS[5][6] ,
         \REGISTERS[5][5] , \REGISTERS[5][4] , \REGISTERS[5][3] ,
         \REGISTERS[5][2] , \REGISTERS[5][1] , \REGISTERS[5][0] ,
         \REGISTERS[4][31] , \REGISTERS[4][30] , \REGISTERS[4][29] ,
         \REGISTERS[4][28] , \REGISTERS[4][27] , \REGISTERS[4][26] ,
         \REGISTERS[4][25] , \REGISTERS[4][24] , \REGISTERS[4][23] ,
         \REGISTERS[4][22] , \REGISTERS[4][21] , \REGISTERS[4][20] ,
         \REGISTERS[4][19] , \REGISTERS[4][18] , \REGISTERS[4][17] ,
         \REGISTERS[4][16] , \REGISTERS[4][15] , \REGISTERS[4][14] ,
         \REGISTERS[4][13] , \REGISTERS[4][12] , \REGISTERS[4][11] ,
         \REGISTERS[4][10] , \REGISTERS[4][9] , \REGISTERS[4][8] ,
         \REGISTERS[4][7] , \REGISTERS[4][6] , \REGISTERS[4][5] ,
         \REGISTERS[4][4] , \REGISTERS[4][3] , \REGISTERS[4][2] ,
         \REGISTERS[4][1] , \REGISTERS[4][0] , \REGISTERS[3][31] ,
         \REGISTERS[3][30] , \REGISTERS[3][29] , \REGISTERS[3][28] ,
         \REGISTERS[3][27] , \REGISTERS[3][26] , \REGISTERS[3][25] ,
         \REGISTERS[3][24] , \REGISTERS[3][23] , \REGISTERS[3][22] ,
         \REGISTERS[3][21] , \REGISTERS[3][20] , \REGISTERS[3][19] ,
         \REGISTERS[3][18] , \REGISTERS[3][17] , \REGISTERS[3][16] ,
         \REGISTERS[3][15] , \REGISTERS[3][14] , \REGISTERS[3][13] ,
         \REGISTERS[3][12] , \REGISTERS[3][11] , \REGISTERS[3][10] ,
         \REGISTERS[3][9] , \REGISTERS[3][8] , \REGISTERS[3][7] ,
         \REGISTERS[3][6] , \REGISTERS[3][5] , \REGISTERS[3][4] ,
         \REGISTERS[3][3] , \REGISTERS[3][2] , \REGISTERS[3][1] ,
         \REGISTERS[3][0] , \REGISTERS[2][31] , \REGISTERS[2][30] ,
         \REGISTERS[2][29] , \REGISTERS[2][28] , \REGISTERS[2][27] ,
         \REGISTERS[2][26] , \REGISTERS[2][25] , \REGISTERS[2][24] ,
         \REGISTERS[2][23] , \REGISTERS[2][22] , \REGISTERS[2][21] ,
         \REGISTERS[2][20] , \REGISTERS[2][19] , \REGISTERS[2][18] ,
         \REGISTERS[2][17] , \REGISTERS[2][16] , \REGISTERS[2][15] ,
         \REGISTERS[2][14] , \REGISTERS[2][13] , \REGISTERS[2][12] ,
         \REGISTERS[2][11] , \REGISTERS[2][10] , \REGISTERS[2][9] ,
         \REGISTERS[2][8] , \REGISTERS[2][7] , \REGISTERS[2][6] ,
         \REGISTERS[2][5] , \REGISTERS[2][4] , \REGISTERS[2][3] ,
         \REGISTERS[2][2] , \REGISTERS[2][1] , \REGISTERS[2][0] ,
         \REGISTERS[1][31] , \REGISTERS[1][30] , \REGISTERS[1][29] ,
         \REGISTERS[1][28] , \REGISTERS[1][27] , \REGISTERS[1][26] ,
         \REGISTERS[1][25] , \REGISTERS[1][24] , \REGISTERS[1][23] ,
         \REGISTERS[1][22] , \REGISTERS[1][21] , \REGISTERS[1][20] ,
         \REGISTERS[1][19] , \REGISTERS[1][18] , \REGISTERS[1][17] ,
         \REGISTERS[1][16] , \REGISTERS[1][15] , \REGISTERS[1][14] ,
         \REGISTERS[1][13] , \REGISTERS[1][12] , \REGISTERS[1][11] ,
         \REGISTERS[1][10] , \REGISTERS[1][9] , \REGISTERS[1][8] ,
         \REGISTERS[1][7] , \REGISTERS[1][6] , \REGISTERS[1][5] ,
         \REGISTERS[1][4] , \REGISTERS[1][3] , \REGISTERS[1][2] ,
         \REGISTERS[1][1] , \REGISTERS[1][0] , \REGISTERS[0][31] ,
         \REGISTERS[0][30] , \REGISTERS[0][29] , \REGISTERS[0][28] ,
         \REGISTERS[0][27] , \REGISTERS[0][26] , \REGISTERS[0][25] ,
         \REGISTERS[0][24] , \REGISTERS[0][23] , \REGISTERS[0][22] ,
         \REGISTERS[0][21] , \REGISTERS[0][20] , \REGISTERS[0][19] ,
         \REGISTERS[0][18] , \REGISTERS[0][17] , \REGISTERS[0][16] ,
         \REGISTERS[0][15] , \REGISTERS[0][14] , \REGISTERS[0][13] ,
         \REGISTERS[0][12] , \REGISTERS[0][11] , \REGISTERS[0][10] ,
         \REGISTERS[0][9] , \REGISTERS[0][8] , \REGISTERS[0][7] ,
         \REGISTERS[0][6] , \REGISTERS[0][5] , \REGISTERS[0][4] ,
         \REGISTERS[0][3] , \REGISTERS[0][2] , \REGISTERS[0][1] ,
         \REGISTERS[0][0] , N1072, N1394, N1458, N1522, N1586, N1650, N1714,
         N1778, N1842, N1906, N1970, N2034, N2098, N2162, N2226, N2290, N2354,
         N2418, N2482, N2546, N2610, N2674, N2738, N2802, N2866, N2930, N2994,
         N3058, N3122, N3186, N3250, N3314, N3317, N3319, N3321, N3323, N3325,
         N3327, N3329, N3331, N3333, N3335, N3337, N3339, N3341, N3343, N3345,
         N3347, N3349, N3351, N3353, N3355, N3357, N3359, N3361, N3363, N3365,
         N3367, N3369, N3371, N3373, N3375, N3377, N3378, N3379, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n1, n1229, n1270, n1876, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306;

  DLH_X1 \REGISTERS_reg[31][31]  ( .G(n2211), .D(N3379), .Q(
        \REGISTERS[31][31] ) );
  DLH_X1 \REGISTERS_reg[31][30]  ( .G(n2211), .D(N3377), .Q(
        \REGISTERS[31][30] ) );
  DLH_X1 \REGISTERS_reg[31][29]  ( .G(n2211), .D(N3375), .Q(
        \REGISTERS[31][29] ) );
  DLH_X1 \REGISTERS_reg[31][28]  ( .G(n2211), .D(N3373), .Q(
        \REGISTERS[31][28] ) );
  DLH_X1 \REGISTERS_reg[31][27]  ( .G(n2211), .D(N3371), .Q(
        \REGISTERS[31][27] ) );
  DLH_X1 \REGISTERS_reg[31][26]  ( .G(n2211), .D(N3369), .Q(
        \REGISTERS[31][26] ) );
  DLH_X1 \REGISTERS_reg[31][25]  ( .G(n2211), .D(N3367), .Q(
        \REGISTERS[31][25] ) );
  DLH_X1 \REGISTERS_reg[31][24]  ( .G(n2211), .D(N3365), .Q(
        \REGISTERS[31][24] ) );
  DLH_X1 \REGISTERS_reg[31][23]  ( .G(n2211), .D(N3363), .Q(
        \REGISTERS[31][23] ) );
  DLH_X1 \REGISTERS_reg[31][22]  ( .G(n2211), .D(N3361), .Q(
        \REGISTERS[31][22] ) );
  DLH_X1 \REGISTERS_reg[31][21]  ( .G(n2211), .D(N3359), .Q(
        \REGISTERS[31][21] ) );
  DLH_X1 \REGISTERS_reg[31][20]  ( .G(n2211), .D(N3357), .Q(
        \REGISTERS[31][20] ) );
  DLH_X1 \REGISTERS_reg[31][19]  ( .G(n2211), .D(N3355), .Q(
        \REGISTERS[31][19] ) );
  DLH_X1 \REGISTERS_reg[31][18]  ( .G(n2212), .D(N3353), .Q(
        \REGISTERS[31][18] ) );
  DLH_X1 \REGISTERS_reg[31][17]  ( .G(n2212), .D(N3351), .Q(
        \REGISTERS[31][17] ) );
  DLH_X1 \REGISTERS_reg[31][16]  ( .G(n2212), .D(N3349), .Q(
        \REGISTERS[31][16] ) );
  DLH_X1 \REGISTERS_reg[31][15]  ( .G(n2212), .D(N3347), .Q(
        \REGISTERS[31][15] ) );
  DLH_X1 \REGISTERS_reg[31][14]  ( .G(n2212), .D(N3345), .Q(
        \REGISTERS[31][14] ) );
  DLH_X1 \REGISTERS_reg[31][13]  ( .G(n2212), .D(N3343), .Q(
        \REGISTERS[31][13] ) );
  DLH_X1 \REGISTERS_reg[31][12]  ( .G(n2212), .D(N3341), .Q(
        \REGISTERS[31][12] ) );
  DLH_X1 \REGISTERS_reg[31][11]  ( .G(n2212), .D(N3339), .Q(
        \REGISTERS[31][11] ) );
  DLH_X1 \REGISTERS_reg[31][10]  ( .G(n2212), .D(N3337), .Q(
        \REGISTERS[31][10] ) );
  DLH_X1 \REGISTERS_reg[31][9]  ( .G(n2212), .D(N3335), .Q(\REGISTERS[31][9] )
         );
  DLH_X1 \REGISTERS_reg[31][8]  ( .G(n2212), .D(N3333), .Q(\REGISTERS[31][8] )
         );
  DLH_X1 \REGISTERS_reg[31][7]  ( .G(n2212), .D(N3331), .Q(\REGISTERS[31][7] )
         );
  DLH_X1 \REGISTERS_reg[31][6]  ( .G(n2212), .D(N3329), .Q(\REGISTERS[31][6] )
         );
  DLH_X1 \REGISTERS_reg[31][5]  ( .G(n2213), .D(N3327), .Q(\REGISTERS[31][5] )
         );
  DLH_X1 \REGISTERS_reg[31][4]  ( .G(n2213), .D(N3325), .Q(\REGISTERS[31][4] )
         );
  DLH_X1 \REGISTERS_reg[31][3]  ( .G(n2213), .D(N3323), .Q(\REGISTERS[31][3] )
         );
  DLH_X1 \REGISTERS_reg[31][2]  ( .G(n2213), .D(N3321), .Q(\REGISTERS[31][2] )
         );
  DLH_X1 \REGISTERS_reg[31][1]  ( .G(n2213), .D(N3319), .Q(\REGISTERS[31][1] )
         );
  DLH_X1 \REGISTERS_reg[31][0]  ( .G(n2213), .D(N3317), .Q(\REGISTERS[31][0] )
         );
  DLH_X1 \REGISTERS_reg[30][31]  ( .G(n2214), .D(n1948), .Q(
        \REGISTERS[30][31] ) );
  DLH_X1 \REGISTERS_reg[30][30]  ( .G(n2214), .D(n1947), .Q(
        \REGISTERS[30][30] ) );
  DLH_X1 \REGISTERS_reg[30][29]  ( .G(n2214), .D(n1946), .Q(
        \REGISTERS[30][29] ) );
  DLH_X1 \REGISTERS_reg[30][28]  ( .G(n2214), .D(n1945), .Q(
        \REGISTERS[30][28] ) );
  DLH_X1 \REGISTERS_reg[30][27]  ( .G(n2214), .D(n1944), .Q(
        \REGISTERS[30][27] ) );
  DLH_X1 \REGISTERS_reg[30][26]  ( .G(n2214), .D(n1943), .Q(
        \REGISTERS[30][26] ) );
  DLH_X1 \REGISTERS_reg[30][25]  ( .G(n2214), .D(n1942), .Q(
        \REGISTERS[30][25] ) );
  DLH_X1 \REGISTERS_reg[30][24]  ( .G(n2214), .D(n1941), .Q(
        \REGISTERS[30][24] ) );
  DLH_X1 \REGISTERS_reg[30][23]  ( .G(n2214), .D(n1940), .Q(
        \REGISTERS[30][23] ) );
  DLH_X1 \REGISTERS_reg[30][22]  ( .G(n2214), .D(n1939), .Q(
        \REGISTERS[30][22] ) );
  DLH_X1 \REGISTERS_reg[30][21]  ( .G(n2214), .D(n1938), .Q(
        \REGISTERS[30][21] ) );
  DLH_X1 \REGISTERS_reg[30][20]  ( .G(n2214), .D(n1937), .Q(
        \REGISTERS[30][20] ) );
  DLH_X1 \REGISTERS_reg[30][19]  ( .G(n2214), .D(n1936), .Q(
        \REGISTERS[30][19] ) );
  DLH_X1 \REGISTERS_reg[30][18]  ( .G(n2215), .D(n1935), .Q(
        \REGISTERS[30][18] ) );
  DLH_X1 \REGISTERS_reg[30][17]  ( .G(n2215), .D(n1934), .Q(
        \REGISTERS[30][17] ) );
  DLH_X1 \REGISTERS_reg[30][16]  ( .G(n2215), .D(n1933), .Q(
        \REGISTERS[30][16] ) );
  DLH_X1 \REGISTERS_reg[30][15]  ( .G(n2215), .D(n1932), .Q(
        \REGISTERS[30][15] ) );
  DLH_X1 \REGISTERS_reg[30][14]  ( .G(n2215), .D(n1931), .Q(
        \REGISTERS[30][14] ) );
  DLH_X1 \REGISTERS_reg[30][13]  ( .G(n2215), .D(n1930), .Q(
        \REGISTERS[30][13] ) );
  DLH_X1 \REGISTERS_reg[30][12]  ( .G(n2215), .D(n1929), .Q(
        \REGISTERS[30][12] ) );
  DLH_X1 \REGISTERS_reg[30][11]  ( .G(n2215), .D(n1928), .Q(
        \REGISTERS[30][11] ) );
  DLH_X1 \REGISTERS_reg[30][10]  ( .G(n2215), .D(n1927), .Q(
        \REGISTERS[30][10] ) );
  DLH_X1 \REGISTERS_reg[30][9]  ( .G(n2215), .D(n1926), .Q(\REGISTERS[30][9] )
         );
  DLH_X1 \REGISTERS_reg[30][8]  ( .G(n2215), .D(n1925), .Q(\REGISTERS[30][8] )
         );
  DLH_X1 \REGISTERS_reg[30][7]  ( .G(n2215), .D(n1924), .Q(\REGISTERS[30][7] )
         );
  DLH_X1 \REGISTERS_reg[30][6]  ( .G(n2215), .D(n1923), .Q(\REGISTERS[30][6] )
         );
  DLH_X1 \REGISTERS_reg[30][5]  ( .G(n2216), .D(n1922), .Q(\REGISTERS[30][5] )
         );
  DLH_X1 \REGISTERS_reg[30][4]  ( .G(n2216), .D(n1921), .Q(\REGISTERS[30][4] )
         );
  DLH_X1 \REGISTERS_reg[30][3]  ( .G(n2216), .D(n1920), .Q(\REGISTERS[30][3] )
         );
  DLH_X1 \REGISTERS_reg[30][2]  ( .G(n2216), .D(n1919), .Q(\REGISTERS[30][2] )
         );
  DLH_X1 \REGISTERS_reg[30][1]  ( .G(n2216), .D(n1918), .Q(\REGISTERS[30][1] )
         );
  DLH_X1 \REGISTERS_reg[30][0]  ( .G(n2216), .D(n1917), .Q(\REGISTERS[30][0] )
         );
  DLH_X1 \REGISTERS_reg[29][31]  ( .G(n2217), .D(N3379), .Q(
        \REGISTERS[29][31] ) );
  DLH_X1 \REGISTERS_reg[29][30]  ( .G(n2217), .D(N3377), .Q(
        \REGISTERS[29][30] ) );
  DLH_X1 \REGISTERS_reg[29][29]  ( .G(n2217), .D(N3375), .Q(
        \REGISTERS[29][29] ) );
  DLH_X1 \REGISTERS_reg[29][28]  ( .G(n2217), .D(N3373), .Q(
        \REGISTERS[29][28] ) );
  DLH_X1 \REGISTERS_reg[29][27]  ( .G(n2217), .D(N3371), .Q(
        \REGISTERS[29][27] ) );
  DLH_X1 \REGISTERS_reg[29][26]  ( .G(n2217), .D(N3369), .Q(
        \REGISTERS[29][26] ) );
  DLH_X1 \REGISTERS_reg[29][25]  ( .G(n2217), .D(N3367), .Q(
        \REGISTERS[29][25] ) );
  DLH_X1 \REGISTERS_reg[29][24]  ( .G(n2217), .D(N3365), .Q(
        \REGISTERS[29][24] ) );
  DLH_X1 \REGISTERS_reg[29][23]  ( .G(n2217), .D(N3363), .Q(
        \REGISTERS[29][23] ) );
  DLH_X1 \REGISTERS_reg[29][22]  ( .G(n2217), .D(N3361), .Q(
        \REGISTERS[29][22] ) );
  DLH_X1 \REGISTERS_reg[29][21]  ( .G(n2217), .D(N3359), .Q(
        \REGISTERS[29][21] ) );
  DLH_X1 \REGISTERS_reg[29][20]  ( .G(n2217), .D(N3357), .Q(
        \REGISTERS[29][20] ) );
  DLH_X1 \REGISTERS_reg[29][19]  ( .G(n2217), .D(N3355), .Q(
        \REGISTERS[29][19] ) );
  DLH_X1 \REGISTERS_reg[29][18]  ( .G(n2218), .D(N3353), .Q(
        \REGISTERS[29][18] ) );
  DLH_X1 \REGISTERS_reg[29][17]  ( .G(n2218), .D(N3351), .Q(
        \REGISTERS[29][17] ) );
  DLH_X1 \REGISTERS_reg[29][16]  ( .G(n2218), .D(N3349), .Q(
        \REGISTERS[29][16] ) );
  DLH_X1 \REGISTERS_reg[29][15]  ( .G(n2218), .D(N3347), .Q(
        \REGISTERS[29][15] ) );
  DLH_X1 \REGISTERS_reg[29][14]  ( .G(n2218), .D(N3345), .Q(
        \REGISTERS[29][14] ) );
  DLH_X1 \REGISTERS_reg[29][13]  ( .G(n2218), .D(N3343), .Q(
        \REGISTERS[29][13] ) );
  DLH_X1 \REGISTERS_reg[29][12]  ( .G(n2218), .D(N3341), .Q(
        \REGISTERS[29][12] ) );
  DLH_X1 \REGISTERS_reg[29][11]  ( .G(n2218), .D(N3339), .Q(
        \REGISTERS[29][11] ) );
  DLH_X1 \REGISTERS_reg[29][10]  ( .G(n2218), .D(N3337), .Q(
        \REGISTERS[29][10] ) );
  DLH_X1 \REGISTERS_reg[29][9]  ( .G(n2218), .D(N3335), .Q(\REGISTERS[29][9] )
         );
  DLH_X1 \REGISTERS_reg[29][8]  ( .G(n2218), .D(N3333), .Q(\REGISTERS[29][8] )
         );
  DLH_X1 \REGISTERS_reg[29][7]  ( .G(n2218), .D(N3331), .Q(\REGISTERS[29][7] )
         );
  DLH_X1 \REGISTERS_reg[29][6]  ( .G(n2218), .D(N3329), .Q(\REGISTERS[29][6] )
         );
  DLH_X1 \REGISTERS_reg[29][5]  ( .G(n2219), .D(N3327), .Q(\REGISTERS[29][5] )
         );
  DLH_X1 \REGISTERS_reg[29][4]  ( .G(n2219), .D(N3325), .Q(\REGISTERS[29][4] )
         );
  DLH_X1 \REGISTERS_reg[29][3]  ( .G(n2219), .D(N3323), .Q(\REGISTERS[29][3] )
         );
  DLH_X1 \REGISTERS_reg[29][2]  ( .G(n2219), .D(N3321), .Q(\REGISTERS[29][2] )
         );
  DLH_X1 \REGISTERS_reg[29][1]  ( .G(n2219), .D(N3319), .Q(\REGISTERS[29][1] )
         );
  DLH_X1 \REGISTERS_reg[29][0]  ( .G(n2219), .D(N3317), .Q(\REGISTERS[29][0] )
         );
  DLH_X1 \REGISTERS_reg[28][31]  ( .G(n2220), .D(n1948), .Q(
        \REGISTERS[28][31] ) );
  DLH_X1 \REGISTERS_reg[28][30]  ( .G(n2220), .D(n1947), .Q(
        \REGISTERS[28][30] ) );
  DLH_X1 \REGISTERS_reg[28][29]  ( .G(n2220), .D(n1946), .Q(
        \REGISTERS[28][29] ) );
  DLH_X1 \REGISTERS_reg[28][28]  ( .G(n2220), .D(n1945), .Q(
        \REGISTERS[28][28] ) );
  DLH_X1 \REGISTERS_reg[28][27]  ( .G(n2220), .D(n1944), .Q(
        \REGISTERS[28][27] ) );
  DLH_X1 \REGISTERS_reg[28][26]  ( .G(n2220), .D(n1943), .Q(
        \REGISTERS[28][26] ) );
  DLH_X1 \REGISTERS_reg[28][25]  ( .G(n2220), .D(n1942), .Q(
        \REGISTERS[28][25] ) );
  DLH_X1 \REGISTERS_reg[28][24]  ( .G(n2220), .D(n1941), .Q(
        \REGISTERS[28][24] ) );
  DLH_X1 \REGISTERS_reg[28][23]  ( .G(n2220), .D(n1940), .Q(
        \REGISTERS[28][23] ) );
  DLH_X1 \REGISTERS_reg[28][22]  ( .G(n2220), .D(n1939), .Q(
        \REGISTERS[28][22] ) );
  DLH_X1 \REGISTERS_reg[28][21]  ( .G(n2220), .D(n1938), .Q(
        \REGISTERS[28][21] ) );
  DLH_X1 \REGISTERS_reg[28][20]  ( .G(n2220), .D(n1937), .Q(
        \REGISTERS[28][20] ) );
  DLH_X1 \REGISTERS_reg[28][19]  ( .G(n2220), .D(n1936), .Q(
        \REGISTERS[28][19] ) );
  DLH_X1 \REGISTERS_reg[28][18]  ( .G(n2221), .D(n1935), .Q(
        \REGISTERS[28][18] ) );
  DLH_X1 \REGISTERS_reg[28][17]  ( .G(n2221), .D(n1934), .Q(
        \REGISTERS[28][17] ) );
  DLH_X1 \REGISTERS_reg[28][16]  ( .G(n2221), .D(n1933), .Q(
        \REGISTERS[28][16] ) );
  DLH_X1 \REGISTERS_reg[28][15]  ( .G(n2221), .D(n1932), .Q(
        \REGISTERS[28][15] ) );
  DLH_X1 \REGISTERS_reg[28][14]  ( .G(n2221), .D(n1931), .Q(
        \REGISTERS[28][14] ) );
  DLH_X1 \REGISTERS_reg[28][13]  ( .G(n2221), .D(n1930), .Q(
        \REGISTERS[28][13] ) );
  DLH_X1 \REGISTERS_reg[28][12]  ( .G(n2221), .D(n1929), .Q(
        \REGISTERS[28][12] ) );
  DLH_X1 \REGISTERS_reg[28][11]  ( .G(n2221), .D(n1928), .Q(
        \REGISTERS[28][11] ) );
  DLH_X1 \REGISTERS_reg[28][10]  ( .G(n2221), .D(n1927), .Q(
        \REGISTERS[28][10] ) );
  DLH_X1 \REGISTERS_reg[28][9]  ( .G(n2221), .D(n1926), .Q(\REGISTERS[28][9] )
         );
  DLH_X1 \REGISTERS_reg[28][8]  ( .G(n2221), .D(n1925), .Q(\REGISTERS[28][8] )
         );
  DLH_X1 \REGISTERS_reg[28][7]  ( .G(n2221), .D(n1924), .Q(\REGISTERS[28][7] )
         );
  DLH_X1 \REGISTERS_reg[28][6]  ( .G(n2221), .D(n1923), .Q(\REGISTERS[28][6] )
         );
  DLH_X1 \REGISTERS_reg[28][5]  ( .G(n2222), .D(n1922), .Q(\REGISTERS[28][5] )
         );
  DLH_X1 \REGISTERS_reg[28][4]  ( .G(n2222), .D(n1921), .Q(\REGISTERS[28][4] )
         );
  DLH_X1 \REGISTERS_reg[28][3]  ( .G(n2222), .D(n1920), .Q(\REGISTERS[28][3] )
         );
  DLH_X1 \REGISTERS_reg[28][2]  ( .G(n2222), .D(n1919), .Q(\REGISTERS[28][2] )
         );
  DLH_X1 \REGISTERS_reg[28][1]  ( .G(n2222), .D(n1918), .Q(\REGISTERS[28][1] )
         );
  DLH_X1 \REGISTERS_reg[28][0]  ( .G(n2222), .D(n1917), .Q(\REGISTERS[28][0] )
         );
  DLH_X1 \REGISTERS_reg[27][31]  ( .G(n2223), .D(N3379), .Q(
        \REGISTERS[27][31] ) );
  DLH_X1 \REGISTERS_reg[27][30]  ( .G(n2223), .D(N3377), .Q(
        \REGISTERS[27][30] ) );
  DLH_X1 \REGISTERS_reg[27][29]  ( .G(n2223), .D(N3375), .Q(
        \REGISTERS[27][29] ) );
  DLH_X1 \REGISTERS_reg[27][28]  ( .G(n2223), .D(N3373), .Q(
        \REGISTERS[27][28] ) );
  DLH_X1 \REGISTERS_reg[27][27]  ( .G(n2223), .D(N3371), .Q(
        \REGISTERS[27][27] ) );
  DLH_X1 \REGISTERS_reg[27][26]  ( .G(n2223), .D(N3369), .Q(
        \REGISTERS[27][26] ) );
  DLH_X1 \REGISTERS_reg[27][25]  ( .G(n2223), .D(N3367), .Q(
        \REGISTERS[27][25] ) );
  DLH_X1 \REGISTERS_reg[27][24]  ( .G(n2223), .D(N3365), .Q(
        \REGISTERS[27][24] ) );
  DLH_X1 \REGISTERS_reg[27][23]  ( .G(n2223), .D(N3363), .Q(
        \REGISTERS[27][23] ) );
  DLH_X1 \REGISTERS_reg[27][22]  ( .G(n2223), .D(N3361), .Q(
        \REGISTERS[27][22] ) );
  DLH_X1 \REGISTERS_reg[27][21]  ( .G(n2223), .D(N3359), .Q(
        \REGISTERS[27][21] ) );
  DLH_X1 \REGISTERS_reg[27][20]  ( .G(n2223), .D(N3357), .Q(
        \REGISTERS[27][20] ) );
  DLH_X1 \REGISTERS_reg[27][19]  ( .G(n2223), .D(N3355), .Q(
        \REGISTERS[27][19] ) );
  DLH_X1 \REGISTERS_reg[27][18]  ( .G(n2224), .D(N3353), .Q(
        \REGISTERS[27][18] ) );
  DLH_X1 \REGISTERS_reg[27][17]  ( .G(n2224), .D(N3351), .Q(
        \REGISTERS[27][17] ) );
  DLH_X1 \REGISTERS_reg[27][16]  ( .G(n2224), .D(N3349), .Q(
        \REGISTERS[27][16] ) );
  DLH_X1 \REGISTERS_reg[27][15]  ( .G(n2224), .D(N3347), .Q(
        \REGISTERS[27][15] ) );
  DLH_X1 \REGISTERS_reg[27][14]  ( .G(n2224), .D(N3345), .Q(
        \REGISTERS[27][14] ) );
  DLH_X1 \REGISTERS_reg[27][13]  ( .G(n2224), .D(N3343), .Q(
        \REGISTERS[27][13] ) );
  DLH_X1 \REGISTERS_reg[27][12]  ( .G(n2224), .D(N3341), .Q(
        \REGISTERS[27][12] ) );
  DLH_X1 \REGISTERS_reg[27][11]  ( .G(n2224), .D(N3339), .Q(
        \REGISTERS[27][11] ) );
  DLH_X1 \REGISTERS_reg[27][10]  ( .G(n2224), .D(N3337), .Q(
        \REGISTERS[27][10] ) );
  DLH_X1 \REGISTERS_reg[27][9]  ( .G(n2224), .D(N3335), .Q(\REGISTERS[27][9] )
         );
  DLH_X1 \REGISTERS_reg[27][8]  ( .G(n2224), .D(N3333), .Q(\REGISTERS[27][8] )
         );
  DLH_X1 \REGISTERS_reg[27][7]  ( .G(n2224), .D(N3331), .Q(\REGISTERS[27][7] )
         );
  DLH_X1 \REGISTERS_reg[27][6]  ( .G(n2224), .D(N3329), .Q(\REGISTERS[27][6] )
         );
  DLH_X1 \REGISTERS_reg[27][5]  ( .G(n2225), .D(N3327), .Q(\REGISTERS[27][5] )
         );
  DLH_X1 \REGISTERS_reg[27][4]  ( .G(n2225), .D(N3325), .Q(\REGISTERS[27][4] )
         );
  DLH_X1 \REGISTERS_reg[27][3]  ( .G(n2225), .D(N3323), .Q(\REGISTERS[27][3] )
         );
  DLH_X1 \REGISTERS_reg[27][2]  ( .G(n2225), .D(N3321), .Q(\REGISTERS[27][2] )
         );
  DLH_X1 \REGISTERS_reg[27][1]  ( .G(n2225), .D(N3319), .Q(\REGISTERS[27][1] )
         );
  DLH_X1 \REGISTERS_reg[27][0]  ( .G(n2225), .D(N3317), .Q(\REGISTERS[27][0] )
         );
  DLH_X1 \REGISTERS_reg[26][31]  ( .G(n2226), .D(n1948), .Q(
        \REGISTERS[26][31] ) );
  DLH_X1 \REGISTERS_reg[26][30]  ( .G(n2226), .D(n1947), .Q(
        \REGISTERS[26][30] ) );
  DLH_X1 \REGISTERS_reg[26][29]  ( .G(n2226), .D(n1946), .Q(
        \REGISTERS[26][29] ) );
  DLH_X1 \REGISTERS_reg[26][28]  ( .G(n2226), .D(n1945), .Q(
        \REGISTERS[26][28] ) );
  DLH_X1 \REGISTERS_reg[26][27]  ( .G(n2226), .D(n1944), .Q(
        \REGISTERS[26][27] ) );
  DLH_X1 \REGISTERS_reg[26][26]  ( .G(n2226), .D(n1943), .Q(
        \REGISTERS[26][26] ) );
  DLH_X1 \REGISTERS_reg[26][25]  ( .G(n2226), .D(n1942), .Q(
        \REGISTERS[26][25] ) );
  DLH_X1 \REGISTERS_reg[26][24]  ( .G(n2226), .D(n1941), .Q(
        \REGISTERS[26][24] ) );
  DLH_X1 \REGISTERS_reg[26][23]  ( .G(n2226), .D(n1940), .Q(
        \REGISTERS[26][23] ) );
  DLH_X1 \REGISTERS_reg[26][22]  ( .G(n2226), .D(n1939), .Q(
        \REGISTERS[26][22] ) );
  DLH_X1 \REGISTERS_reg[26][21]  ( .G(n2226), .D(n1938), .Q(
        \REGISTERS[26][21] ) );
  DLH_X1 \REGISTERS_reg[26][20]  ( .G(n2226), .D(n1937), .Q(
        \REGISTERS[26][20] ) );
  DLH_X1 \REGISTERS_reg[26][19]  ( .G(n2226), .D(n1936), .Q(
        \REGISTERS[26][19] ) );
  DLH_X1 \REGISTERS_reg[26][18]  ( .G(n2227), .D(n1935), .Q(
        \REGISTERS[26][18] ) );
  DLH_X1 \REGISTERS_reg[26][17]  ( .G(n2227), .D(n1934), .Q(
        \REGISTERS[26][17] ) );
  DLH_X1 \REGISTERS_reg[26][16]  ( .G(n2227), .D(n1933), .Q(
        \REGISTERS[26][16] ) );
  DLH_X1 \REGISTERS_reg[26][15]  ( .G(n2227), .D(n1932), .Q(
        \REGISTERS[26][15] ) );
  DLH_X1 \REGISTERS_reg[26][14]  ( .G(n2227), .D(n1931), .Q(
        \REGISTERS[26][14] ) );
  DLH_X1 \REGISTERS_reg[26][13]  ( .G(n2227), .D(n1930), .Q(
        \REGISTERS[26][13] ) );
  DLH_X1 \REGISTERS_reg[26][12]  ( .G(n2227), .D(n1929), .Q(
        \REGISTERS[26][12] ) );
  DLH_X1 \REGISTERS_reg[26][11]  ( .G(n2227), .D(n1928), .Q(
        \REGISTERS[26][11] ) );
  DLH_X1 \REGISTERS_reg[26][10]  ( .G(n2227), .D(n1927), .Q(
        \REGISTERS[26][10] ) );
  DLH_X1 \REGISTERS_reg[26][9]  ( .G(n2227), .D(n1926), .Q(\REGISTERS[26][9] )
         );
  DLH_X1 \REGISTERS_reg[26][8]  ( .G(n2227), .D(n1925), .Q(\REGISTERS[26][8] )
         );
  DLH_X1 \REGISTERS_reg[26][7]  ( .G(n2227), .D(n1924), .Q(\REGISTERS[26][7] )
         );
  DLH_X1 \REGISTERS_reg[26][6]  ( .G(n2227), .D(n1923), .Q(\REGISTERS[26][6] )
         );
  DLH_X1 \REGISTERS_reg[26][5]  ( .G(n2228), .D(n1922), .Q(\REGISTERS[26][5] )
         );
  DLH_X1 \REGISTERS_reg[26][4]  ( .G(n2228), .D(n1921), .Q(\REGISTERS[26][4] )
         );
  DLH_X1 \REGISTERS_reg[26][3]  ( .G(n2228), .D(n1920), .Q(\REGISTERS[26][3] )
         );
  DLH_X1 \REGISTERS_reg[26][2]  ( .G(n2228), .D(n1919), .Q(\REGISTERS[26][2] )
         );
  DLH_X1 \REGISTERS_reg[26][1]  ( .G(n2228), .D(n1918), .Q(\REGISTERS[26][1] )
         );
  DLH_X1 \REGISTERS_reg[26][0]  ( .G(n2228), .D(n1917), .Q(\REGISTERS[26][0] )
         );
  DLH_X1 \REGISTERS_reg[25][31]  ( .G(n2229), .D(N3379), .Q(
        \REGISTERS[25][31] ) );
  DLH_X1 \REGISTERS_reg[25][30]  ( .G(n2229), .D(N3377), .Q(
        \REGISTERS[25][30] ) );
  DLH_X1 \REGISTERS_reg[25][29]  ( .G(n2229), .D(N3375), .Q(
        \REGISTERS[25][29] ) );
  DLH_X1 \REGISTERS_reg[25][28]  ( .G(n2229), .D(N3373), .Q(
        \REGISTERS[25][28] ) );
  DLH_X1 \REGISTERS_reg[25][27]  ( .G(n2229), .D(N3371), .Q(
        \REGISTERS[25][27] ) );
  DLH_X1 \REGISTERS_reg[25][26]  ( .G(n2229), .D(N3369), .Q(
        \REGISTERS[25][26] ) );
  DLH_X1 \REGISTERS_reg[25][25]  ( .G(n2229), .D(N3367), .Q(
        \REGISTERS[25][25] ) );
  DLH_X1 \REGISTERS_reg[25][24]  ( .G(n2229), .D(N3365), .Q(
        \REGISTERS[25][24] ) );
  DLH_X1 \REGISTERS_reg[25][23]  ( .G(n2229), .D(N3363), .Q(
        \REGISTERS[25][23] ) );
  DLH_X1 \REGISTERS_reg[25][22]  ( .G(n2229), .D(N3361), .Q(
        \REGISTERS[25][22] ) );
  DLH_X1 \REGISTERS_reg[25][21]  ( .G(n2229), .D(N3359), .Q(
        \REGISTERS[25][21] ) );
  DLH_X1 \REGISTERS_reg[25][20]  ( .G(n2229), .D(N3357), .Q(
        \REGISTERS[25][20] ) );
  DLH_X1 \REGISTERS_reg[25][19]  ( .G(n2229), .D(N3355), .Q(
        \REGISTERS[25][19] ) );
  DLH_X1 \REGISTERS_reg[25][18]  ( .G(n2230), .D(N3353), .Q(
        \REGISTERS[25][18] ) );
  DLH_X1 \REGISTERS_reg[25][17]  ( .G(n2230), .D(N3351), .Q(
        \REGISTERS[25][17] ) );
  DLH_X1 \REGISTERS_reg[25][16]  ( .G(n2230), .D(N3349), .Q(
        \REGISTERS[25][16] ) );
  DLH_X1 \REGISTERS_reg[25][15]  ( .G(n2230), .D(N3347), .Q(
        \REGISTERS[25][15] ) );
  DLH_X1 \REGISTERS_reg[25][14]  ( .G(n2230), .D(N3345), .Q(
        \REGISTERS[25][14] ) );
  DLH_X1 \REGISTERS_reg[25][13]  ( .G(n2230), .D(N3343), .Q(
        \REGISTERS[25][13] ) );
  DLH_X1 \REGISTERS_reg[25][12]  ( .G(n2230), .D(N3341), .Q(
        \REGISTERS[25][12] ) );
  DLH_X1 \REGISTERS_reg[25][11]  ( .G(n2230), .D(N3339), .Q(
        \REGISTERS[25][11] ) );
  DLH_X1 \REGISTERS_reg[25][10]  ( .G(n2230), .D(N3337), .Q(
        \REGISTERS[25][10] ) );
  DLH_X1 \REGISTERS_reg[25][9]  ( .G(n2230), .D(N3335), .Q(\REGISTERS[25][9] )
         );
  DLH_X1 \REGISTERS_reg[25][8]  ( .G(n2230), .D(N3333), .Q(\REGISTERS[25][8] )
         );
  DLH_X1 \REGISTERS_reg[25][7]  ( .G(n2230), .D(N3331), .Q(\REGISTERS[25][7] )
         );
  DLH_X1 \REGISTERS_reg[25][6]  ( .G(n2230), .D(N3329), .Q(\REGISTERS[25][6] )
         );
  DLH_X1 \REGISTERS_reg[25][5]  ( .G(n2231), .D(N3327), .Q(\REGISTERS[25][5] )
         );
  DLH_X1 \REGISTERS_reg[25][4]  ( .G(n2231), .D(N3325), .Q(\REGISTERS[25][4] )
         );
  DLH_X1 \REGISTERS_reg[25][3]  ( .G(n2231), .D(N3323), .Q(\REGISTERS[25][3] )
         );
  DLH_X1 \REGISTERS_reg[25][2]  ( .G(n2231), .D(N3321), .Q(\REGISTERS[25][2] )
         );
  DLH_X1 \REGISTERS_reg[25][1]  ( .G(n2231), .D(N3319), .Q(\REGISTERS[25][1] )
         );
  DLH_X1 \REGISTERS_reg[25][0]  ( .G(n2231), .D(N3317), .Q(\REGISTERS[25][0] )
         );
  DLH_X1 \REGISTERS_reg[24][31]  ( .G(n2232), .D(n1948), .Q(
        \REGISTERS[24][31] ) );
  DLH_X1 \REGISTERS_reg[24][30]  ( .G(n2232), .D(n1947), .Q(
        \REGISTERS[24][30] ) );
  DLH_X1 \REGISTERS_reg[24][29]  ( .G(n2232), .D(n1946), .Q(
        \REGISTERS[24][29] ) );
  DLH_X1 \REGISTERS_reg[24][28]  ( .G(n2232), .D(n1945), .Q(
        \REGISTERS[24][28] ) );
  DLH_X1 \REGISTERS_reg[24][27]  ( .G(n2232), .D(n1944), .Q(
        \REGISTERS[24][27] ) );
  DLH_X1 \REGISTERS_reg[24][26]  ( .G(n2232), .D(n1943), .Q(
        \REGISTERS[24][26] ) );
  DLH_X1 \REGISTERS_reg[24][25]  ( .G(n2232), .D(n1942), .Q(
        \REGISTERS[24][25] ) );
  DLH_X1 \REGISTERS_reg[24][24]  ( .G(n2232), .D(n1941), .Q(
        \REGISTERS[24][24] ) );
  DLH_X1 \REGISTERS_reg[24][23]  ( .G(n2232), .D(n1940), .Q(
        \REGISTERS[24][23] ) );
  DLH_X1 \REGISTERS_reg[24][22]  ( .G(n2232), .D(n1939), .Q(
        \REGISTERS[24][22] ) );
  DLH_X1 \REGISTERS_reg[24][21]  ( .G(n2232), .D(n1938), .Q(
        \REGISTERS[24][21] ) );
  DLH_X1 \REGISTERS_reg[24][20]  ( .G(n2232), .D(n1937), .Q(
        \REGISTERS[24][20] ) );
  DLH_X1 \REGISTERS_reg[24][19]  ( .G(n2232), .D(n1936), .Q(
        \REGISTERS[24][19] ) );
  DLH_X1 \REGISTERS_reg[24][18]  ( .G(n2233), .D(n1935), .Q(
        \REGISTERS[24][18] ) );
  DLH_X1 \REGISTERS_reg[24][17]  ( .G(n2233), .D(n1934), .Q(
        \REGISTERS[24][17] ) );
  DLH_X1 \REGISTERS_reg[24][16]  ( .G(n2233), .D(n1933), .Q(
        \REGISTERS[24][16] ) );
  DLH_X1 \REGISTERS_reg[24][15]  ( .G(n2233), .D(n1932), .Q(
        \REGISTERS[24][15] ) );
  DLH_X1 \REGISTERS_reg[24][14]  ( .G(n2233), .D(n1931), .Q(
        \REGISTERS[24][14] ) );
  DLH_X1 \REGISTERS_reg[24][13]  ( .G(n2233), .D(n1930), .Q(
        \REGISTERS[24][13] ) );
  DLH_X1 \REGISTERS_reg[24][12]  ( .G(n2233), .D(n1929), .Q(
        \REGISTERS[24][12] ) );
  DLH_X1 \REGISTERS_reg[24][11]  ( .G(n2233), .D(n1928), .Q(
        \REGISTERS[24][11] ) );
  DLH_X1 \REGISTERS_reg[24][10]  ( .G(n2233), .D(n1927), .Q(
        \REGISTERS[24][10] ) );
  DLH_X1 \REGISTERS_reg[24][9]  ( .G(n2233), .D(n1926), .Q(\REGISTERS[24][9] )
         );
  DLH_X1 \REGISTERS_reg[24][8]  ( .G(n2233), .D(n1925), .Q(\REGISTERS[24][8] )
         );
  DLH_X1 \REGISTERS_reg[24][7]  ( .G(n2233), .D(n1924), .Q(\REGISTERS[24][7] )
         );
  DLH_X1 \REGISTERS_reg[24][6]  ( .G(n2233), .D(n1923), .Q(\REGISTERS[24][6] )
         );
  DLH_X1 \REGISTERS_reg[24][5]  ( .G(n2234), .D(n1922), .Q(\REGISTERS[24][5] )
         );
  DLH_X1 \REGISTERS_reg[24][4]  ( .G(n2234), .D(n1921), .Q(\REGISTERS[24][4] )
         );
  DLH_X1 \REGISTERS_reg[24][3]  ( .G(n2234), .D(n1920), .Q(\REGISTERS[24][3] )
         );
  DLH_X1 \REGISTERS_reg[24][2]  ( .G(n2234), .D(n1919), .Q(\REGISTERS[24][2] )
         );
  DLH_X1 \REGISTERS_reg[24][1]  ( .G(n2234), .D(n1918), .Q(\REGISTERS[24][1] )
         );
  DLH_X1 \REGISTERS_reg[24][0]  ( .G(n2234), .D(n1917), .Q(\REGISTERS[24][0] )
         );
  DLH_X1 \REGISTERS_reg[23][31]  ( .G(n2235), .D(N3379), .Q(
        \REGISTERS[23][31] ) );
  DLH_X1 \REGISTERS_reg[23][30]  ( .G(n2235), .D(N3377), .Q(
        \REGISTERS[23][30] ) );
  DLH_X1 \REGISTERS_reg[23][29]  ( .G(n2235), .D(N3375), .Q(
        \REGISTERS[23][29] ) );
  DLH_X1 \REGISTERS_reg[23][28]  ( .G(n2235), .D(N3373), .Q(
        \REGISTERS[23][28] ) );
  DLH_X1 \REGISTERS_reg[23][27]  ( .G(n2235), .D(N3371), .Q(
        \REGISTERS[23][27] ) );
  DLH_X1 \REGISTERS_reg[23][26]  ( .G(n2235), .D(N3369), .Q(
        \REGISTERS[23][26] ) );
  DLH_X1 \REGISTERS_reg[23][25]  ( .G(n2235), .D(N3367), .Q(
        \REGISTERS[23][25] ) );
  DLH_X1 \REGISTERS_reg[23][24]  ( .G(n2235), .D(N3365), .Q(
        \REGISTERS[23][24] ) );
  DLH_X1 \REGISTERS_reg[23][23]  ( .G(n2235), .D(N3363), .Q(
        \REGISTERS[23][23] ) );
  DLH_X1 \REGISTERS_reg[23][22]  ( .G(n2235), .D(N3361), .Q(
        \REGISTERS[23][22] ) );
  DLH_X1 \REGISTERS_reg[23][21]  ( .G(n2235), .D(N3359), .Q(
        \REGISTERS[23][21] ) );
  DLH_X1 \REGISTERS_reg[23][20]  ( .G(n2235), .D(N3357), .Q(
        \REGISTERS[23][20] ) );
  DLH_X1 \REGISTERS_reg[23][19]  ( .G(n2235), .D(N3355), .Q(
        \REGISTERS[23][19] ) );
  DLH_X1 \REGISTERS_reg[23][18]  ( .G(n2236), .D(N3353), .Q(
        \REGISTERS[23][18] ) );
  DLH_X1 \REGISTERS_reg[23][17]  ( .G(n2236), .D(N3351), .Q(
        \REGISTERS[23][17] ) );
  DLH_X1 \REGISTERS_reg[23][16]  ( .G(n2236), .D(N3349), .Q(
        \REGISTERS[23][16] ) );
  DLH_X1 \REGISTERS_reg[23][15]  ( .G(n2236), .D(N3347), .Q(
        \REGISTERS[23][15] ) );
  DLH_X1 \REGISTERS_reg[23][14]  ( .G(n2236), .D(N3345), .Q(
        \REGISTERS[23][14] ) );
  DLH_X1 \REGISTERS_reg[23][13]  ( .G(n2236), .D(N3343), .Q(
        \REGISTERS[23][13] ) );
  DLH_X1 \REGISTERS_reg[23][12]  ( .G(n2236), .D(N3341), .Q(
        \REGISTERS[23][12] ) );
  DLH_X1 \REGISTERS_reg[23][11]  ( .G(n2236), .D(N3339), .Q(
        \REGISTERS[23][11] ) );
  DLH_X1 \REGISTERS_reg[23][10]  ( .G(n2236), .D(N3337), .Q(
        \REGISTERS[23][10] ) );
  DLH_X1 \REGISTERS_reg[23][9]  ( .G(n2236), .D(N3335), .Q(\REGISTERS[23][9] )
         );
  DLH_X1 \REGISTERS_reg[23][8]  ( .G(n2236), .D(N3333), .Q(\REGISTERS[23][8] )
         );
  DLH_X1 \REGISTERS_reg[23][7]  ( .G(n2236), .D(N3331), .Q(\REGISTERS[23][7] )
         );
  DLH_X1 \REGISTERS_reg[23][6]  ( .G(n2236), .D(N3329), .Q(\REGISTERS[23][6] )
         );
  DLH_X1 \REGISTERS_reg[23][5]  ( .G(n2237), .D(N3327), .Q(\REGISTERS[23][5] )
         );
  DLH_X1 \REGISTERS_reg[23][4]  ( .G(n2237), .D(N3325), .Q(\REGISTERS[23][4] )
         );
  DLH_X1 \REGISTERS_reg[23][3]  ( .G(n2237), .D(N3323), .Q(\REGISTERS[23][3] )
         );
  DLH_X1 \REGISTERS_reg[23][2]  ( .G(n2237), .D(N3321), .Q(\REGISTERS[23][2] )
         );
  DLH_X1 \REGISTERS_reg[23][1]  ( .G(n2237), .D(N3319), .Q(\REGISTERS[23][1] )
         );
  DLH_X1 \REGISTERS_reg[23][0]  ( .G(n2237), .D(N3317), .Q(\REGISTERS[23][0] )
         );
  DLH_X1 \REGISTERS_reg[22][31]  ( .G(n2238), .D(n1948), .Q(
        \REGISTERS[22][31] ) );
  DLH_X1 \REGISTERS_reg[22][30]  ( .G(n2238), .D(n1947), .Q(
        \REGISTERS[22][30] ) );
  DLH_X1 \REGISTERS_reg[22][29]  ( .G(n2238), .D(n1946), .Q(
        \REGISTERS[22][29] ) );
  DLH_X1 \REGISTERS_reg[22][28]  ( .G(n2238), .D(n1945), .Q(
        \REGISTERS[22][28] ) );
  DLH_X1 \REGISTERS_reg[22][27]  ( .G(n2238), .D(n1944), .Q(
        \REGISTERS[22][27] ) );
  DLH_X1 \REGISTERS_reg[22][26]  ( .G(n2238), .D(n1943), .Q(
        \REGISTERS[22][26] ) );
  DLH_X1 \REGISTERS_reg[22][25]  ( .G(n2238), .D(n1942), .Q(
        \REGISTERS[22][25] ) );
  DLH_X1 \REGISTERS_reg[22][24]  ( .G(n2238), .D(n1941), .Q(
        \REGISTERS[22][24] ) );
  DLH_X1 \REGISTERS_reg[22][23]  ( .G(n2238), .D(n1940), .Q(
        \REGISTERS[22][23] ) );
  DLH_X1 \REGISTERS_reg[22][22]  ( .G(n2238), .D(n1939), .Q(
        \REGISTERS[22][22] ) );
  DLH_X1 \REGISTERS_reg[22][21]  ( .G(n2238), .D(n1938), .Q(
        \REGISTERS[22][21] ) );
  DLH_X1 \REGISTERS_reg[22][20]  ( .G(n2238), .D(n1937), .Q(
        \REGISTERS[22][20] ) );
  DLH_X1 \REGISTERS_reg[22][19]  ( .G(n2238), .D(n1936), .Q(
        \REGISTERS[22][19] ) );
  DLH_X1 \REGISTERS_reg[22][18]  ( .G(n2239), .D(n1935), .Q(
        \REGISTERS[22][18] ) );
  DLH_X1 \REGISTERS_reg[22][17]  ( .G(n2239), .D(n1934), .Q(
        \REGISTERS[22][17] ) );
  DLH_X1 \REGISTERS_reg[22][16]  ( .G(n2239), .D(n1933), .Q(
        \REGISTERS[22][16] ) );
  DLH_X1 \REGISTERS_reg[22][15]  ( .G(n2239), .D(n1932), .Q(
        \REGISTERS[22][15] ) );
  DLH_X1 \REGISTERS_reg[22][14]  ( .G(n2239), .D(n1931), .Q(
        \REGISTERS[22][14] ) );
  DLH_X1 \REGISTERS_reg[22][13]  ( .G(n2239), .D(n1930), .Q(
        \REGISTERS[22][13] ) );
  DLH_X1 \REGISTERS_reg[22][12]  ( .G(n2239), .D(n1929), .Q(
        \REGISTERS[22][12] ) );
  DLH_X1 \REGISTERS_reg[22][11]  ( .G(n2239), .D(n1928), .Q(
        \REGISTERS[22][11] ) );
  DLH_X1 \REGISTERS_reg[22][10]  ( .G(n2239), .D(n1927), .Q(
        \REGISTERS[22][10] ) );
  DLH_X1 \REGISTERS_reg[22][9]  ( .G(n2239), .D(n1926), .Q(\REGISTERS[22][9] )
         );
  DLH_X1 \REGISTERS_reg[22][8]  ( .G(n2239), .D(n1925), .Q(\REGISTERS[22][8] )
         );
  DLH_X1 \REGISTERS_reg[22][7]  ( .G(n2239), .D(n1924), .Q(\REGISTERS[22][7] )
         );
  DLH_X1 \REGISTERS_reg[22][6]  ( .G(n2239), .D(n1923), .Q(\REGISTERS[22][6] )
         );
  DLH_X1 \REGISTERS_reg[22][5]  ( .G(n2240), .D(n1922), .Q(\REGISTERS[22][5] )
         );
  DLH_X1 \REGISTERS_reg[22][4]  ( .G(n2240), .D(n1921), .Q(\REGISTERS[22][4] )
         );
  DLH_X1 \REGISTERS_reg[22][3]  ( .G(n2240), .D(n1920), .Q(\REGISTERS[22][3] )
         );
  DLH_X1 \REGISTERS_reg[22][2]  ( .G(n2240), .D(n1919), .Q(\REGISTERS[22][2] )
         );
  DLH_X1 \REGISTERS_reg[22][1]  ( .G(n2240), .D(n1918), .Q(\REGISTERS[22][1] )
         );
  DLH_X1 \REGISTERS_reg[22][0]  ( .G(n2240), .D(n1917), .Q(\REGISTERS[22][0] )
         );
  DLH_X1 \REGISTERS_reg[21][31]  ( .G(n2241), .D(N3379), .Q(
        \REGISTERS[21][31] ) );
  DLH_X1 \REGISTERS_reg[21][30]  ( .G(n2241), .D(N3377), .Q(
        \REGISTERS[21][30] ) );
  DLH_X1 \REGISTERS_reg[21][29]  ( .G(n2241), .D(N3375), .Q(
        \REGISTERS[21][29] ) );
  DLH_X1 \REGISTERS_reg[21][28]  ( .G(n2241), .D(N3373), .Q(
        \REGISTERS[21][28] ) );
  DLH_X1 \REGISTERS_reg[21][27]  ( .G(n2241), .D(N3371), .Q(
        \REGISTERS[21][27] ) );
  DLH_X1 \REGISTERS_reg[21][26]  ( .G(n2241), .D(N3369), .Q(
        \REGISTERS[21][26] ) );
  DLH_X1 \REGISTERS_reg[21][25]  ( .G(n2241), .D(N3367), .Q(
        \REGISTERS[21][25] ) );
  DLH_X1 \REGISTERS_reg[21][24]  ( .G(n2241), .D(N3365), .Q(
        \REGISTERS[21][24] ) );
  DLH_X1 \REGISTERS_reg[21][23]  ( .G(n2241), .D(N3363), .Q(
        \REGISTERS[21][23] ) );
  DLH_X1 \REGISTERS_reg[21][22]  ( .G(n2241), .D(N3361), .Q(
        \REGISTERS[21][22] ) );
  DLH_X1 \REGISTERS_reg[21][21]  ( .G(n2241), .D(N3359), .Q(
        \REGISTERS[21][21] ) );
  DLH_X1 \REGISTERS_reg[21][20]  ( .G(n2241), .D(N3357), .Q(
        \REGISTERS[21][20] ) );
  DLH_X1 \REGISTERS_reg[21][19]  ( .G(n2241), .D(N3355), .Q(
        \REGISTERS[21][19] ) );
  DLH_X1 \REGISTERS_reg[21][18]  ( .G(n2242), .D(N3353), .Q(
        \REGISTERS[21][18] ) );
  DLH_X1 \REGISTERS_reg[21][17]  ( .G(n2242), .D(N3351), .Q(
        \REGISTERS[21][17] ) );
  DLH_X1 \REGISTERS_reg[21][16]  ( .G(n2242), .D(N3349), .Q(
        \REGISTERS[21][16] ) );
  DLH_X1 \REGISTERS_reg[21][15]  ( .G(n2242), .D(N3347), .Q(
        \REGISTERS[21][15] ) );
  DLH_X1 \REGISTERS_reg[21][14]  ( .G(n2242), .D(N3345), .Q(
        \REGISTERS[21][14] ) );
  DLH_X1 \REGISTERS_reg[21][13]  ( .G(n2242), .D(N3343), .Q(
        \REGISTERS[21][13] ) );
  DLH_X1 \REGISTERS_reg[21][12]  ( .G(n2242), .D(N3341), .Q(
        \REGISTERS[21][12] ) );
  DLH_X1 \REGISTERS_reg[21][11]  ( .G(n2242), .D(N3339), .Q(
        \REGISTERS[21][11] ) );
  DLH_X1 \REGISTERS_reg[21][10]  ( .G(n2242), .D(N3337), .Q(
        \REGISTERS[21][10] ) );
  DLH_X1 \REGISTERS_reg[21][9]  ( .G(n2242), .D(N3335), .Q(\REGISTERS[21][9] )
         );
  DLH_X1 \REGISTERS_reg[21][8]  ( .G(n2242), .D(N3333), .Q(\REGISTERS[21][8] )
         );
  DLH_X1 \REGISTERS_reg[21][7]  ( .G(n2242), .D(N3331), .Q(\REGISTERS[21][7] )
         );
  DLH_X1 \REGISTERS_reg[21][6]  ( .G(n2242), .D(N3329), .Q(\REGISTERS[21][6] )
         );
  DLH_X1 \REGISTERS_reg[21][5]  ( .G(n2243), .D(N3327), .Q(\REGISTERS[21][5] )
         );
  DLH_X1 \REGISTERS_reg[21][4]  ( .G(n2243), .D(N3325), .Q(\REGISTERS[21][4] )
         );
  DLH_X1 \REGISTERS_reg[21][3]  ( .G(n2243), .D(N3323), .Q(\REGISTERS[21][3] )
         );
  DLH_X1 \REGISTERS_reg[21][2]  ( .G(n2243), .D(N3321), .Q(\REGISTERS[21][2] )
         );
  DLH_X1 \REGISTERS_reg[21][1]  ( .G(n2243), .D(N3319), .Q(\REGISTERS[21][1] )
         );
  DLH_X1 \REGISTERS_reg[21][0]  ( .G(n2243), .D(N3317), .Q(\REGISTERS[21][0] )
         );
  DLH_X1 \REGISTERS_reg[20][31]  ( .G(n2244), .D(n1948), .Q(
        \REGISTERS[20][31] ) );
  DLH_X1 \REGISTERS_reg[20][30]  ( .G(n2244), .D(n1947), .Q(
        \REGISTERS[20][30] ) );
  DLH_X1 \REGISTERS_reg[20][29]  ( .G(n2244), .D(n1946), .Q(
        \REGISTERS[20][29] ) );
  DLH_X1 \REGISTERS_reg[20][28]  ( .G(n2244), .D(n1945), .Q(
        \REGISTERS[20][28] ) );
  DLH_X1 \REGISTERS_reg[20][27]  ( .G(n2244), .D(n1944), .Q(
        \REGISTERS[20][27] ) );
  DLH_X1 \REGISTERS_reg[20][26]  ( .G(n2244), .D(n1943), .Q(
        \REGISTERS[20][26] ) );
  DLH_X1 \REGISTERS_reg[20][25]  ( .G(n2244), .D(n1942), .Q(
        \REGISTERS[20][25] ) );
  DLH_X1 \REGISTERS_reg[20][24]  ( .G(n2244), .D(n1941), .Q(
        \REGISTERS[20][24] ) );
  DLH_X1 \REGISTERS_reg[20][23]  ( .G(n2244), .D(n1940), .Q(
        \REGISTERS[20][23] ) );
  DLH_X1 \REGISTERS_reg[20][22]  ( .G(n2244), .D(n1939), .Q(
        \REGISTERS[20][22] ) );
  DLH_X1 \REGISTERS_reg[20][21]  ( .G(n2244), .D(n1938), .Q(
        \REGISTERS[20][21] ) );
  DLH_X1 \REGISTERS_reg[20][20]  ( .G(n2244), .D(n1937), .Q(
        \REGISTERS[20][20] ) );
  DLH_X1 \REGISTERS_reg[20][19]  ( .G(n2244), .D(n1936), .Q(
        \REGISTERS[20][19] ) );
  DLH_X1 \REGISTERS_reg[20][18]  ( .G(n2245), .D(n1935), .Q(
        \REGISTERS[20][18] ) );
  DLH_X1 \REGISTERS_reg[20][17]  ( .G(n2245), .D(n1934), .Q(
        \REGISTERS[20][17] ) );
  DLH_X1 \REGISTERS_reg[20][16]  ( .G(n2245), .D(n1933), .Q(
        \REGISTERS[20][16] ) );
  DLH_X1 \REGISTERS_reg[20][15]  ( .G(n2245), .D(n1932), .Q(
        \REGISTERS[20][15] ) );
  DLH_X1 \REGISTERS_reg[20][14]  ( .G(n2245), .D(n1931), .Q(
        \REGISTERS[20][14] ) );
  DLH_X1 \REGISTERS_reg[20][13]  ( .G(n2245), .D(n1930), .Q(
        \REGISTERS[20][13] ) );
  DLH_X1 \REGISTERS_reg[20][12]  ( .G(n2245), .D(n1929), .Q(
        \REGISTERS[20][12] ) );
  DLH_X1 \REGISTERS_reg[20][11]  ( .G(n2245), .D(n1928), .Q(
        \REGISTERS[20][11] ) );
  DLH_X1 \REGISTERS_reg[20][10]  ( .G(n2245), .D(n1927), .Q(
        \REGISTERS[20][10] ) );
  DLH_X1 \REGISTERS_reg[20][9]  ( .G(n2245), .D(n1926), .Q(\REGISTERS[20][9] )
         );
  DLH_X1 \REGISTERS_reg[20][8]  ( .G(n2245), .D(n1925), .Q(\REGISTERS[20][8] )
         );
  DLH_X1 \REGISTERS_reg[20][7]  ( .G(n2245), .D(n1924), .Q(\REGISTERS[20][7] )
         );
  DLH_X1 \REGISTERS_reg[20][6]  ( .G(n2245), .D(n1923), .Q(\REGISTERS[20][6] )
         );
  DLH_X1 \REGISTERS_reg[20][5]  ( .G(n2246), .D(n1922), .Q(\REGISTERS[20][5] )
         );
  DLH_X1 \REGISTERS_reg[20][4]  ( .G(n2246), .D(n1921), .Q(\REGISTERS[20][4] )
         );
  DLH_X1 \REGISTERS_reg[20][3]  ( .G(n2246), .D(n1920), .Q(\REGISTERS[20][3] )
         );
  DLH_X1 \REGISTERS_reg[20][2]  ( .G(n2246), .D(n1919), .Q(\REGISTERS[20][2] )
         );
  DLH_X1 \REGISTERS_reg[20][1]  ( .G(n2246), .D(n1918), .Q(\REGISTERS[20][1] )
         );
  DLH_X1 \REGISTERS_reg[20][0]  ( .G(n2246), .D(n1917), .Q(\REGISTERS[20][0] )
         );
  DLH_X1 \REGISTERS_reg[19][31]  ( .G(n2247), .D(N3379), .Q(
        \REGISTERS[19][31] ) );
  DLH_X1 \REGISTERS_reg[19][30]  ( .G(n2247), .D(N3377), .Q(
        \REGISTERS[19][30] ) );
  DLH_X1 \REGISTERS_reg[19][29]  ( .G(n2247), .D(N3375), .Q(
        \REGISTERS[19][29] ) );
  DLH_X1 \REGISTERS_reg[19][28]  ( .G(n2247), .D(N3373), .Q(
        \REGISTERS[19][28] ) );
  DLH_X1 \REGISTERS_reg[19][27]  ( .G(n2247), .D(N3371), .Q(
        \REGISTERS[19][27] ) );
  DLH_X1 \REGISTERS_reg[19][26]  ( .G(n2247), .D(N3369), .Q(
        \REGISTERS[19][26] ) );
  DLH_X1 \REGISTERS_reg[19][25]  ( .G(n2247), .D(N3367), .Q(
        \REGISTERS[19][25] ) );
  DLH_X1 \REGISTERS_reg[19][24]  ( .G(n2247), .D(N3365), .Q(
        \REGISTERS[19][24] ) );
  DLH_X1 \REGISTERS_reg[19][23]  ( .G(n2247), .D(N3363), .Q(
        \REGISTERS[19][23] ) );
  DLH_X1 \REGISTERS_reg[19][22]  ( .G(n2247), .D(N3361), .Q(
        \REGISTERS[19][22] ) );
  DLH_X1 \REGISTERS_reg[19][21]  ( .G(n2247), .D(N3359), .Q(
        \REGISTERS[19][21] ) );
  DLH_X1 \REGISTERS_reg[19][20]  ( .G(n2247), .D(N3357), .Q(
        \REGISTERS[19][20] ) );
  DLH_X1 \REGISTERS_reg[19][19]  ( .G(n2247), .D(N3355), .Q(
        \REGISTERS[19][19] ) );
  DLH_X1 \REGISTERS_reg[19][18]  ( .G(n2248), .D(N3353), .Q(
        \REGISTERS[19][18] ) );
  DLH_X1 \REGISTERS_reg[19][17]  ( .G(n2248), .D(N3351), .Q(
        \REGISTERS[19][17] ) );
  DLH_X1 \REGISTERS_reg[19][16]  ( .G(n2248), .D(N3349), .Q(
        \REGISTERS[19][16] ) );
  DLH_X1 \REGISTERS_reg[19][15]  ( .G(n2248), .D(N3347), .Q(
        \REGISTERS[19][15] ) );
  DLH_X1 \REGISTERS_reg[19][14]  ( .G(n2248), .D(N3345), .Q(
        \REGISTERS[19][14] ) );
  DLH_X1 \REGISTERS_reg[19][13]  ( .G(n2248), .D(N3343), .Q(
        \REGISTERS[19][13] ) );
  DLH_X1 \REGISTERS_reg[19][12]  ( .G(n2248), .D(N3341), .Q(
        \REGISTERS[19][12] ) );
  DLH_X1 \REGISTERS_reg[19][11]  ( .G(n2248), .D(N3339), .Q(
        \REGISTERS[19][11] ) );
  DLH_X1 \REGISTERS_reg[19][10]  ( .G(n2248), .D(N3337), .Q(
        \REGISTERS[19][10] ) );
  DLH_X1 \REGISTERS_reg[19][9]  ( .G(n2248), .D(N3335), .Q(\REGISTERS[19][9] )
         );
  DLH_X1 \REGISTERS_reg[19][8]  ( .G(n2248), .D(N3333), .Q(\REGISTERS[19][8] )
         );
  DLH_X1 \REGISTERS_reg[19][7]  ( .G(n2248), .D(N3331), .Q(\REGISTERS[19][7] )
         );
  DLH_X1 \REGISTERS_reg[19][6]  ( .G(n2248), .D(N3329), .Q(\REGISTERS[19][6] )
         );
  DLH_X1 \REGISTERS_reg[19][5]  ( .G(n2249), .D(N3327), .Q(\REGISTERS[19][5] )
         );
  DLH_X1 \REGISTERS_reg[19][4]  ( .G(n2249), .D(N3325), .Q(\REGISTERS[19][4] )
         );
  DLH_X1 \REGISTERS_reg[19][3]  ( .G(n2249), .D(N3323), .Q(\REGISTERS[19][3] )
         );
  DLH_X1 \REGISTERS_reg[19][2]  ( .G(n2249), .D(N3321), .Q(\REGISTERS[19][2] )
         );
  DLH_X1 \REGISTERS_reg[19][1]  ( .G(n2249), .D(N3319), .Q(\REGISTERS[19][1] )
         );
  DLH_X1 \REGISTERS_reg[19][0]  ( .G(n2249), .D(N3317), .Q(\REGISTERS[19][0] )
         );
  DLH_X1 \REGISTERS_reg[18][31]  ( .G(n2250), .D(n1948), .Q(
        \REGISTERS[18][31] ) );
  DLH_X1 \REGISTERS_reg[18][30]  ( .G(n2250), .D(n1947), .Q(
        \REGISTERS[18][30] ) );
  DLH_X1 \REGISTERS_reg[18][29]  ( .G(n2250), .D(n1946), .Q(
        \REGISTERS[18][29] ) );
  DLH_X1 \REGISTERS_reg[18][28]  ( .G(n2250), .D(n1945), .Q(
        \REGISTERS[18][28] ) );
  DLH_X1 \REGISTERS_reg[18][27]  ( .G(n2250), .D(n1944), .Q(
        \REGISTERS[18][27] ) );
  DLH_X1 \REGISTERS_reg[18][26]  ( .G(n2250), .D(n1943), .Q(
        \REGISTERS[18][26] ) );
  DLH_X1 \REGISTERS_reg[18][25]  ( .G(n2250), .D(n1942), .Q(
        \REGISTERS[18][25] ) );
  DLH_X1 \REGISTERS_reg[18][24]  ( .G(n2250), .D(n1941), .Q(
        \REGISTERS[18][24] ) );
  DLH_X1 \REGISTERS_reg[18][23]  ( .G(n2250), .D(n1940), .Q(
        \REGISTERS[18][23] ) );
  DLH_X1 \REGISTERS_reg[18][22]  ( .G(n2250), .D(n1939), .Q(
        \REGISTERS[18][22] ) );
  DLH_X1 \REGISTERS_reg[18][21]  ( .G(n2250), .D(n1938), .Q(
        \REGISTERS[18][21] ) );
  DLH_X1 \REGISTERS_reg[18][20]  ( .G(n2250), .D(n1937), .Q(
        \REGISTERS[18][20] ) );
  DLH_X1 \REGISTERS_reg[18][19]  ( .G(n2250), .D(n1936), .Q(
        \REGISTERS[18][19] ) );
  DLH_X1 \REGISTERS_reg[18][18]  ( .G(n2251), .D(n1935), .Q(
        \REGISTERS[18][18] ) );
  DLH_X1 \REGISTERS_reg[18][17]  ( .G(n2251), .D(n1934), .Q(
        \REGISTERS[18][17] ) );
  DLH_X1 \REGISTERS_reg[18][16]  ( .G(n2251), .D(n1933), .Q(
        \REGISTERS[18][16] ) );
  DLH_X1 \REGISTERS_reg[18][15]  ( .G(n2251), .D(n1932), .Q(
        \REGISTERS[18][15] ) );
  DLH_X1 \REGISTERS_reg[18][14]  ( .G(n2251), .D(n1931), .Q(
        \REGISTERS[18][14] ) );
  DLH_X1 \REGISTERS_reg[18][13]  ( .G(n2251), .D(n1930), .Q(
        \REGISTERS[18][13] ) );
  DLH_X1 \REGISTERS_reg[18][12]  ( .G(n2251), .D(n1929), .Q(
        \REGISTERS[18][12] ) );
  DLH_X1 \REGISTERS_reg[18][11]  ( .G(n2251), .D(n1928), .Q(
        \REGISTERS[18][11] ) );
  DLH_X1 \REGISTERS_reg[18][10]  ( .G(n2251), .D(n1927), .Q(
        \REGISTERS[18][10] ) );
  DLH_X1 \REGISTERS_reg[18][9]  ( .G(n2251), .D(n1926), .Q(\REGISTERS[18][9] )
         );
  DLH_X1 \REGISTERS_reg[18][8]  ( .G(n2251), .D(n1925), .Q(\REGISTERS[18][8] )
         );
  DLH_X1 \REGISTERS_reg[18][7]  ( .G(n2251), .D(n1924), .Q(\REGISTERS[18][7] )
         );
  DLH_X1 \REGISTERS_reg[18][6]  ( .G(n2251), .D(n1923), .Q(\REGISTERS[18][6] )
         );
  DLH_X1 \REGISTERS_reg[18][5]  ( .G(n2252), .D(n1922), .Q(\REGISTERS[18][5] )
         );
  DLH_X1 \REGISTERS_reg[18][4]  ( .G(n2252), .D(n1921), .Q(\REGISTERS[18][4] )
         );
  DLH_X1 \REGISTERS_reg[18][3]  ( .G(n2252), .D(n1920), .Q(\REGISTERS[18][3] )
         );
  DLH_X1 \REGISTERS_reg[18][2]  ( .G(n2252), .D(n1919), .Q(\REGISTERS[18][2] )
         );
  DLH_X1 \REGISTERS_reg[18][1]  ( .G(n2252), .D(n1918), .Q(\REGISTERS[18][1] )
         );
  DLH_X1 \REGISTERS_reg[18][0]  ( .G(n2252), .D(n1917), .Q(\REGISTERS[18][0] )
         );
  DLH_X1 \REGISTERS_reg[17][31]  ( .G(n2253), .D(N3379), .Q(
        \REGISTERS[17][31] ) );
  DLH_X1 \REGISTERS_reg[17][30]  ( .G(n2253), .D(N3377), .Q(
        \REGISTERS[17][30] ) );
  DLH_X1 \REGISTERS_reg[17][29]  ( .G(n2253), .D(N3375), .Q(
        \REGISTERS[17][29] ) );
  DLH_X1 \REGISTERS_reg[17][28]  ( .G(n2253), .D(N3373), .Q(
        \REGISTERS[17][28] ) );
  DLH_X1 \REGISTERS_reg[17][27]  ( .G(n2253), .D(N3371), .Q(
        \REGISTERS[17][27] ) );
  DLH_X1 \REGISTERS_reg[17][26]  ( .G(n2253), .D(N3369), .Q(
        \REGISTERS[17][26] ) );
  DLH_X1 \REGISTERS_reg[17][25]  ( .G(n2253), .D(N3367), .Q(
        \REGISTERS[17][25] ) );
  DLH_X1 \REGISTERS_reg[17][24]  ( .G(n2253), .D(N3365), .Q(
        \REGISTERS[17][24] ) );
  DLH_X1 \REGISTERS_reg[17][23]  ( .G(n2253), .D(N3363), .Q(
        \REGISTERS[17][23] ) );
  DLH_X1 \REGISTERS_reg[17][22]  ( .G(n2253), .D(N3361), .Q(
        \REGISTERS[17][22] ) );
  DLH_X1 \REGISTERS_reg[17][21]  ( .G(n2253), .D(N3359), .Q(
        \REGISTERS[17][21] ) );
  DLH_X1 \REGISTERS_reg[17][20]  ( .G(n2253), .D(N3357), .Q(
        \REGISTERS[17][20] ) );
  DLH_X1 \REGISTERS_reg[17][19]  ( .G(n2253), .D(N3355), .Q(
        \REGISTERS[17][19] ) );
  DLH_X1 \REGISTERS_reg[17][18]  ( .G(n2254), .D(N3353), .Q(
        \REGISTERS[17][18] ) );
  DLH_X1 \REGISTERS_reg[17][17]  ( .G(n2254), .D(N3351), .Q(
        \REGISTERS[17][17] ) );
  DLH_X1 \REGISTERS_reg[17][16]  ( .G(n2254), .D(N3349), .Q(
        \REGISTERS[17][16] ) );
  DLH_X1 \REGISTERS_reg[17][15]  ( .G(n2254), .D(N3347), .Q(
        \REGISTERS[17][15] ) );
  DLH_X1 \REGISTERS_reg[17][14]  ( .G(n2254), .D(N3345), .Q(
        \REGISTERS[17][14] ) );
  DLH_X1 \REGISTERS_reg[17][13]  ( .G(n2254), .D(N3343), .Q(
        \REGISTERS[17][13] ) );
  DLH_X1 \REGISTERS_reg[17][12]  ( .G(n2254), .D(N3341), .Q(
        \REGISTERS[17][12] ) );
  DLH_X1 \REGISTERS_reg[17][11]  ( .G(n2254), .D(N3339), .Q(
        \REGISTERS[17][11] ) );
  DLH_X1 \REGISTERS_reg[17][10]  ( .G(n2254), .D(N3337), .Q(
        \REGISTERS[17][10] ) );
  DLH_X1 \REGISTERS_reg[17][9]  ( .G(n2254), .D(N3335), .Q(\REGISTERS[17][9] )
         );
  DLH_X1 \REGISTERS_reg[17][8]  ( .G(n2254), .D(N3333), .Q(\REGISTERS[17][8] )
         );
  DLH_X1 \REGISTERS_reg[17][7]  ( .G(n2254), .D(N3331), .Q(\REGISTERS[17][7] )
         );
  DLH_X1 \REGISTERS_reg[17][6]  ( .G(n2254), .D(N3329), .Q(\REGISTERS[17][6] )
         );
  DLH_X1 \REGISTERS_reg[17][5]  ( .G(n2255), .D(N3327), .Q(\REGISTERS[17][5] )
         );
  DLH_X1 \REGISTERS_reg[17][4]  ( .G(n2255), .D(N3325), .Q(\REGISTERS[17][4] )
         );
  DLH_X1 \REGISTERS_reg[17][3]  ( .G(n2255), .D(N3323), .Q(\REGISTERS[17][3] )
         );
  DLH_X1 \REGISTERS_reg[17][2]  ( .G(n2255), .D(N3321), .Q(\REGISTERS[17][2] )
         );
  DLH_X1 \REGISTERS_reg[17][1]  ( .G(n2255), .D(N3319), .Q(\REGISTERS[17][1] )
         );
  DLH_X1 \REGISTERS_reg[17][0]  ( .G(n2255), .D(N3317), .Q(\REGISTERS[17][0] )
         );
  DLH_X1 \REGISTERS_reg[16][31]  ( .G(n2256), .D(n1948), .Q(
        \REGISTERS[16][31] ) );
  DLH_X1 \REGISTERS_reg[16][30]  ( .G(n2256), .D(n1947), .Q(
        \REGISTERS[16][30] ) );
  DLH_X1 \REGISTERS_reg[16][29]  ( .G(n2256), .D(n1946), .Q(
        \REGISTERS[16][29] ) );
  DLH_X1 \REGISTERS_reg[16][28]  ( .G(n2256), .D(n1945), .Q(
        \REGISTERS[16][28] ) );
  DLH_X1 \REGISTERS_reg[16][27]  ( .G(n2256), .D(n1944), .Q(
        \REGISTERS[16][27] ) );
  DLH_X1 \REGISTERS_reg[16][26]  ( .G(n2256), .D(n1943), .Q(
        \REGISTERS[16][26] ) );
  DLH_X1 \REGISTERS_reg[16][25]  ( .G(n2256), .D(n1942), .Q(
        \REGISTERS[16][25] ) );
  DLH_X1 \REGISTERS_reg[16][24]  ( .G(n2256), .D(n1941), .Q(
        \REGISTERS[16][24] ) );
  DLH_X1 \REGISTERS_reg[16][23]  ( .G(n2256), .D(n1940), .Q(
        \REGISTERS[16][23] ) );
  DLH_X1 \REGISTERS_reg[16][22]  ( .G(n2256), .D(n1939), .Q(
        \REGISTERS[16][22] ) );
  DLH_X1 \REGISTERS_reg[16][21]  ( .G(n2256), .D(n1938), .Q(
        \REGISTERS[16][21] ) );
  DLH_X1 \REGISTERS_reg[16][20]  ( .G(n2256), .D(n1937), .Q(
        \REGISTERS[16][20] ) );
  DLH_X1 \REGISTERS_reg[16][19]  ( .G(n2256), .D(n1936), .Q(
        \REGISTERS[16][19] ) );
  DLH_X1 \REGISTERS_reg[16][18]  ( .G(n2257), .D(n1935), .Q(
        \REGISTERS[16][18] ) );
  DLH_X1 \REGISTERS_reg[16][17]  ( .G(n2257), .D(n1934), .Q(
        \REGISTERS[16][17] ) );
  DLH_X1 \REGISTERS_reg[16][16]  ( .G(n2257), .D(n1933), .Q(
        \REGISTERS[16][16] ) );
  DLH_X1 \REGISTERS_reg[16][15]  ( .G(n2257), .D(n1932), .Q(
        \REGISTERS[16][15] ) );
  DLH_X1 \REGISTERS_reg[16][14]  ( .G(n2257), .D(n1931), .Q(
        \REGISTERS[16][14] ) );
  DLH_X1 \REGISTERS_reg[16][13]  ( .G(n2257), .D(n1930), .Q(
        \REGISTERS[16][13] ) );
  DLH_X1 \REGISTERS_reg[16][12]  ( .G(n2257), .D(n1929), .Q(
        \REGISTERS[16][12] ) );
  DLH_X1 \REGISTERS_reg[16][11]  ( .G(n2257), .D(n1928), .Q(
        \REGISTERS[16][11] ) );
  DLH_X1 \REGISTERS_reg[16][10]  ( .G(n2257), .D(n1927), .Q(
        \REGISTERS[16][10] ) );
  DLH_X1 \REGISTERS_reg[16][9]  ( .G(n2257), .D(n1926), .Q(\REGISTERS[16][9] )
         );
  DLH_X1 \REGISTERS_reg[16][8]  ( .G(n2257), .D(n1925), .Q(\REGISTERS[16][8] )
         );
  DLH_X1 \REGISTERS_reg[16][7]  ( .G(n2257), .D(n1924), .Q(\REGISTERS[16][7] )
         );
  DLH_X1 \REGISTERS_reg[16][6]  ( .G(n2257), .D(n1923), .Q(\REGISTERS[16][6] )
         );
  DLH_X1 \REGISTERS_reg[16][5]  ( .G(n2258), .D(n1922), .Q(\REGISTERS[16][5] )
         );
  DLH_X1 \REGISTERS_reg[16][4]  ( .G(n2258), .D(n1921), .Q(\REGISTERS[16][4] )
         );
  DLH_X1 \REGISTERS_reg[16][3]  ( .G(n2258), .D(n1920), .Q(\REGISTERS[16][3] )
         );
  DLH_X1 \REGISTERS_reg[16][2]  ( .G(n2258), .D(n1919), .Q(\REGISTERS[16][2] )
         );
  DLH_X1 \REGISTERS_reg[16][1]  ( .G(n2258), .D(n1918), .Q(\REGISTERS[16][1] )
         );
  DLH_X1 \REGISTERS_reg[16][0]  ( .G(n2258), .D(n1917), .Q(\REGISTERS[16][0] )
         );
  DLH_X1 \REGISTERS_reg[15][31]  ( .G(n2259), .D(N3379), .Q(
        \REGISTERS[15][31] ) );
  DLH_X1 \REGISTERS_reg[15][30]  ( .G(n2259), .D(N3377), .Q(
        \REGISTERS[15][30] ) );
  DLH_X1 \REGISTERS_reg[15][29]  ( .G(n2259), .D(N3375), .Q(
        \REGISTERS[15][29] ) );
  DLH_X1 \REGISTERS_reg[15][28]  ( .G(n2259), .D(N3373), .Q(
        \REGISTERS[15][28] ) );
  DLH_X1 \REGISTERS_reg[15][27]  ( .G(n2259), .D(N3371), .Q(
        \REGISTERS[15][27] ) );
  DLH_X1 \REGISTERS_reg[15][26]  ( .G(n2259), .D(N3369), .Q(
        \REGISTERS[15][26] ) );
  DLH_X1 \REGISTERS_reg[15][25]  ( .G(n2259), .D(N3367), .Q(
        \REGISTERS[15][25] ) );
  DLH_X1 \REGISTERS_reg[15][24]  ( .G(n2259), .D(N3365), .Q(
        \REGISTERS[15][24] ) );
  DLH_X1 \REGISTERS_reg[15][23]  ( .G(n2259), .D(N3363), .Q(
        \REGISTERS[15][23] ) );
  DLH_X1 \REGISTERS_reg[15][22]  ( .G(n2259), .D(N3361), .Q(
        \REGISTERS[15][22] ) );
  DLH_X1 \REGISTERS_reg[15][21]  ( .G(n2259), .D(N3359), .Q(
        \REGISTERS[15][21] ) );
  DLH_X1 \REGISTERS_reg[15][20]  ( .G(n2259), .D(N3357), .Q(
        \REGISTERS[15][20] ) );
  DLH_X1 \REGISTERS_reg[15][19]  ( .G(n2259), .D(N3355), .Q(
        \REGISTERS[15][19] ) );
  DLH_X1 \REGISTERS_reg[15][18]  ( .G(n2260), .D(N3353), .Q(
        \REGISTERS[15][18] ) );
  DLH_X1 \REGISTERS_reg[15][17]  ( .G(n2260), .D(N3351), .Q(
        \REGISTERS[15][17] ) );
  DLH_X1 \REGISTERS_reg[15][16]  ( .G(n2260), .D(N3349), .Q(
        \REGISTERS[15][16] ) );
  DLH_X1 \REGISTERS_reg[15][15]  ( .G(n2260), .D(N3347), .Q(
        \REGISTERS[15][15] ) );
  DLH_X1 \REGISTERS_reg[15][14]  ( .G(n2260), .D(N3345), .Q(
        \REGISTERS[15][14] ) );
  DLH_X1 \REGISTERS_reg[15][13]  ( .G(n2260), .D(N3343), .Q(
        \REGISTERS[15][13] ) );
  DLH_X1 \REGISTERS_reg[15][12]  ( .G(n2260), .D(N3341), .Q(
        \REGISTERS[15][12] ) );
  DLH_X1 \REGISTERS_reg[15][11]  ( .G(n2260), .D(N3339), .Q(
        \REGISTERS[15][11] ) );
  DLH_X1 \REGISTERS_reg[15][10]  ( .G(n2260), .D(N3337), .Q(
        \REGISTERS[15][10] ) );
  DLH_X1 \REGISTERS_reg[15][9]  ( .G(n2260), .D(N3335), .Q(\REGISTERS[15][9] )
         );
  DLH_X1 \REGISTERS_reg[15][8]  ( .G(n2260), .D(N3333), .Q(\REGISTERS[15][8] )
         );
  DLH_X1 \REGISTERS_reg[15][7]  ( .G(n2260), .D(N3331), .Q(\REGISTERS[15][7] )
         );
  DLH_X1 \REGISTERS_reg[15][6]  ( .G(n2260), .D(N3329), .Q(\REGISTERS[15][6] )
         );
  DLH_X1 \REGISTERS_reg[15][5]  ( .G(n2261), .D(N3327), .Q(\REGISTERS[15][5] )
         );
  DLH_X1 \REGISTERS_reg[15][4]  ( .G(n2261), .D(N3325), .Q(\REGISTERS[15][4] )
         );
  DLH_X1 \REGISTERS_reg[15][3]  ( .G(n2261), .D(N3323), .Q(\REGISTERS[15][3] )
         );
  DLH_X1 \REGISTERS_reg[15][2]  ( .G(n2261), .D(N3321), .Q(\REGISTERS[15][2] )
         );
  DLH_X1 \REGISTERS_reg[15][1]  ( .G(n2261), .D(N3319), .Q(\REGISTERS[15][1] )
         );
  DLH_X1 \REGISTERS_reg[15][0]  ( .G(n2261), .D(N3317), .Q(\REGISTERS[15][0] )
         );
  DLH_X1 \REGISTERS_reg[14][31]  ( .G(n2262), .D(n1948), .Q(
        \REGISTERS[14][31] ) );
  DLH_X1 \REGISTERS_reg[14][30]  ( .G(n2262), .D(n1947), .Q(
        \REGISTERS[14][30] ) );
  DLH_X1 \REGISTERS_reg[14][29]  ( .G(n2262), .D(n1946), .Q(
        \REGISTERS[14][29] ) );
  DLH_X1 \REGISTERS_reg[14][28]  ( .G(n2262), .D(n1945), .Q(
        \REGISTERS[14][28] ) );
  DLH_X1 \REGISTERS_reg[14][27]  ( .G(n2262), .D(n1944), .Q(
        \REGISTERS[14][27] ) );
  DLH_X1 \REGISTERS_reg[14][26]  ( .G(n2262), .D(n1943), .Q(
        \REGISTERS[14][26] ) );
  DLH_X1 \REGISTERS_reg[14][25]  ( .G(n2262), .D(n1942), .Q(
        \REGISTERS[14][25] ) );
  DLH_X1 \REGISTERS_reg[14][24]  ( .G(n2262), .D(n1941), .Q(
        \REGISTERS[14][24] ) );
  DLH_X1 \REGISTERS_reg[14][23]  ( .G(n2262), .D(n1940), .Q(
        \REGISTERS[14][23] ) );
  DLH_X1 \REGISTERS_reg[14][22]  ( .G(n2262), .D(n1939), .Q(
        \REGISTERS[14][22] ) );
  DLH_X1 \REGISTERS_reg[14][21]  ( .G(n2262), .D(n1938), .Q(
        \REGISTERS[14][21] ) );
  DLH_X1 \REGISTERS_reg[14][20]  ( .G(n2262), .D(n1937), .Q(
        \REGISTERS[14][20] ) );
  DLH_X1 \REGISTERS_reg[14][19]  ( .G(n2262), .D(n1936), .Q(
        \REGISTERS[14][19] ) );
  DLH_X1 \REGISTERS_reg[14][18]  ( .G(n2263), .D(n1935), .Q(
        \REGISTERS[14][18] ) );
  DLH_X1 \REGISTERS_reg[14][17]  ( .G(n2263), .D(n1934), .Q(
        \REGISTERS[14][17] ) );
  DLH_X1 \REGISTERS_reg[14][16]  ( .G(n2263), .D(n1933), .Q(
        \REGISTERS[14][16] ) );
  DLH_X1 \REGISTERS_reg[14][15]  ( .G(n2263), .D(n1932), .Q(
        \REGISTERS[14][15] ) );
  DLH_X1 \REGISTERS_reg[14][14]  ( .G(n2263), .D(n1931), .Q(
        \REGISTERS[14][14] ) );
  DLH_X1 \REGISTERS_reg[14][13]  ( .G(n2263), .D(n1930), .Q(
        \REGISTERS[14][13] ) );
  DLH_X1 \REGISTERS_reg[14][12]  ( .G(n2263), .D(n1929), .Q(
        \REGISTERS[14][12] ) );
  DLH_X1 \REGISTERS_reg[14][11]  ( .G(n2263), .D(n1928), .Q(
        \REGISTERS[14][11] ) );
  DLH_X1 \REGISTERS_reg[14][10]  ( .G(n2263), .D(n1927), .Q(
        \REGISTERS[14][10] ) );
  DLH_X1 \REGISTERS_reg[14][9]  ( .G(n2263), .D(n1926), .Q(\REGISTERS[14][9] )
         );
  DLH_X1 \REGISTERS_reg[14][8]  ( .G(n2263), .D(n1925), .Q(\REGISTERS[14][8] )
         );
  DLH_X1 \REGISTERS_reg[14][7]  ( .G(n2263), .D(n1924), .Q(\REGISTERS[14][7] )
         );
  DLH_X1 \REGISTERS_reg[14][6]  ( .G(n2263), .D(n1923), .Q(\REGISTERS[14][6] )
         );
  DLH_X1 \REGISTERS_reg[14][5]  ( .G(n2264), .D(n1922), .Q(\REGISTERS[14][5] )
         );
  DLH_X1 \REGISTERS_reg[14][4]  ( .G(n2264), .D(n1921), .Q(\REGISTERS[14][4] )
         );
  DLH_X1 \REGISTERS_reg[14][3]  ( .G(n2264), .D(n1920), .Q(\REGISTERS[14][3] )
         );
  DLH_X1 \REGISTERS_reg[14][2]  ( .G(n2264), .D(n1919), .Q(\REGISTERS[14][2] )
         );
  DLH_X1 \REGISTERS_reg[14][1]  ( .G(n2264), .D(n1918), .Q(\REGISTERS[14][1] )
         );
  DLH_X1 \REGISTERS_reg[14][0]  ( .G(n2264), .D(n1917), .Q(\REGISTERS[14][0] )
         );
  DLH_X1 \REGISTERS_reg[13][31]  ( .G(n2265), .D(N3379), .Q(
        \REGISTERS[13][31] ) );
  DLH_X1 \REGISTERS_reg[13][30]  ( .G(n2265), .D(N3377), .Q(
        \REGISTERS[13][30] ) );
  DLH_X1 \REGISTERS_reg[13][29]  ( .G(n2265), .D(N3375), .Q(
        \REGISTERS[13][29] ) );
  DLH_X1 \REGISTERS_reg[13][28]  ( .G(n2265), .D(N3373), .Q(
        \REGISTERS[13][28] ) );
  DLH_X1 \REGISTERS_reg[13][27]  ( .G(n2265), .D(N3371), .Q(
        \REGISTERS[13][27] ) );
  DLH_X1 \REGISTERS_reg[13][26]  ( .G(n2265), .D(N3369), .Q(
        \REGISTERS[13][26] ) );
  DLH_X1 \REGISTERS_reg[13][25]  ( .G(n2265), .D(N3367), .Q(
        \REGISTERS[13][25] ) );
  DLH_X1 \REGISTERS_reg[13][24]  ( .G(n2265), .D(N3365), .Q(
        \REGISTERS[13][24] ) );
  DLH_X1 \REGISTERS_reg[13][23]  ( .G(n2265), .D(N3363), .Q(
        \REGISTERS[13][23] ) );
  DLH_X1 \REGISTERS_reg[13][22]  ( .G(n2265), .D(N3361), .Q(
        \REGISTERS[13][22] ) );
  DLH_X1 \REGISTERS_reg[13][21]  ( .G(n2265), .D(N3359), .Q(
        \REGISTERS[13][21] ) );
  DLH_X1 \REGISTERS_reg[13][20]  ( .G(n2265), .D(N3357), .Q(
        \REGISTERS[13][20] ) );
  DLH_X1 \REGISTERS_reg[13][19]  ( .G(n2265), .D(N3355), .Q(
        \REGISTERS[13][19] ) );
  DLH_X1 \REGISTERS_reg[13][18]  ( .G(n2266), .D(N3353), .Q(
        \REGISTERS[13][18] ) );
  DLH_X1 \REGISTERS_reg[13][17]  ( .G(n2266), .D(N3351), .Q(
        \REGISTERS[13][17] ) );
  DLH_X1 \REGISTERS_reg[13][16]  ( .G(n2266), .D(N3349), .Q(
        \REGISTERS[13][16] ) );
  DLH_X1 \REGISTERS_reg[13][15]  ( .G(n2266), .D(N3347), .Q(
        \REGISTERS[13][15] ) );
  DLH_X1 \REGISTERS_reg[13][14]  ( .G(n2266), .D(N3345), .Q(
        \REGISTERS[13][14] ) );
  DLH_X1 \REGISTERS_reg[13][13]  ( .G(n2266), .D(N3343), .Q(
        \REGISTERS[13][13] ) );
  DLH_X1 \REGISTERS_reg[13][12]  ( .G(n2266), .D(N3341), .Q(
        \REGISTERS[13][12] ) );
  DLH_X1 \REGISTERS_reg[13][11]  ( .G(n2266), .D(N3339), .Q(
        \REGISTERS[13][11] ) );
  DLH_X1 \REGISTERS_reg[13][10]  ( .G(n2266), .D(N3337), .Q(
        \REGISTERS[13][10] ) );
  DLH_X1 \REGISTERS_reg[13][9]  ( .G(n2266), .D(N3335), .Q(\REGISTERS[13][9] )
         );
  DLH_X1 \REGISTERS_reg[13][8]  ( .G(n2266), .D(N3333), .Q(\REGISTERS[13][8] )
         );
  DLH_X1 \REGISTERS_reg[13][7]  ( .G(n2266), .D(N3331), .Q(\REGISTERS[13][7] )
         );
  DLH_X1 \REGISTERS_reg[13][6]  ( .G(n2266), .D(N3329), .Q(\REGISTERS[13][6] )
         );
  DLH_X1 \REGISTERS_reg[13][5]  ( .G(n2267), .D(N3327), .Q(\REGISTERS[13][5] )
         );
  DLH_X1 \REGISTERS_reg[13][4]  ( .G(n2267), .D(N3325), .Q(\REGISTERS[13][4] )
         );
  DLH_X1 \REGISTERS_reg[13][3]  ( .G(n2267), .D(N3323), .Q(\REGISTERS[13][3] )
         );
  DLH_X1 \REGISTERS_reg[13][2]  ( .G(n2267), .D(N3321), .Q(\REGISTERS[13][2] )
         );
  DLH_X1 \REGISTERS_reg[13][1]  ( .G(n2267), .D(N3319), .Q(\REGISTERS[13][1] )
         );
  DLH_X1 \REGISTERS_reg[13][0]  ( .G(n2267), .D(N3317), .Q(\REGISTERS[13][0] )
         );
  DLH_X1 \REGISTERS_reg[12][31]  ( .G(n2268), .D(n1948), .Q(
        \REGISTERS[12][31] ) );
  DLH_X1 \REGISTERS_reg[12][30]  ( .G(n2268), .D(n1947), .Q(
        \REGISTERS[12][30] ) );
  DLH_X1 \REGISTERS_reg[12][29]  ( .G(n2268), .D(n1946), .Q(
        \REGISTERS[12][29] ) );
  DLH_X1 \REGISTERS_reg[12][28]  ( .G(n2268), .D(n1945), .Q(
        \REGISTERS[12][28] ) );
  DLH_X1 \REGISTERS_reg[12][27]  ( .G(n2268), .D(n1944), .Q(
        \REGISTERS[12][27] ) );
  DLH_X1 \REGISTERS_reg[12][26]  ( .G(n2268), .D(n1943), .Q(
        \REGISTERS[12][26] ) );
  DLH_X1 \REGISTERS_reg[12][25]  ( .G(n2268), .D(n1942), .Q(
        \REGISTERS[12][25] ) );
  DLH_X1 \REGISTERS_reg[12][24]  ( .G(n2268), .D(n1941), .Q(
        \REGISTERS[12][24] ) );
  DLH_X1 \REGISTERS_reg[12][23]  ( .G(n2268), .D(n1940), .Q(
        \REGISTERS[12][23] ) );
  DLH_X1 \REGISTERS_reg[12][22]  ( .G(n2268), .D(n1939), .Q(
        \REGISTERS[12][22] ) );
  DLH_X1 \REGISTERS_reg[12][21]  ( .G(n2268), .D(n1938), .Q(
        \REGISTERS[12][21] ) );
  DLH_X1 \REGISTERS_reg[12][20]  ( .G(n2268), .D(n1937), .Q(
        \REGISTERS[12][20] ) );
  DLH_X1 \REGISTERS_reg[12][19]  ( .G(n2268), .D(n1936), .Q(
        \REGISTERS[12][19] ) );
  DLH_X1 \REGISTERS_reg[12][18]  ( .G(n2269), .D(n1935), .Q(
        \REGISTERS[12][18] ) );
  DLH_X1 \REGISTERS_reg[12][17]  ( .G(n2269), .D(n1934), .Q(
        \REGISTERS[12][17] ) );
  DLH_X1 \REGISTERS_reg[12][16]  ( .G(n2269), .D(n1933), .Q(
        \REGISTERS[12][16] ) );
  DLH_X1 \REGISTERS_reg[12][15]  ( .G(n2269), .D(n1932), .Q(
        \REGISTERS[12][15] ) );
  DLH_X1 \REGISTERS_reg[12][14]  ( .G(n2269), .D(n1931), .Q(
        \REGISTERS[12][14] ) );
  DLH_X1 \REGISTERS_reg[12][13]  ( .G(n2269), .D(n1930), .Q(
        \REGISTERS[12][13] ) );
  DLH_X1 \REGISTERS_reg[12][12]  ( .G(n2269), .D(n1929), .Q(
        \REGISTERS[12][12] ) );
  DLH_X1 \REGISTERS_reg[12][11]  ( .G(n2269), .D(n1928), .Q(
        \REGISTERS[12][11] ) );
  DLH_X1 \REGISTERS_reg[12][10]  ( .G(n2269), .D(n1927), .Q(
        \REGISTERS[12][10] ) );
  DLH_X1 \REGISTERS_reg[12][9]  ( .G(n2269), .D(n1926), .Q(\REGISTERS[12][9] )
         );
  DLH_X1 \REGISTERS_reg[12][8]  ( .G(n2269), .D(n1925), .Q(\REGISTERS[12][8] )
         );
  DLH_X1 \REGISTERS_reg[12][7]  ( .G(n2269), .D(n1924), .Q(\REGISTERS[12][7] )
         );
  DLH_X1 \REGISTERS_reg[12][6]  ( .G(n2269), .D(n1923), .Q(\REGISTERS[12][6] )
         );
  DLH_X1 \REGISTERS_reg[12][5]  ( .G(n2270), .D(n1922), .Q(\REGISTERS[12][5] )
         );
  DLH_X1 \REGISTERS_reg[12][4]  ( .G(n2270), .D(n1921), .Q(\REGISTERS[12][4] )
         );
  DLH_X1 \REGISTERS_reg[12][3]  ( .G(n2270), .D(n1920), .Q(\REGISTERS[12][3] )
         );
  DLH_X1 \REGISTERS_reg[12][2]  ( .G(n2270), .D(n1919), .Q(\REGISTERS[12][2] )
         );
  DLH_X1 \REGISTERS_reg[12][1]  ( .G(n2270), .D(n1918), .Q(\REGISTERS[12][1] )
         );
  DLH_X1 \REGISTERS_reg[12][0]  ( .G(n2270), .D(n1917), .Q(\REGISTERS[12][0] )
         );
  DLH_X1 \REGISTERS_reg[11][31]  ( .G(n2271), .D(N3379), .Q(
        \REGISTERS[11][31] ) );
  DLH_X1 \REGISTERS_reg[11][30]  ( .G(n2271), .D(N3377), .Q(
        \REGISTERS[11][30] ) );
  DLH_X1 \REGISTERS_reg[11][29]  ( .G(n2271), .D(N3375), .Q(
        \REGISTERS[11][29] ) );
  DLH_X1 \REGISTERS_reg[11][28]  ( .G(n2271), .D(N3373), .Q(
        \REGISTERS[11][28] ) );
  DLH_X1 \REGISTERS_reg[11][27]  ( .G(n2271), .D(N3371), .Q(
        \REGISTERS[11][27] ) );
  DLH_X1 \REGISTERS_reg[11][26]  ( .G(n2271), .D(N3369), .Q(
        \REGISTERS[11][26] ) );
  DLH_X1 \REGISTERS_reg[11][25]  ( .G(n2271), .D(N3367), .Q(
        \REGISTERS[11][25] ) );
  DLH_X1 \REGISTERS_reg[11][24]  ( .G(n2271), .D(N3365), .Q(
        \REGISTERS[11][24] ) );
  DLH_X1 \REGISTERS_reg[11][23]  ( .G(n2271), .D(N3363), .Q(
        \REGISTERS[11][23] ) );
  DLH_X1 \REGISTERS_reg[11][22]  ( .G(n2271), .D(N3361), .Q(
        \REGISTERS[11][22] ) );
  DLH_X1 \REGISTERS_reg[11][21]  ( .G(n2271), .D(N3359), .Q(
        \REGISTERS[11][21] ) );
  DLH_X1 \REGISTERS_reg[11][20]  ( .G(n2271), .D(N3357), .Q(
        \REGISTERS[11][20] ) );
  DLH_X1 \REGISTERS_reg[11][19]  ( .G(n2271), .D(N3355), .Q(
        \REGISTERS[11][19] ) );
  DLH_X1 \REGISTERS_reg[11][18]  ( .G(n2272), .D(N3353), .Q(
        \REGISTERS[11][18] ) );
  DLH_X1 \REGISTERS_reg[11][17]  ( .G(n2272), .D(N3351), .Q(
        \REGISTERS[11][17] ) );
  DLH_X1 \REGISTERS_reg[11][16]  ( .G(n2272), .D(N3349), .Q(
        \REGISTERS[11][16] ) );
  DLH_X1 \REGISTERS_reg[11][15]  ( .G(n2272), .D(N3347), .Q(
        \REGISTERS[11][15] ) );
  DLH_X1 \REGISTERS_reg[11][14]  ( .G(n2272), .D(N3345), .Q(
        \REGISTERS[11][14] ) );
  DLH_X1 \REGISTERS_reg[11][13]  ( .G(n2272), .D(N3343), .Q(
        \REGISTERS[11][13] ) );
  DLH_X1 \REGISTERS_reg[11][12]  ( .G(n2272), .D(N3341), .Q(
        \REGISTERS[11][12] ) );
  DLH_X1 \REGISTERS_reg[11][11]  ( .G(n2272), .D(N3339), .Q(
        \REGISTERS[11][11] ) );
  DLH_X1 \REGISTERS_reg[11][10]  ( .G(n2272), .D(N3337), .Q(
        \REGISTERS[11][10] ) );
  DLH_X1 \REGISTERS_reg[11][9]  ( .G(n2272), .D(N3335), .Q(\REGISTERS[11][9] )
         );
  DLH_X1 \REGISTERS_reg[11][8]  ( .G(n2272), .D(N3333), .Q(\REGISTERS[11][8] )
         );
  DLH_X1 \REGISTERS_reg[11][7]  ( .G(n2272), .D(N3331), .Q(\REGISTERS[11][7] )
         );
  DLH_X1 \REGISTERS_reg[11][6]  ( .G(n2272), .D(N3329), .Q(\REGISTERS[11][6] )
         );
  DLH_X1 \REGISTERS_reg[11][5]  ( .G(n2273), .D(N3327), .Q(\REGISTERS[11][5] )
         );
  DLH_X1 \REGISTERS_reg[11][4]  ( .G(n2273), .D(N3325), .Q(\REGISTERS[11][4] )
         );
  DLH_X1 \REGISTERS_reg[11][3]  ( .G(n2273), .D(N3323), .Q(\REGISTERS[11][3] )
         );
  DLH_X1 \REGISTERS_reg[11][2]  ( .G(n2273), .D(N3321), .Q(\REGISTERS[11][2] )
         );
  DLH_X1 \REGISTERS_reg[11][1]  ( .G(n2273), .D(N3319), .Q(\REGISTERS[11][1] )
         );
  DLH_X1 \REGISTERS_reg[11][0]  ( .G(n2273), .D(N3317), .Q(\REGISTERS[11][0] )
         );
  DLH_X1 \REGISTERS_reg[10][31]  ( .G(n2274), .D(n1948), .Q(
        \REGISTERS[10][31] ) );
  DLH_X1 \REGISTERS_reg[10][30]  ( .G(n2274), .D(n1947), .Q(
        \REGISTERS[10][30] ) );
  DLH_X1 \REGISTERS_reg[10][29]  ( .G(n2274), .D(n1946), .Q(
        \REGISTERS[10][29] ) );
  DLH_X1 \REGISTERS_reg[10][28]  ( .G(n2274), .D(n1945), .Q(
        \REGISTERS[10][28] ) );
  DLH_X1 \REGISTERS_reg[10][27]  ( .G(n2274), .D(n1944), .Q(
        \REGISTERS[10][27] ) );
  DLH_X1 \REGISTERS_reg[10][26]  ( .G(n2274), .D(n1943), .Q(
        \REGISTERS[10][26] ) );
  DLH_X1 \REGISTERS_reg[10][25]  ( .G(n2274), .D(n1942), .Q(
        \REGISTERS[10][25] ) );
  DLH_X1 \REGISTERS_reg[10][24]  ( .G(n2274), .D(n1941), .Q(
        \REGISTERS[10][24] ) );
  DLH_X1 \REGISTERS_reg[10][23]  ( .G(n2274), .D(n1940), .Q(
        \REGISTERS[10][23] ) );
  DLH_X1 \REGISTERS_reg[10][22]  ( .G(n2274), .D(n1939), .Q(
        \REGISTERS[10][22] ) );
  DLH_X1 \REGISTERS_reg[10][21]  ( .G(n2274), .D(n1938), .Q(
        \REGISTERS[10][21] ) );
  DLH_X1 \REGISTERS_reg[10][20]  ( .G(n2274), .D(n1937), .Q(
        \REGISTERS[10][20] ) );
  DLH_X1 \REGISTERS_reg[10][19]  ( .G(n2274), .D(n1936), .Q(
        \REGISTERS[10][19] ) );
  DLH_X1 \REGISTERS_reg[10][18]  ( .G(n2275), .D(n1935), .Q(
        \REGISTERS[10][18] ) );
  DLH_X1 \REGISTERS_reg[10][17]  ( .G(n2275), .D(n1934), .Q(
        \REGISTERS[10][17] ) );
  DLH_X1 \REGISTERS_reg[10][16]  ( .G(n2275), .D(n1933), .Q(
        \REGISTERS[10][16] ) );
  DLH_X1 \REGISTERS_reg[10][15]  ( .G(n2275), .D(n1932), .Q(
        \REGISTERS[10][15] ) );
  DLH_X1 \REGISTERS_reg[10][14]  ( .G(n2275), .D(n1931), .Q(
        \REGISTERS[10][14] ) );
  DLH_X1 \REGISTERS_reg[10][13]  ( .G(n2275), .D(n1930), .Q(
        \REGISTERS[10][13] ) );
  DLH_X1 \REGISTERS_reg[10][12]  ( .G(n2275), .D(n1929), .Q(
        \REGISTERS[10][12] ) );
  DLH_X1 \REGISTERS_reg[10][11]  ( .G(n2275), .D(n1928), .Q(
        \REGISTERS[10][11] ) );
  DLH_X1 \REGISTERS_reg[10][10]  ( .G(n2275), .D(n1927), .Q(
        \REGISTERS[10][10] ) );
  DLH_X1 \REGISTERS_reg[10][9]  ( .G(n2275), .D(n1926), .Q(\REGISTERS[10][9] )
         );
  DLH_X1 \REGISTERS_reg[10][8]  ( .G(n2275), .D(n1925), .Q(\REGISTERS[10][8] )
         );
  DLH_X1 \REGISTERS_reg[10][7]  ( .G(n2275), .D(n1924), .Q(\REGISTERS[10][7] )
         );
  DLH_X1 \REGISTERS_reg[10][6]  ( .G(n2275), .D(n1923), .Q(\REGISTERS[10][6] )
         );
  DLH_X1 \REGISTERS_reg[10][5]  ( .G(n2276), .D(n1922), .Q(\REGISTERS[10][5] )
         );
  DLH_X1 \REGISTERS_reg[10][4]  ( .G(n2276), .D(n1921), .Q(\REGISTERS[10][4] )
         );
  DLH_X1 \REGISTERS_reg[10][3]  ( .G(n2276), .D(n1920), .Q(\REGISTERS[10][3] )
         );
  DLH_X1 \REGISTERS_reg[10][2]  ( .G(n2276), .D(n1919), .Q(\REGISTERS[10][2] )
         );
  DLH_X1 \REGISTERS_reg[10][1]  ( .G(n2276), .D(n1918), .Q(\REGISTERS[10][1] )
         );
  DLH_X1 \REGISTERS_reg[10][0]  ( .G(n2276), .D(n1917), .Q(\REGISTERS[10][0] )
         );
  DLH_X1 \REGISTERS_reg[9][31]  ( .G(n2277), .D(N3379), .Q(\REGISTERS[9][31] )
         );
  DLH_X1 \REGISTERS_reg[9][30]  ( .G(n2277), .D(N3377), .Q(\REGISTERS[9][30] )
         );
  DLH_X1 \REGISTERS_reg[9][29]  ( .G(n2277), .D(N3375), .Q(\REGISTERS[9][29] )
         );
  DLH_X1 \REGISTERS_reg[9][28]  ( .G(n2277), .D(N3373), .Q(\REGISTERS[9][28] )
         );
  DLH_X1 \REGISTERS_reg[9][27]  ( .G(n2277), .D(N3371), .Q(\REGISTERS[9][27] )
         );
  DLH_X1 \REGISTERS_reg[9][26]  ( .G(n2277), .D(N3369), .Q(\REGISTERS[9][26] )
         );
  DLH_X1 \REGISTERS_reg[9][25]  ( .G(n2277), .D(N3367), .Q(\REGISTERS[9][25] )
         );
  DLH_X1 \REGISTERS_reg[9][24]  ( .G(n2277), .D(N3365), .Q(\REGISTERS[9][24] )
         );
  DLH_X1 \REGISTERS_reg[9][23]  ( .G(n2277), .D(N3363), .Q(\REGISTERS[9][23] )
         );
  DLH_X1 \REGISTERS_reg[9][22]  ( .G(n2277), .D(N3361), .Q(\REGISTERS[9][22] )
         );
  DLH_X1 \REGISTERS_reg[9][21]  ( .G(n2277), .D(N3359), .Q(\REGISTERS[9][21] )
         );
  DLH_X1 \REGISTERS_reg[9][20]  ( .G(n2277), .D(N3357), .Q(\REGISTERS[9][20] )
         );
  DLH_X1 \REGISTERS_reg[9][19]  ( .G(n2277), .D(N3355), .Q(\REGISTERS[9][19] )
         );
  DLH_X1 \REGISTERS_reg[9][18]  ( .G(n2278), .D(N3353), .Q(\REGISTERS[9][18] )
         );
  DLH_X1 \REGISTERS_reg[9][17]  ( .G(n2278), .D(N3351), .Q(\REGISTERS[9][17] )
         );
  DLH_X1 \REGISTERS_reg[9][16]  ( .G(n2278), .D(N3349), .Q(\REGISTERS[9][16] )
         );
  DLH_X1 \REGISTERS_reg[9][15]  ( .G(n2278), .D(N3347), .Q(\REGISTERS[9][15] )
         );
  DLH_X1 \REGISTERS_reg[9][14]  ( .G(n2278), .D(N3345), .Q(\REGISTERS[9][14] )
         );
  DLH_X1 \REGISTERS_reg[9][13]  ( .G(n2278), .D(N3343), .Q(\REGISTERS[9][13] )
         );
  DLH_X1 \REGISTERS_reg[9][12]  ( .G(n2278), .D(N3341), .Q(\REGISTERS[9][12] )
         );
  DLH_X1 \REGISTERS_reg[9][11]  ( .G(n2278), .D(N3339), .Q(\REGISTERS[9][11] )
         );
  DLH_X1 \REGISTERS_reg[9][10]  ( .G(n2278), .D(N3337), .Q(\REGISTERS[9][10] )
         );
  DLH_X1 \REGISTERS_reg[9][9]  ( .G(n2278), .D(N3335), .Q(\REGISTERS[9][9] )
         );
  DLH_X1 \REGISTERS_reg[9][8]  ( .G(n2278), .D(N3333), .Q(\REGISTERS[9][8] )
         );
  DLH_X1 \REGISTERS_reg[9][7]  ( .G(n2278), .D(N3331), .Q(\REGISTERS[9][7] )
         );
  DLH_X1 \REGISTERS_reg[9][6]  ( .G(n2278), .D(N3329), .Q(\REGISTERS[9][6] )
         );
  DLH_X1 \REGISTERS_reg[9][5]  ( .G(n2279), .D(N3327), .Q(\REGISTERS[9][5] )
         );
  DLH_X1 \REGISTERS_reg[9][4]  ( .G(n2279), .D(N3325), .Q(\REGISTERS[9][4] )
         );
  DLH_X1 \REGISTERS_reg[9][3]  ( .G(n2279), .D(N3323), .Q(\REGISTERS[9][3] )
         );
  DLH_X1 \REGISTERS_reg[9][2]  ( .G(n2279), .D(N3321), .Q(\REGISTERS[9][2] )
         );
  DLH_X1 \REGISTERS_reg[9][1]  ( .G(n2279), .D(N3319), .Q(\REGISTERS[9][1] )
         );
  DLH_X1 \REGISTERS_reg[9][0]  ( .G(n2279), .D(N3317), .Q(\REGISTERS[9][0] )
         );
  DLH_X1 \REGISTERS_reg[8][31]  ( .G(n2280), .D(n1948), .Q(\REGISTERS[8][31] )
         );
  DLH_X1 \REGISTERS_reg[8][30]  ( .G(n2280), .D(n1947), .Q(\REGISTERS[8][30] )
         );
  DLH_X1 \REGISTERS_reg[8][29]  ( .G(n2280), .D(n1946), .Q(\REGISTERS[8][29] )
         );
  DLH_X1 \REGISTERS_reg[8][28]  ( .G(n2280), .D(n1945), .Q(\REGISTERS[8][28] )
         );
  DLH_X1 \REGISTERS_reg[8][27]  ( .G(n2280), .D(n1944), .Q(\REGISTERS[8][27] )
         );
  DLH_X1 \REGISTERS_reg[8][26]  ( .G(n2280), .D(n1943), .Q(\REGISTERS[8][26] )
         );
  DLH_X1 \REGISTERS_reg[8][25]  ( .G(n2280), .D(n1942), .Q(\REGISTERS[8][25] )
         );
  DLH_X1 \REGISTERS_reg[8][24]  ( .G(n2280), .D(n1941), .Q(\REGISTERS[8][24] )
         );
  DLH_X1 \REGISTERS_reg[8][23]  ( .G(n2280), .D(n1940), .Q(\REGISTERS[8][23] )
         );
  DLH_X1 \REGISTERS_reg[8][22]  ( .G(n2280), .D(n1939), .Q(\REGISTERS[8][22] )
         );
  DLH_X1 \REGISTERS_reg[8][21]  ( .G(n2280), .D(n1938), .Q(\REGISTERS[8][21] )
         );
  DLH_X1 \REGISTERS_reg[8][20]  ( .G(n2280), .D(n1937), .Q(\REGISTERS[8][20] )
         );
  DLH_X1 \REGISTERS_reg[8][19]  ( .G(n2280), .D(n1936), .Q(\REGISTERS[8][19] )
         );
  DLH_X1 \REGISTERS_reg[8][18]  ( .G(n2281), .D(n1935), .Q(\REGISTERS[8][18] )
         );
  DLH_X1 \REGISTERS_reg[8][17]  ( .G(n2281), .D(n1934), .Q(\REGISTERS[8][17] )
         );
  DLH_X1 \REGISTERS_reg[8][16]  ( .G(n2281), .D(n1933), .Q(\REGISTERS[8][16] )
         );
  DLH_X1 \REGISTERS_reg[8][15]  ( .G(n2281), .D(n1932), .Q(\REGISTERS[8][15] )
         );
  DLH_X1 \REGISTERS_reg[8][14]  ( .G(n2281), .D(n1931), .Q(\REGISTERS[8][14] )
         );
  DLH_X1 \REGISTERS_reg[8][13]  ( .G(n2281), .D(n1930), .Q(\REGISTERS[8][13] )
         );
  DLH_X1 \REGISTERS_reg[8][12]  ( .G(n2281), .D(n1929), .Q(\REGISTERS[8][12] )
         );
  DLH_X1 \REGISTERS_reg[8][11]  ( .G(n2281), .D(n1928), .Q(\REGISTERS[8][11] )
         );
  DLH_X1 \REGISTERS_reg[8][10]  ( .G(n2281), .D(n1927), .Q(\REGISTERS[8][10] )
         );
  DLH_X1 \REGISTERS_reg[8][9]  ( .G(n2281), .D(n1926), .Q(\REGISTERS[8][9] )
         );
  DLH_X1 \REGISTERS_reg[8][8]  ( .G(n2281), .D(n1925), .Q(\REGISTERS[8][8] )
         );
  DLH_X1 \REGISTERS_reg[8][7]  ( .G(n2281), .D(n1924), .Q(\REGISTERS[8][7] )
         );
  DLH_X1 \REGISTERS_reg[8][6]  ( .G(n2281), .D(n1923), .Q(\REGISTERS[8][6] )
         );
  DLH_X1 \REGISTERS_reg[8][5]  ( .G(n2282), .D(n1922), .Q(\REGISTERS[8][5] )
         );
  DLH_X1 \REGISTERS_reg[8][4]  ( .G(n2282), .D(n1921), .Q(\REGISTERS[8][4] )
         );
  DLH_X1 \REGISTERS_reg[8][3]  ( .G(n2282), .D(n1920), .Q(\REGISTERS[8][3] )
         );
  DLH_X1 \REGISTERS_reg[8][2]  ( .G(n2282), .D(n1919), .Q(\REGISTERS[8][2] )
         );
  DLH_X1 \REGISTERS_reg[8][1]  ( .G(n2282), .D(n1918), .Q(\REGISTERS[8][1] )
         );
  DLH_X1 \REGISTERS_reg[8][0]  ( .G(n2282), .D(n1917), .Q(\REGISTERS[8][0] )
         );
  DLH_X1 \REGISTERS_reg[7][31]  ( .G(n2283), .D(N3379), .Q(\REGISTERS[7][31] )
         );
  DLH_X1 \REGISTERS_reg[7][30]  ( .G(n2283), .D(N3377), .Q(\REGISTERS[7][30] )
         );
  DLH_X1 \REGISTERS_reg[7][29]  ( .G(n2283), .D(N3375), .Q(\REGISTERS[7][29] )
         );
  DLH_X1 \REGISTERS_reg[7][28]  ( .G(n2283), .D(N3373), .Q(\REGISTERS[7][28] )
         );
  DLH_X1 \REGISTERS_reg[7][27]  ( .G(n2283), .D(N3371), .Q(\REGISTERS[7][27] )
         );
  DLH_X1 \REGISTERS_reg[7][26]  ( .G(n2283), .D(N3369), .Q(\REGISTERS[7][26] )
         );
  DLH_X1 \REGISTERS_reg[7][25]  ( .G(n2283), .D(N3367), .Q(\REGISTERS[7][25] )
         );
  DLH_X1 \REGISTERS_reg[7][24]  ( .G(n2283), .D(N3365), .Q(\REGISTERS[7][24] )
         );
  DLH_X1 \REGISTERS_reg[7][23]  ( .G(n2283), .D(N3363), .Q(\REGISTERS[7][23] )
         );
  DLH_X1 \REGISTERS_reg[7][22]  ( .G(n2283), .D(N3361), .Q(\REGISTERS[7][22] )
         );
  DLH_X1 \REGISTERS_reg[7][21]  ( .G(n2283), .D(N3359), .Q(\REGISTERS[7][21] )
         );
  DLH_X1 \REGISTERS_reg[7][20]  ( .G(n2283), .D(N3357), .Q(\REGISTERS[7][20] )
         );
  DLH_X1 \REGISTERS_reg[7][19]  ( .G(n2283), .D(N3355), .Q(\REGISTERS[7][19] )
         );
  DLH_X1 \REGISTERS_reg[7][18]  ( .G(n2284), .D(N3353), .Q(\REGISTERS[7][18] )
         );
  DLH_X1 \REGISTERS_reg[7][17]  ( .G(n2284), .D(N3351), .Q(\REGISTERS[7][17] )
         );
  DLH_X1 \REGISTERS_reg[7][16]  ( .G(n2284), .D(N3349), .Q(\REGISTERS[7][16] )
         );
  DLH_X1 \REGISTERS_reg[7][15]  ( .G(n2284), .D(N3347), .Q(\REGISTERS[7][15] )
         );
  DLH_X1 \REGISTERS_reg[7][14]  ( .G(n2284), .D(N3345), .Q(\REGISTERS[7][14] )
         );
  DLH_X1 \REGISTERS_reg[7][13]  ( .G(n2284), .D(N3343), .Q(\REGISTERS[7][13] )
         );
  DLH_X1 \REGISTERS_reg[7][12]  ( .G(n2284), .D(N3341), .Q(\REGISTERS[7][12] )
         );
  DLH_X1 \REGISTERS_reg[7][11]  ( .G(n2284), .D(N3339), .Q(\REGISTERS[7][11] )
         );
  DLH_X1 \REGISTERS_reg[7][10]  ( .G(n2284), .D(N3337), .Q(\REGISTERS[7][10] )
         );
  DLH_X1 \REGISTERS_reg[7][9]  ( .G(n2284), .D(N3335), .Q(\REGISTERS[7][9] )
         );
  DLH_X1 \REGISTERS_reg[7][8]  ( .G(n2284), .D(N3333), .Q(\REGISTERS[7][8] )
         );
  DLH_X1 \REGISTERS_reg[7][7]  ( .G(n2284), .D(N3331), .Q(\REGISTERS[7][7] )
         );
  DLH_X1 \REGISTERS_reg[7][6]  ( .G(n2284), .D(N3329), .Q(\REGISTERS[7][6] )
         );
  DLH_X1 \REGISTERS_reg[7][5]  ( .G(n2285), .D(N3327), .Q(\REGISTERS[7][5] )
         );
  DLH_X1 \REGISTERS_reg[7][4]  ( .G(n2285), .D(N3325), .Q(\REGISTERS[7][4] )
         );
  DLH_X1 \REGISTERS_reg[7][3]  ( .G(n2285), .D(N3323), .Q(\REGISTERS[7][3] )
         );
  DLH_X1 \REGISTERS_reg[7][2]  ( .G(n2285), .D(N3321), .Q(\REGISTERS[7][2] )
         );
  DLH_X1 \REGISTERS_reg[7][1]  ( .G(n2285), .D(N3319), .Q(\REGISTERS[7][1] )
         );
  DLH_X1 \REGISTERS_reg[7][0]  ( .G(n2285), .D(N3317), .Q(\REGISTERS[7][0] )
         );
  DLH_X1 \REGISTERS_reg[6][31]  ( .G(n2286), .D(n1948), .Q(\REGISTERS[6][31] )
         );
  DLH_X1 \REGISTERS_reg[6][30]  ( .G(n2286), .D(n1947), .Q(\REGISTERS[6][30] )
         );
  DLH_X1 \REGISTERS_reg[6][29]  ( .G(n2286), .D(n1946), .Q(\REGISTERS[6][29] )
         );
  DLH_X1 \REGISTERS_reg[6][28]  ( .G(n2286), .D(n1945), .Q(\REGISTERS[6][28] )
         );
  DLH_X1 \REGISTERS_reg[6][27]  ( .G(n2286), .D(n1944), .Q(\REGISTERS[6][27] )
         );
  DLH_X1 \REGISTERS_reg[6][26]  ( .G(n2286), .D(n1943), .Q(\REGISTERS[6][26] )
         );
  DLH_X1 \REGISTERS_reg[6][25]  ( .G(n2286), .D(n1942), .Q(\REGISTERS[6][25] )
         );
  DLH_X1 \REGISTERS_reg[6][24]  ( .G(n2286), .D(n1941), .Q(\REGISTERS[6][24] )
         );
  DLH_X1 \REGISTERS_reg[6][23]  ( .G(n2286), .D(n1940), .Q(\REGISTERS[6][23] )
         );
  DLH_X1 \REGISTERS_reg[6][22]  ( .G(n2286), .D(n1939), .Q(\REGISTERS[6][22] )
         );
  DLH_X1 \REGISTERS_reg[6][21]  ( .G(n2286), .D(n1938), .Q(\REGISTERS[6][21] )
         );
  DLH_X1 \REGISTERS_reg[6][20]  ( .G(n2286), .D(n1937), .Q(\REGISTERS[6][20] )
         );
  DLH_X1 \REGISTERS_reg[6][19]  ( .G(n2286), .D(n1936), .Q(\REGISTERS[6][19] )
         );
  DLH_X1 \REGISTERS_reg[6][18]  ( .G(n2287), .D(n1935), .Q(\REGISTERS[6][18] )
         );
  DLH_X1 \REGISTERS_reg[6][17]  ( .G(n2287), .D(n1934), .Q(\REGISTERS[6][17] )
         );
  DLH_X1 \REGISTERS_reg[6][16]  ( .G(n2287), .D(n1933), .Q(\REGISTERS[6][16] )
         );
  DLH_X1 \REGISTERS_reg[6][15]  ( .G(n2287), .D(n1932), .Q(\REGISTERS[6][15] )
         );
  DLH_X1 \REGISTERS_reg[6][14]  ( .G(n2287), .D(n1931), .Q(\REGISTERS[6][14] )
         );
  DLH_X1 \REGISTERS_reg[6][13]  ( .G(n2287), .D(n1930), .Q(\REGISTERS[6][13] )
         );
  DLH_X1 \REGISTERS_reg[6][12]  ( .G(n2287), .D(n1929), .Q(\REGISTERS[6][12] )
         );
  DLH_X1 \REGISTERS_reg[6][11]  ( .G(n2287), .D(n1928), .Q(\REGISTERS[6][11] )
         );
  DLH_X1 \REGISTERS_reg[6][10]  ( .G(n2287), .D(n1927), .Q(\REGISTERS[6][10] )
         );
  DLH_X1 \REGISTERS_reg[6][9]  ( .G(n2287), .D(n1926), .Q(\REGISTERS[6][9] )
         );
  DLH_X1 \REGISTERS_reg[6][8]  ( .G(n2287), .D(n1925), .Q(\REGISTERS[6][8] )
         );
  DLH_X1 \REGISTERS_reg[6][7]  ( .G(n2287), .D(n1924), .Q(\REGISTERS[6][7] )
         );
  DLH_X1 \REGISTERS_reg[6][6]  ( .G(n2287), .D(n1923), .Q(\REGISTERS[6][6] )
         );
  DLH_X1 \REGISTERS_reg[6][5]  ( .G(n2288), .D(n1922), .Q(\REGISTERS[6][5] )
         );
  DLH_X1 \REGISTERS_reg[6][4]  ( .G(n2288), .D(n1921), .Q(\REGISTERS[6][4] )
         );
  DLH_X1 \REGISTERS_reg[6][3]  ( .G(n2288), .D(n1920), .Q(\REGISTERS[6][3] )
         );
  DLH_X1 \REGISTERS_reg[6][2]  ( .G(n2288), .D(n1919), .Q(\REGISTERS[6][2] )
         );
  DLH_X1 \REGISTERS_reg[6][1]  ( .G(n2288), .D(n1918), .Q(\REGISTERS[6][1] )
         );
  DLH_X1 \REGISTERS_reg[6][0]  ( .G(n2288), .D(n1917), .Q(\REGISTERS[6][0] )
         );
  DLH_X1 \REGISTERS_reg[5][31]  ( .G(n2289), .D(N3379), .Q(\REGISTERS[5][31] )
         );
  DLH_X1 \REGISTERS_reg[5][30]  ( .G(n2289), .D(N3377), .Q(\REGISTERS[5][30] )
         );
  DLH_X1 \REGISTERS_reg[5][29]  ( .G(n2289), .D(N3375), .Q(\REGISTERS[5][29] )
         );
  DLH_X1 \REGISTERS_reg[5][28]  ( .G(n2289), .D(N3373), .Q(\REGISTERS[5][28] )
         );
  DLH_X1 \REGISTERS_reg[5][27]  ( .G(n2289), .D(N3371), .Q(\REGISTERS[5][27] )
         );
  DLH_X1 \REGISTERS_reg[5][26]  ( .G(n2289), .D(N3369), .Q(\REGISTERS[5][26] )
         );
  DLH_X1 \REGISTERS_reg[5][25]  ( .G(n2289), .D(N3367), .Q(\REGISTERS[5][25] )
         );
  DLH_X1 \REGISTERS_reg[5][24]  ( .G(n2289), .D(N3365), .Q(\REGISTERS[5][24] )
         );
  DLH_X1 \REGISTERS_reg[5][23]  ( .G(n2289), .D(N3363), .Q(\REGISTERS[5][23] )
         );
  DLH_X1 \REGISTERS_reg[5][22]  ( .G(n2289), .D(N3361), .Q(\REGISTERS[5][22] )
         );
  DLH_X1 \REGISTERS_reg[5][21]  ( .G(n2289), .D(N3359), .Q(\REGISTERS[5][21] )
         );
  DLH_X1 \REGISTERS_reg[5][20]  ( .G(n2289), .D(N3357), .Q(\REGISTERS[5][20] )
         );
  DLH_X1 \REGISTERS_reg[5][19]  ( .G(n2289), .D(N3355), .Q(\REGISTERS[5][19] )
         );
  DLH_X1 \REGISTERS_reg[5][18]  ( .G(n2290), .D(N3353), .Q(\REGISTERS[5][18] )
         );
  DLH_X1 \REGISTERS_reg[5][17]  ( .G(n2290), .D(N3351), .Q(\REGISTERS[5][17] )
         );
  DLH_X1 \REGISTERS_reg[5][16]  ( .G(n2290), .D(N3349), .Q(\REGISTERS[5][16] )
         );
  DLH_X1 \REGISTERS_reg[5][15]  ( .G(n2290), .D(N3347), .Q(\REGISTERS[5][15] )
         );
  DLH_X1 \REGISTERS_reg[5][14]  ( .G(n2290), .D(N3345), .Q(\REGISTERS[5][14] )
         );
  DLH_X1 \REGISTERS_reg[5][13]  ( .G(n2290), .D(N3343), .Q(\REGISTERS[5][13] )
         );
  DLH_X1 \REGISTERS_reg[5][12]  ( .G(n2290), .D(N3341), .Q(\REGISTERS[5][12] )
         );
  DLH_X1 \REGISTERS_reg[5][11]  ( .G(n2290), .D(N3339), .Q(\REGISTERS[5][11] )
         );
  DLH_X1 \REGISTERS_reg[5][10]  ( .G(n2290), .D(N3337), .Q(\REGISTERS[5][10] )
         );
  DLH_X1 \REGISTERS_reg[5][9]  ( .G(n2290), .D(N3335), .Q(\REGISTERS[5][9] )
         );
  DLH_X1 \REGISTERS_reg[5][8]  ( .G(n2290), .D(N3333), .Q(\REGISTERS[5][8] )
         );
  DLH_X1 \REGISTERS_reg[5][7]  ( .G(n2290), .D(N3331), .Q(\REGISTERS[5][7] )
         );
  DLH_X1 \REGISTERS_reg[5][6]  ( .G(n2290), .D(N3329), .Q(\REGISTERS[5][6] )
         );
  DLH_X1 \REGISTERS_reg[5][5]  ( .G(n2291), .D(N3327), .Q(\REGISTERS[5][5] )
         );
  DLH_X1 \REGISTERS_reg[5][4]  ( .G(n2291), .D(N3325), .Q(\REGISTERS[5][4] )
         );
  DLH_X1 \REGISTERS_reg[5][3]  ( .G(n2291), .D(N3323), .Q(\REGISTERS[5][3] )
         );
  DLH_X1 \REGISTERS_reg[5][2]  ( .G(n2291), .D(N3321), .Q(\REGISTERS[5][2] )
         );
  DLH_X1 \REGISTERS_reg[5][1]  ( .G(n2291), .D(N3319), .Q(\REGISTERS[5][1] )
         );
  DLH_X1 \REGISTERS_reg[5][0]  ( .G(n2291), .D(N3317), .Q(\REGISTERS[5][0] )
         );
  DLH_X1 \REGISTERS_reg[4][31]  ( .G(n2292), .D(n1948), .Q(\REGISTERS[4][31] )
         );
  DLH_X1 \REGISTERS_reg[4][30]  ( .G(n2292), .D(n1947), .Q(\REGISTERS[4][30] )
         );
  DLH_X1 \REGISTERS_reg[4][29]  ( .G(n2292), .D(n1946), .Q(\REGISTERS[4][29] )
         );
  DLH_X1 \REGISTERS_reg[4][28]  ( .G(n2292), .D(n1945), .Q(\REGISTERS[4][28] )
         );
  DLH_X1 \REGISTERS_reg[4][27]  ( .G(n2292), .D(n1944), .Q(\REGISTERS[4][27] )
         );
  DLH_X1 \REGISTERS_reg[4][26]  ( .G(n2292), .D(n1943), .Q(\REGISTERS[4][26] )
         );
  DLH_X1 \REGISTERS_reg[4][25]  ( .G(n2292), .D(n1942), .Q(\REGISTERS[4][25] )
         );
  DLH_X1 \REGISTERS_reg[4][24]  ( .G(n2292), .D(n1941), .Q(\REGISTERS[4][24] )
         );
  DLH_X1 \REGISTERS_reg[4][23]  ( .G(n2292), .D(n1940), .Q(\REGISTERS[4][23] )
         );
  DLH_X1 \REGISTERS_reg[4][22]  ( .G(n2292), .D(n1939), .Q(\REGISTERS[4][22] )
         );
  DLH_X1 \REGISTERS_reg[4][21]  ( .G(n2292), .D(n1938), .Q(\REGISTERS[4][21] )
         );
  DLH_X1 \REGISTERS_reg[4][20]  ( .G(n2292), .D(n1937), .Q(\REGISTERS[4][20] )
         );
  DLH_X1 \REGISTERS_reg[4][19]  ( .G(n2292), .D(n1936), .Q(\REGISTERS[4][19] )
         );
  DLH_X1 \REGISTERS_reg[4][18]  ( .G(n2293), .D(n1935), .Q(\REGISTERS[4][18] )
         );
  DLH_X1 \REGISTERS_reg[4][17]  ( .G(n2293), .D(n1934), .Q(\REGISTERS[4][17] )
         );
  DLH_X1 \REGISTERS_reg[4][16]  ( .G(n2293), .D(n1933), .Q(\REGISTERS[4][16] )
         );
  DLH_X1 \REGISTERS_reg[4][15]  ( .G(n2293), .D(n1932), .Q(\REGISTERS[4][15] )
         );
  DLH_X1 \REGISTERS_reg[4][14]  ( .G(n2293), .D(n1931), .Q(\REGISTERS[4][14] )
         );
  DLH_X1 \REGISTERS_reg[4][13]  ( .G(n2293), .D(n1930), .Q(\REGISTERS[4][13] )
         );
  DLH_X1 \REGISTERS_reg[4][12]  ( .G(n2293), .D(n1929), .Q(\REGISTERS[4][12] )
         );
  DLH_X1 \REGISTERS_reg[4][11]  ( .G(n2293), .D(n1928), .Q(\REGISTERS[4][11] )
         );
  DLH_X1 \REGISTERS_reg[4][10]  ( .G(n2293), .D(n1927), .Q(\REGISTERS[4][10] )
         );
  DLH_X1 \REGISTERS_reg[4][9]  ( .G(n2293), .D(n1926), .Q(\REGISTERS[4][9] )
         );
  DLH_X1 \REGISTERS_reg[4][8]  ( .G(n2293), .D(n1925), .Q(\REGISTERS[4][8] )
         );
  DLH_X1 \REGISTERS_reg[4][7]  ( .G(n2293), .D(n1924), .Q(\REGISTERS[4][7] )
         );
  DLH_X1 \REGISTERS_reg[4][6]  ( .G(n2293), .D(n1923), .Q(\REGISTERS[4][6] )
         );
  DLH_X1 \REGISTERS_reg[4][5]  ( .G(n2294), .D(n1922), .Q(\REGISTERS[4][5] )
         );
  DLH_X1 \REGISTERS_reg[4][4]  ( .G(n2294), .D(n1921), .Q(\REGISTERS[4][4] )
         );
  DLH_X1 \REGISTERS_reg[4][3]  ( .G(n2294), .D(n1920), .Q(\REGISTERS[4][3] )
         );
  DLH_X1 \REGISTERS_reg[4][2]  ( .G(n2294), .D(n1919), .Q(\REGISTERS[4][2] )
         );
  DLH_X1 \REGISTERS_reg[4][1]  ( .G(n2294), .D(n1918), .Q(\REGISTERS[4][1] )
         );
  DLH_X1 \REGISTERS_reg[4][0]  ( .G(n2294), .D(n1917), .Q(\REGISTERS[4][0] )
         );
  DLH_X1 \REGISTERS_reg[3][31]  ( .G(n2295), .D(N3379), .Q(\REGISTERS[3][31] )
         );
  DLH_X1 \REGISTERS_reg[3][30]  ( .G(n2295), .D(N3377), .Q(\REGISTERS[3][30] )
         );
  DLH_X1 \REGISTERS_reg[3][29]  ( .G(n2295), .D(N3375), .Q(\REGISTERS[3][29] )
         );
  DLH_X1 \REGISTERS_reg[3][28]  ( .G(n2295), .D(N3373), .Q(\REGISTERS[3][28] )
         );
  DLH_X1 \REGISTERS_reg[3][27]  ( .G(n2295), .D(N3371), .Q(\REGISTERS[3][27] )
         );
  DLH_X1 \REGISTERS_reg[3][26]  ( .G(n2295), .D(N3369), .Q(\REGISTERS[3][26] )
         );
  DLH_X1 \REGISTERS_reg[3][25]  ( .G(n2295), .D(N3367), .Q(\REGISTERS[3][25] )
         );
  DLH_X1 \REGISTERS_reg[3][24]  ( .G(n2295), .D(N3365), .Q(\REGISTERS[3][24] )
         );
  DLH_X1 \REGISTERS_reg[3][23]  ( .G(n2295), .D(N3363), .Q(\REGISTERS[3][23] )
         );
  DLH_X1 \REGISTERS_reg[3][22]  ( .G(n2295), .D(N3361), .Q(\REGISTERS[3][22] )
         );
  DLH_X1 \REGISTERS_reg[3][21]  ( .G(n2295), .D(N3359), .Q(\REGISTERS[3][21] )
         );
  DLH_X1 \REGISTERS_reg[3][20]  ( .G(n2295), .D(N3357), .Q(\REGISTERS[3][20] )
         );
  DLH_X1 \REGISTERS_reg[3][19]  ( .G(n2295), .D(N3355), .Q(\REGISTERS[3][19] )
         );
  DLH_X1 \REGISTERS_reg[3][18]  ( .G(n2296), .D(N3353), .Q(\REGISTERS[3][18] )
         );
  DLH_X1 \REGISTERS_reg[3][17]  ( .G(n2296), .D(N3351), .Q(\REGISTERS[3][17] )
         );
  DLH_X1 \REGISTERS_reg[3][16]  ( .G(n2296), .D(N3349), .Q(\REGISTERS[3][16] )
         );
  DLH_X1 \REGISTERS_reg[3][15]  ( .G(n2296), .D(N3347), .Q(\REGISTERS[3][15] )
         );
  DLH_X1 \REGISTERS_reg[3][14]  ( .G(n2296), .D(N3345), .Q(\REGISTERS[3][14] )
         );
  DLH_X1 \REGISTERS_reg[3][13]  ( .G(n2296), .D(N3343), .Q(\REGISTERS[3][13] )
         );
  DLH_X1 \REGISTERS_reg[3][12]  ( .G(n2296), .D(N3341), .Q(\REGISTERS[3][12] )
         );
  DLH_X1 \REGISTERS_reg[3][11]  ( .G(n2296), .D(N3339), .Q(\REGISTERS[3][11] )
         );
  DLH_X1 \REGISTERS_reg[3][10]  ( .G(n2296), .D(N3337), .Q(\REGISTERS[3][10] )
         );
  DLH_X1 \REGISTERS_reg[3][9]  ( .G(n2296), .D(N3335), .Q(\REGISTERS[3][9] )
         );
  DLH_X1 \REGISTERS_reg[3][8]  ( .G(n2296), .D(N3333), .Q(\REGISTERS[3][8] )
         );
  DLH_X1 \REGISTERS_reg[3][7]  ( .G(n2296), .D(N3331), .Q(\REGISTERS[3][7] )
         );
  DLH_X1 \REGISTERS_reg[3][6]  ( .G(n2296), .D(N3329), .Q(\REGISTERS[3][6] )
         );
  DLH_X1 \REGISTERS_reg[3][5]  ( .G(n2297), .D(N3327), .Q(\REGISTERS[3][5] )
         );
  DLH_X1 \REGISTERS_reg[3][4]  ( .G(n2297), .D(N3325), .Q(\REGISTERS[3][4] )
         );
  DLH_X1 \REGISTERS_reg[3][3]  ( .G(n2297), .D(N3323), .Q(\REGISTERS[3][3] )
         );
  DLH_X1 \REGISTERS_reg[3][2]  ( .G(n2297), .D(N3321), .Q(\REGISTERS[3][2] )
         );
  DLH_X1 \REGISTERS_reg[3][1]  ( .G(n2297), .D(N3319), .Q(\REGISTERS[3][1] )
         );
  DLH_X1 \REGISTERS_reg[3][0]  ( .G(n2297), .D(N3317), .Q(\REGISTERS[3][0] )
         );
  DLH_X1 \REGISTERS_reg[2][31]  ( .G(n2298), .D(n1948), .Q(\REGISTERS[2][31] )
         );
  DLH_X1 \REGISTERS_reg[2][30]  ( .G(n2298), .D(n1947), .Q(\REGISTERS[2][30] )
         );
  DLH_X1 \REGISTERS_reg[2][29]  ( .G(n2298), .D(n1946), .Q(\REGISTERS[2][29] )
         );
  DLH_X1 \REGISTERS_reg[2][28]  ( .G(n2298), .D(n1945), .Q(\REGISTERS[2][28] )
         );
  DLH_X1 \REGISTERS_reg[2][27]  ( .G(n2298), .D(n1944), .Q(\REGISTERS[2][27] )
         );
  DLH_X1 \REGISTERS_reg[2][26]  ( .G(n2298), .D(n1943), .Q(\REGISTERS[2][26] )
         );
  DLH_X1 \REGISTERS_reg[2][25]  ( .G(n2298), .D(n1942), .Q(\REGISTERS[2][25] )
         );
  DLH_X1 \REGISTERS_reg[2][24]  ( .G(n2298), .D(n1941), .Q(\REGISTERS[2][24] )
         );
  DLH_X1 \REGISTERS_reg[2][23]  ( .G(n2298), .D(n1940), .Q(\REGISTERS[2][23] )
         );
  DLH_X1 \REGISTERS_reg[2][22]  ( .G(n2298), .D(n1939), .Q(\REGISTERS[2][22] )
         );
  DLH_X1 \REGISTERS_reg[2][21]  ( .G(n2298), .D(n1938), .Q(\REGISTERS[2][21] )
         );
  DLH_X1 \REGISTERS_reg[2][20]  ( .G(n2298), .D(n1937), .Q(\REGISTERS[2][20] )
         );
  DLH_X1 \REGISTERS_reg[2][19]  ( .G(n2298), .D(n1936), .Q(\REGISTERS[2][19] )
         );
  DLH_X1 \REGISTERS_reg[2][18]  ( .G(n2299), .D(n1935), .Q(\REGISTERS[2][18] )
         );
  DLH_X1 \REGISTERS_reg[2][17]  ( .G(n2299), .D(n1934), .Q(\REGISTERS[2][17] )
         );
  DLH_X1 \REGISTERS_reg[2][16]  ( .G(n2299), .D(n1933), .Q(\REGISTERS[2][16] )
         );
  DLH_X1 \REGISTERS_reg[2][15]  ( .G(n2299), .D(n1932), .Q(\REGISTERS[2][15] )
         );
  DLH_X1 \REGISTERS_reg[2][14]  ( .G(n2299), .D(n1931), .Q(\REGISTERS[2][14] )
         );
  DLH_X1 \REGISTERS_reg[2][13]  ( .G(n2299), .D(n1930), .Q(\REGISTERS[2][13] )
         );
  DLH_X1 \REGISTERS_reg[2][12]  ( .G(n2299), .D(n1929), .Q(\REGISTERS[2][12] )
         );
  DLH_X1 \REGISTERS_reg[2][11]  ( .G(n2299), .D(n1928), .Q(\REGISTERS[2][11] )
         );
  DLH_X1 \REGISTERS_reg[2][10]  ( .G(n2299), .D(n1927), .Q(\REGISTERS[2][10] )
         );
  DLH_X1 \REGISTERS_reg[2][9]  ( .G(n2299), .D(n1926), .Q(\REGISTERS[2][9] )
         );
  DLH_X1 \REGISTERS_reg[2][8]  ( .G(n2299), .D(n1925), .Q(\REGISTERS[2][8] )
         );
  DLH_X1 \REGISTERS_reg[2][7]  ( .G(n2299), .D(n1924), .Q(\REGISTERS[2][7] )
         );
  DLH_X1 \REGISTERS_reg[2][6]  ( .G(n2299), .D(n1923), .Q(\REGISTERS[2][6] )
         );
  DLH_X1 \REGISTERS_reg[2][5]  ( .G(n2300), .D(n1922), .Q(\REGISTERS[2][5] )
         );
  DLH_X1 \REGISTERS_reg[2][4]  ( .G(n2300), .D(n1921), .Q(\REGISTERS[2][4] )
         );
  DLH_X1 \REGISTERS_reg[2][3]  ( .G(n2300), .D(n1920), .Q(\REGISTERS[2][3] )
         );
  DLH_X1 \REGISTERS_reg[2][2]  ( .G(n2300), .D(n1919), .Q(\REGISTERS[2][2] )
         );
  DLH_X1 \REGISTERS_reg[2][1]  ( .G(n2300), .D(n1918), .Q(\REGISTERS[2][1] )
         );
  DLH_X1 \REGISTERS_reg[2][0]  ( .G(n2300), .D(n1917), .Q(\REGISTERS[2][0] )
         );
  DLH_X1 \REGISTERS_reg[1][31]  ( .G(n2301), .D(N3379), .Q(\REGISTERS[1][31] )
         );
  DLH_X1 \REGISTERS_reg[1][30]  ( .G(n2301), .D(N3377), .Q(\REGISTERS[1][30] )
         );
  DLH_X1 \REGISTERS_reg[1][29]  ( .G(n2301), .D(N3375), .Q(\REGISTERS[1][29] )
         );
  DLH_X1 \REGISTERS_reg[1][28]  ( .G(n2301), .D(N3373), .Q(\REGISTERS[1][28] )
         );
  DLH_X1 \REGISTERS_reg[1][27]  ( .G(n2301), .D(N3371), .Q(\REGISTERS[1][27] )
         );
  DLH_X1 \REGISTERS_reg[1][26]  ( .G(n2301), .D(N3369), .Q(\REGISTERS[1][26] )
         );
  DLH_X1 \REGISTERS_reg[1][25]  ( .G(n2301), .D(N3367), .Q(\REGISTERS[1][25] )
         );
  DLH_X1 \REGISTERS_reg[1][24]  ( .G(n2301), .D(N3365), .Q(\REGISTERS[1][24] )
         );
  DLH_X1 \REGISTERS_reg[1][23]  ( .G(n2301), .D(N3363), .Q(\REGISTERS[1][23] )
         );
  DLH_X1 \REGISTERS_reg[1][22]  ( .G(n2301), .D(N3361), .Q(\REGISTERS[1][22] )
         );
  DLH_X1 \REGISTERS_reg[1][21]  ( .G(n2301), .D(N3359), .Q(\REGISTERS[1][21] )
         );
  DLH_X1 \REGISTERS_reg[1][20]  ( .G(n2301), .D(N3357), .Q(\REGISTERS[1][20] )
         );
  DLH_X1 \REGISTERS_reg[1][19]  ( .G(n2301), .D(N3355), .Q(\REGISTERS[1][19] )
         );
  DLH_X1 \REGISTERS_reg[1][18]  ( .G(n2302), .D(N3353), .Q(\REGISTERS[1][18] )
         );
  DLH_X1 \REGISTERS_reg[1][17]  ( .G(n2302), .D(N3351), .Q(\REGISTERS[1][17] )
         );
  DLH_X1 \REGISTERS_reg[1][16]  ( .G(n2302), .D(N3349), .Q(\REGISTERS[1][16] )
         );
  DLH_X1 \REGISTERS_reg[1][15]  ( .G(n2302), .D(N3347), .Q(\REGISTERS[1][15] )
         );
  DLH_X1 \REGISTERS_reg[1][14]  ( .G(n2302), .D(N3345), .Q(\REGISTERS[1][14] )
         );
  DLH_X1 \REGISTERS_reg[1][13]  ( .G(n2302), .D(N3343), .Q(\REGISTERS[1][13] )
         );
  DLH_X1 \REGISTERS_reg[1][12]  ( .G(n2302), .D(N3341), .Q(\REGISTERS[1][12] )
         );
  DLH_X1 \REGISTERS_reg[1][11]  ( .G(n2302), .D(N3339), .Q(\REGISTERS[1][11] )
         );
  DLH_X1 \REGISTERS_reg[1][10]  ( .G(n2302), .D(N3337), .Q(\REGISTERS[1][10] )
         );
  DLH_X1 \REGISTERS_reg[1][9]  ( .G(n2302), .D(N3335), .Q(\REGISTERS[1][9] )
         );
  DLH_X1 \REGISTERS_reg[1][8]  ( .G(n2302), .D(N3333), .Q(\REGISTERS[1][8] )
         );
  DLH_X1 \REGISTERS_reg[1][7]  ( .G(n2302), .D(N3331), .Q(\REGISTERS[1][7] )
         );
  DLH_X1 \REGISTERS_reg[1][6]  ( .G(n2302), .D(N3329), .Q(\REGISTERS[1][6] )
         );
  DLH_X1 \REGISTERS_reg[1][5]  ( .G(n2303), .D(N3327), .Q(\REGISTERS[1][5] )
         );
  DLH_X1 \REGISTERS_reg[1][4]  ( .G(n2303), .D(N3325), .Q(\REGISTERS[1][4] )
         );
  DLH_X1 \REGISTERS_reg[1][3]  ( .G(n2303), .D(N3323), .Q(\REGISTERS[1][3] )
         );
  DLH_X1 \REGISTERS_reg[1][2]  ( .G(n2303), .D(N3321), .Q(\REGISTERS[1][2] )
         );
  DLH_X1 \REGISTERS_reg[1][1]  ( .G(n2303), .D(N3319), .Q(\REGISTERS[1][1] )
         );
  DLH_X1 \REGISTERS_reg[1][0]  ( .G(n2303), .D(N3317), .Q(\REGISTERS[1][0] )
         );
  DLH_X1 \REGISTERS_reg[0][31]  ( .G(n2304), .D(n1948), .Q(\REGISTERS[0][31] )
         );
  DFF_X1 \DATA_OUT_1_reg[31]  ( .D(n2043), .CK(N1072), .Q(DATA_OUT_1[31]) );
  DLH_X1 \REGISTERS_reg[0][30]  ( .G(n2304), .D(n1947), .Q(\REGISTERS[0][30] )
         );
  DFF_X1 \DATA_OUT_1_reg[30]  ( .D(n2042), .CK(N1072), .Q(DATA_OUT_1[30]) );
  DLH_X1 \REGISTERS_reg[0][29]  ( .G(n2304), .D(n1946), .Q(\REGISTERS[0][29] )
         );
  DFF_X1 \DATA_OUT_1_reg[29]  ( .D(n2041), .CK(N1072), .Q(DATA_OUT_1[29]) );
  DLH_X1 \REGISTERS_reg[0][28]  ( .G(n2304), .D(n1945), .Q(\REGISTERS[0][28] )
         );
  DFF_X1 \DATA_OUT_1_reg[28]  ( .D(n2040), .CK(N1072), .Q(DATA_OUT_1[28]) );
  DLH_X1 \REGISTERS_reg[0][27]  ( .G(n2304), .D(n1944), .Q(\REGISTERS[0][27] )
         );
  DFF_X1 \DATA_OUT_1_reg[27]  ( .D(n2039), .CK(N1072), .Q(DATA_OUT_1[27]) );
  DLH_X1 \REGISTERS_reg[0][26]  ( .G(n2304), .D(n1943), .Q(\REGISTERS[0][26] )
         );
  DFF_X1 \DATA_OUT_1_reg[26]  ( .D(n2038), .CK(N1072), .Q(DATA_OUT_1[26]) );
  DLH_X1 \REGISTERS_reg[0][25]  ( .G(n2304), .D(n1942), .Q(\REGISTERS[0][25] )
         );
  DFF_X1 \DATA_OUT_1_reg[25]  ( .D(n2037), .CK(N1072), .Q(DATA_OUT_1[25]) );
  DLH_X1 \REGISTERS_reg[0][24]  ( .G(n2304), .D(n1941), .Q(\REGISTERS[0][24] )
         );
  DFF_X1 \DATA_OUT_1_reg[24]  ( .D(n2036), .CK(N1072), .Q(DATA_OUT_1[24]) );
  DLH_X1 \REGISTERS_reg[0][23]  ( .G(n2304), .D(n1940), .Q(\REGISTERS[0][23] )
         );
  DFF_X1 \DATA_OUT_1_reg[23]  ( .D(n2035), .CK(N1072), .Q(DATA_OUT_1[23]) );
  DLH_X1 \REGISTERS_reg[0][22]  ( .G(n2304), .D(n1939), .Q(\REGISTERS[0][22] )
         );
  DFF_X1 \DATA_OUT_1_reg[22]  ( .D(n2034), .CK(N1072), .Q(DATA_OUT_1[22]) );
  DLH_X1 \REGISTERS_reg[0][21]  ( .G(n2304), .D(n1938), .Q(\REGISTERS[0][21] )
         );
  DFF_X1 \DATA_OUT_1_reg[21]  ( .D(n2033), .CK(N1072), .Q(DATA_OUT_1[21]) );
  DLH_X1 \REGISTERS_reg[0][20]  ( .G(n2304), .D(n1937), .Q(\REGISTERS[0][20] )
         );
  DFF_X1 \DATA_OUT_1_reg[20]  ( .D(n2032), .CK(N1072), .Q(DATA_OUT_1[20]) );
  DLH_X1 \REGISTERS_reg[0][19]  ( .G(n2304), .D(n1936), .Q(\REGISTERS[0][19] )
         );
  DFF_X1 \DATA_OUT_1_reg[19]  ( .D(n2031), .CK(N1072), .Q(DATA_OUT_1[19]) );
  DLH_X1 \REGISTERS_reg[0][18]  ( .G(n2305), .D(n1935), .Q(\REGISTERS[0][18] )
         );
  DFF_X1 \DATA_OUT_1_reg[18]  ( .D(n2030), .CK(N1072), .Q(DATA_OUT_1[18]) );
  DLH_X1 \REGISTERS_reg[0][17]  ( .G(n2305), .D(n1934), .Q(\REGISTERS[0][17] )
         );
  DFF_X1 \DATA_OUT_1_reg[17]  ( .D(n2029), .CK(N1072), .Q(DATA_OUT_1[17]) );
  DLH_X1 \REGISTERS_reg[0][16]  ( .G(n2305), .D(n1933), .Q(\REGISTERS[0][16] )
         );
  DFF_X1 \DATA_OUT_1_reg[16]  ( .D(n2028), .CK(N1072), .Q(DATA_OUT_1[16]) );
  DLH_X1 \REGISTERS_reg[0][15]  ( .G(n2305), .D(n1932), .Q(\REGISTERS[0][15] )
         );
  DFF_X1 \DATA_OUT_1_reg[15]  ( .D(n2027), .CK(N1072), .Q(DATA_OUT_1[15]) );
  DLH_X1 \REGISTERS_reg[0][14]  ( .G(n2305), .D(n1931), .Q(\REGISTERS[0][14] )
         );
  DFF_X1 \DATA_OUT_1_reg[14]  ( .D(n2026), .CK(N1072), .Q(DATA_OUT_1[14]) );
  DLH_X1 \REGISTERS_reg[0][13]  ( .G(n2305), .D(n1930), .Q(\REGISTERS[0][13] )
         );
  DFF_X1 \DATA_OUT_1_reg[13]  ( .D(n2025), .CK(N1072), .Q(DATA_OUT_1[13]) );
  DLH_X1 \REGISTERS_reg[0][12]  ( .G(n2305), .D(n1929), .Q(\REGISTERS[0][12] )
         );
  DFF_X1 \DATA_OUT_1_reg[12]  ( .D(n2024), .CK(N1072), .Q(DATA_OUT_1[12]) );
  DLH_X1 \REGISTERS_reg[0][11]  ( .G(n2305), .D(n1928), .Q(\REGISTERS[0][11] )
         );
  DFF_X1 \DATA_OUT_1_reg[11]  ( .D(n2023), .CK(N1072), .Q(DATA_OUT_1[11]) );
  DLH_X1 \REGISTERS_reg[0][10]  ( .G(n2305), .D(n1927), .Q(\REGISTERS[0][10] )
         );
  DFF_X1 \DATA_OUT_1_reg[10]  ( .D(n2022), .CK(N1072), .Q(DATA_OUT_1[10]) );
  DLH_X1 \REGISTERS_reg[0][9]  ( .G(n2305), .D(n1926), .Q(\REGISTERS[0][9] )
         );
  DFF_X1 \DATA_OUT_1_reg[9]  ( .D(n2021), .CK(N1072), .Q(DATA_OUT_1[9]) );
  DLH_X1 \REGISTERS_reg[0][8]  ( .G(n2305), .D(n1925), .Q(\REGISTERS[0][8] )
         );
  DFF_X1 \DATA_OUT_1_reg[8]  ( .D(n2020), .CK(N1072), .Q(DATA_OUT_1[8]) );
  DLH_X1 \REGISTERS_reg[0][7]  ( .G(n2305), .D(n1924), .Q(\REGISTERS[0][7] )
         );
  DFF_X1 \DATA_OUT_1_reg[7]  ( .D(n2019), .CK(N1072), .Q(DATA_OUT_1[7]) );
  DLH_X1 \REGISTERS_reg[0][6]  ( .G(n2305), .D(n1923), .Q(\REGISTERS[0][6] )
         );
  DFF_X1 \DATA_OUT_1_reg[6]  ( .D(n2018), .CK(N1072), .Q(DATA_OUT_1[6]) );
  DLH_X1 \REGISTERS_reg[0][5]  ( .G(n2306), .D(n1922), .Q(\REGISTERS[0][5] )
         );
  DFF_X1 \DATA_OUT_1_reg[5]  ( .D(n2017), .CK(N1072), .Q(DATA_OUT_1[5]) );
  DLH_X1 \REGISTERS_reg[0][4]  ( .G(n2306), .D(n1921), .Q(\REGISTERS[0][4] )
         );
  DFF_X1 \DATA_OUT_1_reg[4]  ( .D(n2016), .CK(N1072), .Q(DATA_OUT_1[4]) );
  DLH_X1 \REGISTERS_reg[0][3]  ( .G(n2306), .D(n1920), .Q(\REGISTERS[0][3] )
         );
  DFF_X1 \DATA_OUT_1_reg[3]  ( .D(n2015), .CK(N1072), .Q(DATA_OUT_1[3]) );
  DLH_X1 \REGISTERS_reg[0][2]  ( .G(n2306), .D(n1919), .Q(\REGISTERS[0][2] )
         );
  DFF_X1 \DATA_OUT_1_reg[2]  ( .D(n2014), .CK(N1072), .Q(DATA_OUT_1[2]) );
  DLH_X1 \REGISTERS_reg[0][1]  ( .G(n2306), .D(n1918), .Q(\REGISTERS[0][1] )
         );
  DFF_X1 \DATA_OUT_1_reg[1]  ( .D(n2013), .CK(N1072), .Q(DATA_OUT_1[1]) );
  DLH_X1 \REGISTERS_reg[0][0]  ( .G(n2306), .D(n1917), .Q(\REGISTERS[0][0] )
         );
  DFF_X1 \DATA_OUT_1_reg[0]  ( .D(n2012), .CK(N1072), .Q(DATA_OUT_1[0]) );
  DFF_X1 \DATA_OUT_2_reg[31]  ( .D(n2011), .CK(N1072), .Q(DATA_OUT_2[31]) );
  DFF_X1 \DATA_OUT_2_reg[30]  ( .D(n2010), .CK(N1072), .Q(DATA_OUT_2[30]) );
  DFF_X1 \DATA_OUT_2_reg[29]  ( .D(n2009), .CK(N1072), .Q(DATA_OUT_2[29]) );
  DFF_X1 \DATA_OUT_2_reg[28]  ( .D(n2008), .CK(N1072), .Q(DATA_OUT_2[28]) );
  DFF_X1 \DATA_OUT_2_reg[27]  ( .D(n2007), .CK(N1072), .Q(DATA_OUT_2[27]) );
  DFF_X1 \DATA_OUT_2_reg[26]  ( .D(n2006), .CK(N1072), .Q(DATA_OUT_2[26]) );
  DFF_X1 \DATA_OUT_2_reg[25]  ( .D(n2005), .CK(N1072), .Q(DATA_OUT_2[25]) );
  DFF_X1 \DATA_OUT_2_reg[24]  ( .D(n2004), .CK(N1072), .Q(DATA_OUT_2[24]) );
  DFF_X1 \DATA_OUT_2_reg[23]  ( .D(n2003), .CK(N1072), .Q(DATA_OUT_2[23]) );
  DFF_X1 \DATA_OUT_2_reg[22]  ( .D(n2002), .CK(N1072), .Q(DATA_OUT_2[22]) );
  DFF_X1 \DATA_OUT_2_reg[21]  ( .D(n2001), .CK(N1072), .Q(DATA_OUT_2[21]) );
  DFF_X1 \DATA_OUT_2_reg[20]  ( .D(n2000), .CK(N1072), .Q(DATA_OUT_2[20]) );
  DFF_X1 \DATA_OUT_2_reg[19]  ( .D(n1999), .CK(N1072), .Q(DATA_OUT_2[19]) );
  DFF_X1 \DATA_OUT_2_reg[18]  ( .D(n1998), .CK(N1072), .Q(DATA_OUT_2[18]) );
  DFF_X1 \DATA_OUT_2_reg[17]  ( .D(n1997), .CK(N1072), .Q(DATA_OUT_2[17]) );
  DFF_X1 \DATA_OUT_2_reg[16]  ( .D(n1996), .CK(N1072), .Q(DATA_OUT_2[16]) );
  DFF_X1 \DATA_OUT_2_reg[15]  ( .D(n1995), .CK(N1072), .Q(DATA_OUT_2[15]) );
  DFF_X1 \DATA_OUT_2_reg[14]  ( .D(n1994), .CK(N1072), .Q(DATA_OUT_2[14]) );
  DFF_X1 \DATA_OUT_2_reg[13]  ( .D(n1993), .CK(N1072), .Q(DATA_OUT_2[13]) );
  DFF_X1 \DATA_OUT_2_reg[12]  ( .D(n1992), .CK(N1072), .Q(DATA_OUT_2[12]) );
  DFF_X1 \DATA_OUT_2_reg[11]  ( .D(n1991), .CK(N1072), .Q(DATA_OUT_2[11]) );
  DFF_X1 \DATA_OUT_2_reg[10]  ( .D(n1990), .CK(N1072), .Q(DATA_OUT_2[10]) );
  DFF_X1 \DATA_OUT_2_reg[9]  ( .D(n1989), .CK(N1072), .Q(DATA_OUT_2[9]) );
  DFF_X1 \DATA_OUT_2_reg[8]  ( .D(n1988), .CK(N1072), .Q(DATA_OUT_2[8]) );
  DFF_X1 \DATA_OUT_2_reg[7]  ( .D(n1987), .CK(N1072), .Q(DATA_OUT_2[7]) );
  DFF_X1 \DATA_OUT_2_reg[6]  ( .D(n1986), .CK(N1072), .Q(DATA_OUT_2[6]) );
  DFF_X1 \DATA_OUT_2_reg[5]  ( .D(n1985), .CK(N1072), .Q(DATA_OUT_2[5]) );
  DFF_X1 \DATA_OUT_2_reg[4]  ( .D(n1984), .CK(N1072), .Q(DATA_OUT_2[4]) );
  DFF_X1 \DATA_OUT_2_reg[3]  ( .D(n1983), .CK(N1072), .Q(DATA_OUT_2[3]) );
  DFF_X1 \DATA_OUT_2_reg[2]  ( .D(n1982), .CK(N1072), .Q(DATA_OUT_2[2]) );
  DFF_X1 \DATA_OUT_2_reg[1]  ( .D(n1981), .CK(N1072), .Q(DATA_OUT_2[1]) );
  DFF_X1 \DATA_OUT_2_reg[0]  ( .D(n1980), .CK(N1072), .Q(DATA_OUT_2[0]) );
  NAND3_X1 U598 ( .A1(n1228), .A2(n2120), .A3(n1230), .ZN(n12) );
  NAND2_X1 U599 ( .A1(n1224), .A2(n1227), .ZN(n10) );
  NAND2_X1 U604 ( .A1(n1226), .A2(n1225), .ZN(n19) );
  NAND2_X1 U605 ( .A1(n1234), .A2(n1227), .ZN(n17) );
  NAND2_X1 U610 ( .A1(n1235), .A2(n1225), .ZN(n26) );
  NAND2_X1 U611 ( .A1(n1239), .A2(n1227), .ZN(n24) );
  NAND2_X1 U618 ( .A1(n1241), .A2(n1240), .ZN(n33) );
  NAND2_X1 U620 ( .A1(n1245), .A2(n1227), .ZN(n31) );
  NAND3_X1 U624 ( .A1(n2122), .A2(n1246), .A3(n1239), .ZN(n45) );
  NAND3_X1 U625 ( .A1(n1235), .A2(n2120), .A3(n1230), .ZN(n43) );
  NAND3_X1 U627 ( .A1(n1239), .A2(n2121), .A3(n1230), .ZN(n49) );
  NAND3_X1 U629 ( .A1(n2122), .A2(n1246), .A3(n1241), .ZN(n47) );
  NAND3_X1 U632 ( .A1(n1245), .A2(n2122), .A3(n1247), .ZN(n53) );
  NAND3_X1 U633 ( .A1(n1241), .A2(n2120), .A3(n1230), .ZN(n51) );
  NAND3_X1 U636 ( .A1(n1245), .A2(n2120), .A3(n1230), .ZN(n57) );
  NAND3_X1 U638 ( .A1(n1228), .A2(n2121), .A3(n1247), .ZN(n55) );
  NAND3_X1 U642 ( .A1(n1234), .A2(n2121), .A3(n1230), .ZN(n64) );
  NAND3_X1 U643 ( .A1(n1247), .A2(n2121), .A3(n1235), .ZN(n62) );
  NAND3_X1 U650 ( .A1(n1224), .A2(n2122), .A3(n1230), .ZN(n71) );
  NAND3_X1 U652 ( .A1(n1247), .A2(n2121), .A3(n1226), .ZN(n69) );
  NAND3_X1 U1878 ( .A1(n1875), .A2(n1957), .A3(n1877), .ZN(n1280) );
  NAND2_X1 U1880 ( .A1(n1871), .A2(n1874), .ZN(n1279) );
  NAND2_X1 U1886 ( .A1(n1873), .A2(n1872), .ZN(n1285) );
  NAND2_X1 U1888 ( .A1(n1879), .A2(n1874), .ZN(n1284) );
  NAND2_X1 U1894 ( .A1(n1880), .A2(n1872), .ZN(n1290) );
  NAND2_X1 U1896 ( .A1(n1882), .A2(n1874), .ZN(n1289) );
  NAND2_X1 U1904 ( .A1(n1884), .A2(n1883), .ZN(n1295) );
  NAND2_X1 U1907 ( .A1(n1886), .A2(n1874), .ZN(n1294) );
  NAND3_X1 U1912 ( .A1(n1959), .A2(n1887), .A3(n1882), .ZN(n1305) );
  NAND3_X1 U1914 ( .A1(n1880), .A2(n1957), .A3(n1877), .ZN(n1304) );
  NAND3_X1 U1917 ( .A1(n1882), .A2(n1958), .A3(n1877), .ZN(n1307) );
  NAND3_X1 U1920 ( .A1(n1959), .A2(n1887), .A3(n1884), .ZN(n1306) );
  NAND3_X1 U1924 ( .A1(n1886), .A2(n1959), .A3(n1888), .ZN(n1309) );
  NAND3_X1 U1926 ( .A1(n1884), .A2(n1957), .A3(n1877), .ZN(n1308) );
  NAND3_X1 U1930 ( .A1(n1886), .A2(n1957), .A3(n1877), .ZN(n1311) );
  NAND3_X1 U1933 ( .A1(n1875), .A2(n1958), .A3(n1888), .ZN(n1310) );
  NAND3_X1 U1938 ( .A1(n1879), .A2(n1958), .A3(n1877), .ZN(n1316) );
  NAND3_X1 U1940 ( .A1(n1888), .A2(n1958), .A3(n1880), .ZN(n1315) );
  NAND3_X1 U1948 ( .A1(n1871), .A2(n1959), .A3(n1877), .ZN(n1321) );
  NAND3_X1 U1951 ( .A1(n1888), .A2(n1958), .A3(n1873), .ZN(n1320) );
  NAND3_X1 U1959 ( .A1(EN), .A2(n1876), .A3(RD1), .ZN(n1318) );
  NAND3_X1 U2003 ( .A1(ADDR_WR[4]), .A2(ADDR_WR[3]), .A3(WR), .ZN(n1899) );
  NAND3_X1 U2012 ( .A1(ADDR_WR[4]), .A2(n1909), .A3(WR), .ZN(n1908) );
  NAND3_X1 U2021 ( .A1(ADDR_WR[3]), .A2(n1911), .A3(WR), .ZN(n1910) );
  NAND3_X1 U2023 ( .A1(ADDR_WR[1]), .A2(ADDR_WR[0]), .A3(ADDR_WR[2]), .ZN(
        n1900) );
  NAND3_X1 U2025 ( .A1(ADDR_WR[1]), .A2(n1913), .A3(ADDR_WR[2]), .ZN(n1901) );
  NAND3_X1 U2027 ( .A1(ADDR_WR[0]), .A2(n1914), .A3(ADDR_WR[2]), .ZN(n1902) );
  NAND3_X1 U2029 ( .A1(n1913), .A2(n1914), .A3(ADDR_WR[2]), .ZN(n1903) );
  NAND3_X1 U2031 ( .A1(ADDR_WR[0]), .A2(n1915), .A3(ADDR_WR[1]), .ZN(n1904) );
  NAND3_X1 U2033 ( .A1(n1913), .A2(n1915), .A3(ADDR_WR[1]), .ZN(n1905) );
  NAND3_X1 U2035 ( .A1(n1914), .A2(n1915), .A3(ADDR_WR[0]), .ZN(n1906) );
  NAND3_X1 U2038 ( .A1(n1909), .A2(n1911), .A3(WR), .ZN(n1912) );
  NAND3_X1 U2041 ( .A1(n1914), .A2(n1915), .A3(n1913), .ZN(n1907) );
  INV_X2 U2045 ( .A(CLK), .ZN(N1072) );
  NOR4_X2 U3 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .ZN(n5) );
  CLKBUF_X3 U4 ( .A(n23), .Z(n2187) );
  NOR4_X2 U5 ( .A1(n761), .A2(n762), .A3(n763), .A4(n764), .ZN(n760) );
  NOR4_X2 U6 ( .A1(n723), .A2(n724), .A3(n725), .A4(n726), .ZN(n722) );
  NOR4_X2 U7 ( .A1(n685), .A2(n686), .A3(n687), .A4(n688), .ZN(n684) );
  NOR4_X2 U8 ( .A1(n647), .A2(n648), .A3(n649), .A4(n650), .ZN(n646) );
  NOR4_X2 U9 ( .A1(n609), .A2(n610), .A3(n611), .A4(n612), .ZN(n608) );
  NOR4_X2 U10 ( .A1(n571), .A2(n572), .A3(n573), .A4(n574), .ZN(n570) );
  NOR4_X2 U11 ( .A1(n533), .A2(n534), .A3(n535), .A4(n536), .ZN(n532) );
  NOR4_X2 U12 ( .A1(n495), .A2(n496), .A3(n497), .A4(n498), .ZN(n494) );
  NOR4_X2 U13 ( .A1(n457), .A2(n458), .A3(n459), .A4(n460), .ZN(n456) );
  NOR4_X2 U14 ( .A1(n419), .A2(n420), .A3(n421), .A4(n422), .ZN(n418) );
  NOR4_X2 U15 ( .A1(n381), .A2(n382), .A3(n383), .A4(n384), .ZN(n380) );
  NOR4_X2 U16 ( .A1(n343), .A2(n344), .A3(n345), .A4(n346), .ZN(n342) );
  NOR4_X2 U17 ( .A1(n305), .A2(n306), .A3(n307), .A4(n308), .ZN(n304) );
  BUF_X8 U18 ( .A(n1298), .Z(n2066) );
  AND2_X2 U19 ( .A1(n1224), .A2(n1225), .ZN(n16) );
  NOR4_X2 U20 ( .A1(n267), .A2(n268), .A3(n269), .A4(n270), .ZN(n266) );
  AND2_X2 U21 ( .A1(n1875), .A2(n1872), .ZN(n1298) );
  BUF_X8 U22 ( .A(n37), .Z(n2165) );
  AND2_X2 U23 ( .A1(n1228), .A2(n1225), .ZN(n37) );
  AND2_X1 U24 ( .A1(n1227), .A2(n1228), .ZN(n38) );
  NOR3_X1 U25 ( .A1(ADDR_RD1[1]), .A2(ADDR_RD1[2]), .A3(n1318), .ZN(n1874) );
  NAND3_X1 U26 ( .A1(EN), .A2(n1), .A3(RD2), .ZN(n67) );
  AND2_X1 U27 ( .A1(n2120), .A2(n1246), .ZN(n1225) );
  AND2_X1 U28 ( .A1(n1957), .A2(n1887), .ZN(n1872) );
  CLKBUF_X1 U29 ( .A(n36), .Z(n2168) );
  CLKBUF_X1 U30 ( .A(n15), .Z(n2204) );
  CLKBUF_X1 U31 ( .A(n22), .Z(n2192) );
  CLKBUF_X1 U32 ( .A(n29), .Z(n2180) );
  CLKBUF_X1 U33 ( .A(n1282), .Z(n2105) );
  CLKBUF_X1 U34 ( .A(n1287), .Z(n2093) );
  CLKBUF_X1 U35 ( .A(n1292), .Z(n2081) );
  CLKBUF_X1 U36 ( .A(n10), .Z(n2210) );
  CLKBUF_X1 U37 ( .A(n1297), .Z(n2069) );
  CLKBUF_X1 U38 ( .A(n16), .Z(n2201) );
  CLKBUF_X1 U39 ( .A(n23), .Z(n2189) );
  CLKBUF_X1 U40 ( .A(n1279), .Z(n2111) );
  CLKBUF_X1 U41 ( .A(n1284), .Z(n2099) );
  CLKBUF_X1 U42 ( .A(n1289), .Z(n2087) );
  CLKBUF_X1 U43 ( .A(n38), .Z(n2164) );
  CLKBUF_X1 U44 ( .A(n1293), .Z(n2078) );
  CLKBUF_X1 U45 ( .A(n1283), .Z(n2102) );
  CLKBUF_X1 U46 ( .A(n1288), .Z(n2090) );
  CLKBUF_X1 U47 ( .A(n1299), .Z(n2065) );
  INV_X1 U48 ( .A(n1958), .ZN(n1956) );
  INV_X1 U49 ( .A(n1959), .ZN(n1955) );
  INV_X1 U50 ( .A(n2121), .ZN(n2119) );
  INV_X1 U51 ( .A(n2122), .ZN(n2118) );
  BUF_X1 U52 ( .A(N1394), .Z(n2305) );
  BUF_X1 U53 ( .A(N1394), .Z(n2304) );
  BUF_X1 U54 ( .A(N1394), .Z(n2306) );
  BUF_X1 U55 ( .A(n1304), .Z(n2060) );
  BUF_X1 U56 ( .A(n1308), .Z(n2048) );
  BUF_X1 U57 ( .A(n1315), .Z(n1966) );
  BUF_X1 U58 ( .A(n1320), .Z(n1952) );
  BUF_X1 U59 ( .A(n1304), .Z(n2061) );
  BUF_X1 U60 ( .A(n1308), .Z(n2049) );
  BUF_X1 U61 ( .A(n1315), .Z(n1967) );
  BUF_X1 U62 ( .A(n1320), .Z(n1953) );
  BUF_X1 U63 ( .A(n1306), .Z(n2054) );
  BUF_X1 U64 ( .A(n1310), .Z(n1978) );
  BUF_X1 U65 ( .A(n1306), .Z(n2055) );
  BUF_X1 U66 ( .A(n1310), .Z(n1979) );
  BUF_X1 U67 ( .A(n1307), .Z(n2051) );
  BUF_X1 U68 ( .A(n1311), .Z(n1975) );
  BUF_X1 U69 ( .A(n1316), .Z(n1963) );
  BUF_X1 U70 ( .A(n1321), .Z(n1949) );
  BUF_X1 U71 ( .A(n1307), .Z(n2052) );
  BUF_X1 U72 ( .A(n1311), .Z(n1976) );
  BUF_X1 U73 ( .A(n1316), .Z(n1964) );
  BUF_X1 U74 ( .A(n1321), .Z(n1950) );
  BUF_X1 U75 ( .A(n1305), .Z(n2057) );
  BUF_X1 U76 ( .A(n1309), .Z(n2045) );
  BUF_X1 U77 ( .A(n1305), .Z(n2058) );
  BUF_X1 U78 ( .A(n1309), .Z(n2046) );
  BUF_X1 U79 ( .A(n1280), .Z(n2106) );
  BUF_X1 U80 ( .A(n1280), .Z(n2107) );
  BUF_X1 U81 ( .A(n49), .Z(n2150) );
  BUF_X1 U82 ( .A(n57), .Z(n2138) );
  BUF_X1 U83 ( .A(n64), .Z(n2126) );
  BUF_X1 U84 ( .A(n71), .Z(n2112) );
  BUF_X1 U85 ( .A(n49), .Z(n2151) );
  BUF_X1 U86 ( .A(n57), .Z(n2139) );
  BUF_X1 U87 ( .A(n64), .Z(n2127) );
  BUF_X1 U88 ( .A(n71), .Z(n2113) );
  BUF_X1 U89 ( .A(n45), .Z(n2156) );
  BUF_X1 U90 ( .A(n53), .Z(n2144) );
  BUF_X1 U91 ( .A(n45), .Z(n2157) );
  BUF_X1 U92 ( .A(n53), .Z(n2145) );
  BUF_X1 U93 ( .A(n43), .Z(n2159) );
  BUF_X1 U94 ( .A(n51), .Z(n2147) );
  BUF_X1 U95 ( .A(n62), .Z(n2129) );
  BUF_X1 U96 ( .A(n69), .Z(n2115) );
  BUF_X1 U97 ( .A(n43), .Z(n2160) );
  BUF_X1 U98 ( .A(n51), .Z(n2148) );
  BUF_X1 U99 ( .A(n62), .Z(n2130) );
  BUF_X1 U100 ( .A(n69), .Z(n2116) );
  BUF_X1 U101 ( .A(n47), .Z(n2153) );
  BUF_X1 U102 ( .A(n55), .Z(n2141) );
  BUF_X1 U103 ( .A(n47), .Z(n2154) );
  BUF_X1 U104 ( .A(n55), .Z(n2142) );
  BUF_X1 U105 ( .A(n12), .Z(n2205) );
  BUF_X1 U106 ( .A(n12), .Z(n2206) );
  BUF_X1 U107 ( .A(n31), .Z(n2174) );
  BUF_X1 U108 ( .A(n17), .Z(n2198) );
  BUF_X1 U109 ( .A(n24), .Z(n2186) );
  BUF_X1 U110 ( .A(n60), .Z(n2134) );
  BUF_X1 U111 ( .A(n30), .Z(n2177) );
  BUF_X1 U112 ( .A(n1304), .Z(n2062) );
  BUF_X1 U113 ( .A(n1308), .Z(n2050) );
  BUF_X1 U114 ( .A(n1315), .Z(n1968) );
  BUF_X1 U115 ( .A(n1320), .Z(n1954) );
  BUF_X1 U116 ( .A(n1306), .Z(n2056) );
  BUF_X1 U117 ( .A(n1310), .Z(n2044) );
  BUF_X1 U118 ( .A(n1307), .Z(n2053) );
  BUF_X1 U119 ( .A(n1311), .Z(n1977) );
  BUF_X1 U120 ( .A(n1316), .Z(n1965) );
  BUF_X1 U121 ( .A(n1321), .Z(n1951) );
  BUF_X1 U122 ( .A(n1305), .Z(n2059) );
  BUF_X1 U123 ( .A(n1309), .Z(n2047) );
  BUF_X1 U124 ( .A(n1295), .Z(n2072) );
  BUF_X1 U125 ( .A(n1285), .Z(n2096) );
  BUF_X1 U126 ( .A(n1290), .Z(n2084) );
  BUF_X1 U127 ( .A(n1280), .Z(n2108) );
  BUF_X1 U128 ( .A(n1312), .Z(n1974) );
  BUF_X1 U129 ( .A(n1317), .Z(n1962) );
  BUF_X1 U130 ( .A(n1294), .Z(n2075) );
  BUF_X1 U131 ( .A(n49), .Z(n2152) );
  BUF_X1 U132 ( .A(n57), .Z(n2140) );
  BUF_X1 U133 ( .A(n64), .Z(n2128) );
  BUF_X1 U134 ( .A(n71), .Z(n2114) );
  BUF_X1 U135 ( .A(n45), .Z(n2158) );
  BUF_X1 U136 ( .A(n53), .Z(n2146) );
  BUF_X1 U137 ( .A(n43), .Z(n2161) );
  BUF_X1 U138 ( .A(n51), .Z(n2149) );
  BUF_X1 U139 ( .A(n62), .Z(n2131) );
  BUF_X1 U140 ( .A(n69), .Z(n2117) );
  BUF_X1 U141 ( .A(n47), .Z(n2155) );
  BUF_X1 U142 ( .A(n55), .Z(n2143) );
  BUF_X1 U143 ( .A(n1313), .Z(n1971) );
  BUF_X1 U144 ( .A(n59), .Z(n2137) );
  BUF_X1 U145 ( .A(n66), .Z(n2125) );
  BUF_X1 U146 ( .A(n33), .Z(n2171) );
  BUF_X1 U147 ( .A(n19), .Z(n2195) );
  BUF_X1 U148 ( .A(n26), .Z(n2183) );
  BUF_X1 U149 ( .A(n12), .Z(n2207) );
  BUF_X1 U150 ( .A(n10), .Z(n2208) );
  BUF_X1 U151 ( .A(n17), .Z(n2196) );
  BUF_X1 U152 ( .A(n24), .Z(n2184) );
  BUF_X1 U153 ( .A(n31), .Z(n2173) );
  BUF_X1 U154 ( .A(n10), .Z(n2209) );
  BUF_X1 U155 ( .A(n17), .Z(n2197) );
  BUF_X1 U156 ( .A(n24), .Z(n2185) );
  BUF_X1 U157 ( .A(n60), .Z(n2133) );
  BUF_X1 U158 ( .A(n60), .Z(n2132) );
  BUF_X1 U159 ( .A(n15), .Z(n2203) );
  BUF_X1 U160 ( .A(n22), .Z(n2191) );
  BUF_X1 U161 ( .A(n15), .Z(n2202) );
  BUF_X1 U162 ( .A(n22), .Z(n2190) );
  BUF_X1 U163 ( .A(n29), .Z(n2179) );
  BUF_X1 U164 ( .A(n29), .Z(n2178) );
  BUF_X1 U165 ( .A(n16), .Z(n2200) );
  BUF_X1 U166 ( .A(n23), .Z(n2188) );
  BUF_X1 U167 ( .A(n16), .Z(n2199) );
  BUF_X1 U168 ( .A(n30), .Z(n2176) );
  BUF_X1 U169 ( .A(n30), .Z(n2175) );
  BUF_X1 U170 ( .A(n31), .Z(n2172) );
  BUF_X1 U171 ( .A(n38), .Z(n2163) );
  BUF_X1 U172 ( .A(n38), .Z(n2162) );
  BUF_X1 U173 ( .A(n1285), .Z(n2094) );
  BUF_X1 U174 ( .A(n1290), .Z(n2082) );
  BUF_X1 U175 ( .A(n1295), .Z(n2071) );
  BUF_X1 U176 ( .A(n1285), .Z(n2095) );
  BUF_X1 U177 ( .A(n1290), .Z(n2083) );
  BUF_X1 U178 ( .A(n1312), .Z(n1973) );
  BUF_X1 U179 ( .A(n1317), .Z(n1961) );
  BUF_X1 U180 ( .A(n1312), .Z(n1972) );
  BUF_X1 U181 ( .A(n1317), .Z(n1960) );
  BUF_X1 U182 ( .A(n36), .Z(n2167) );
  BUF_X1 U183 ( .A(n36), .Z(n2166) );
  BUF_X1 U184 ( .A(n1279), .Z(n2109) );
  BUF_X1 U185 ( .A(n1284), .Z(n2097) );
  BUF_X1 U186 ( .A(n1289), .Z(n2085) );
  BUF_X1 U187 ( .A(n1294), .Z(n2074) );
  BUF_X1 U188 ( .A(n1279), .Z(n2110) );
  BUF_X1 U189 ( .A(n1284), .Z(n2098) );
  BUF_X1 U190 ( .A(n1289), .Z(n2086) );
  BUF_X1 U191 ( .A(n1295), .Z(n2070) );
  BUF_X1 U192 ( .A(n1297), .Z(n2068) );
  BUF_X1 U193 ( .A(n1297), .Z(n2067) );
  BUF_X1 U194 ( .A(n1313), .Z(n1970) );
  BUF_X1 U195 ( .A(n1313), .Z(n1969) );
  BUF_X1 U196 ( .A(n1282), .Z(n2104) );
  BUF_X1 U197 ( .A(n1287), .Z(n2092) );
  BUF_X1 U198 ( .A(n1282), .Z(n2103) );
  BUF_X1 U199 ( .A(n1287), .Z(n2091) );
  BUF_X1 U200 ( .A(n1292), .Z(n2080) );
  BUF_X1 U201 ( .A(n1292), .Z(n2079) );
  BUF_X1 U202 ( .A(n59), .Z(n2136) );
  BUF_X1 U203 ( .A(n66), .Z(n2124) );
  BUF_X1 U204 ( .A(n59), .Z(n2135) );
  BUF_X1 U205 ( .A(n66), .Z(n2123) );
  BUF_X1 U206 ( .A(n1294), .Z(n2073) );
  BUF_X1 U207 ( .A(n19), .Z(n2193) );
  BUF_X1 U208 ( .A(n26), .Z(n2181) );
  BUF_X1 U209 ( .A(n33), .Z(n2170) );
  BUF_X1 U210 ( .A(n19), .Z(n2194) );
  BUF_X1 U211 ( .A(n26), .Z(n2182) );
  BUF_X1 U212 ( .A(n1283), .Z(n2101) );
  BUF_X1 U213 ( .A(n1288), .Z(n2089) );
  BUF_X1 U214 ( .A(n1283), .Z(n2100) );
  BUF_X1 U215 ( .A(n1288), .Z(n2088) );
  BUF_X1 U216 ( .A(n1293), .Z(n2077) );
  BUF_X1 U217 ( .A(n1293), .Z(n2076) );
  BUF_X1 U218 ( .A(n1299), .Z(n2064) );
  BUF_X1 U219 ( .A(n1299), .Z(n2063) );
  BUF_X1 U220 ( .A(n33), .Z(n2169) );
  AND2_X1 U221 ( .A1(n1247), .A2(n2122), .ZN(n1240) );
  AND2_X1 U222 ( .A1(n1888), .A2(n1959), .ZN(n1883) );
  BUF_X1 U223 ( .A(n1916), .Z(n1) );
  BUF_X1 U224 ( .A(n1916), .Z(n1876) );
  BUF_X1 U225 ( .A(n1229), .Z(n1270) );
  BUF_X1 U226 ( .A(n1916), .Z(n1229) );
  OAI21_X1 U227 ( .B1(n1907), .B2(n1912), .A(n1876), .ZN(N1394) );
  BUF_X1 U228 ( .A(N2930), .Z(n2233) );
  BUF_X1 U229 ( .A(N2930), .Z(n2232) );
  BUF_X1 U230 ( .A(N2994), .Z(n2230) );
  BUF_X1 U231 ( .A(N2994), .Z(n2229) );
  BUF_X1 U232 ( .A(N3058), .Z(n2227) );
  BUF_X1 U233 ( .A(N3058), .Z(n2226) );
  BUF_X1 U234 ( .A(N3122), .Z(n2224) );
  BUF_X1 U235 ( .A(N3122), .Z(n2223) );
  BUF_X1 U236 ( .A(N3186), .Z(n2221) );
  BUF_X1 U237 ( .A(N3186), .Z(n2220) );
  BUF_X1 U238 ( .A(N3250), .Z(n2218) );
  BUF_X1 U239 ( .A(N3250), .Z(n2217) );
  BUF_X1 U240 ( .A(N3314), .Z(n2215) );
  BUF_X1 U241 ( .A(N3314), .Z(n2214) );
  BUF_X1 U242 ( .A(N3378), .Z(n2212) );
  BUF_X1 U243 ( .A(N3378), .Z(n2211) );
  BUF_X1 U244 ( .A(N1458), .Z(n2302) );
  BUF_X1 U245 ( .A(N1458), .Z(n2301) );
  BUF_X1 U246 ( .A(N1522), .Z(n2299) );
  BUF_X1 U247 ( .A(N1522), .Z(n2298) );
  BUF_X1 U248 ( .A(N1586), .Z(n2296) );
  BUF_X1 U249 ( .A(N1586), .Z(n2295) );
  BUF_X1 U250 ( .A(N1650), .Z(n2293) );
  BUF_X1 U251 ( .A(N1650), .Z(n2292) );
  BUF_X1 U252 ( .A(N1714), .Z(n2290) );
  BUF_X1 U253 ( .A(N1714), .Z(n2289) );
  BUF_X1 U254 ( .A(N1778), .Z(n2287) );
  BUF_X1 U255 ( .A(N1778), .Z(n2286) );
  BUF_X1 U256 ( .A(N1842), .Z(n2284) );
  BUF_X1 U257 ( .A(N1842), .Z(n2283) );
  BUF_X1 U258 ( .A(N1906), .Z(n2281) );
  BUF_X1 U259 ( .A(N1906), .Z(n2280) );
  BUF_X1 U260 ( .A(N1970), .Z(n2278) );
  BUF_X1 U261 ( .A(N1970), .Z(n2277) );
  BUF_X1 U262 ( .A(N2034), .Z(n2275) );
  BUF_X1 U263 ( .A(N2034), .Z(n2274) );
  BUF_X1 U264 ( .A(N2098), .Z(n2272) );
  BUF_X1 U265 ( .A(N2098), .Z(n2271) );
  BUF_X1 U266 ( .A(N2162), .Z(n2269) );
  BUF_X1 U267 ( .A(N2162), .Z(n2268) );
  BUF_X1 U268 ( .A(N2226), .Z(n2266) );
  BUF_X1 U269 ( .A(N2226), .Z(n2265) );
  BUF_X1 U270 ( .A(N2290), .Z(n2263) );
  BUF_X1 U271 ( .A(N2290), .Z(n2262) );
  BUF_X1 U272 ( .A(N2354), .Z(n2260) );
  BUF_X1 U273 ( .A(N2354), .Z(n2259) );
  BUF_X1 U274 ( .A(N2418), .Z(n2257) );
  BUF_X1 U275 ( .A(N2418), .Z(n2256) );
  BUF_X1 U276 ( .A(N2482), .Z(n2254) );
  BUF_X1 U277 ( .A(N2482), .Z(n2253) );
  BUF_X1 U278 ( .A(N2546), .Z(n2251) );
  BUF_X1 U279 ( .A(N2546), .Z(n2250) );
  BUF_X1 U280 ( .A(N2610), .Z(n2248) );
  BUF_X1 U281 ( .A(N2610), .Z(n2247) );
  BUF_X1 U282 ( .A(N2674), .Z(n2245) );
  BUF_X1 U283 ( .A(N2674), .Z(n2244) );
  BUF_X1 U284 ( .A(N2738), .Z(n2242) );
  BUF_X1 U285 ( .A(N2738), .Z(n2241) );
  BUF_X1 U286 ( .A(N2802), .Z(n2239) );
  BUF_X1 U287 ( .A(N2802), .Z(n2238) );
  BUF_X1 U288 ( .A(N2866), .Z(n2236) );
  BUF_X1 U289 ( .A(N2866), .Z(n2235) );
  BUF_X1 U290 ( .A(N2930), .Z(n2234) );
  BUF_X1 U291 ( .A(N2994), .Z(n2231) );
  BUF_X1 U292 ( .A(N3058), .Z(n2228) );
  BUF_X1 U293 ( .A(N3122), .Z(n2225) );
  BUF_X1 U294 ( .A(N3186), .Z(n2222) );
  BUF_X1 U295 ( .A(N3250), .Z(n2219) );
  BUF_X1 U296 ( .A(N3314), .Z(n2216) );
  BUF_X1 U297 ( .A(N3378), .Z(n2213) );
  BUF_X1 U298 ( .A(N1458), .Z(n2303) );
  BUF_X1 U299 ( .A(N1522), .Z(n2300) );
  BUF_X1 U300 ( .A(N1586), .Z(n2297) );
  BUF_X1 U301 ( .A(N1650), .Z(n2294) );
  BUF_X1 U302 ( .A(N1714), .Z(n2291) );
  BUF_X1 U303 ( .A(N1778), .Z(n2288) );
  BUF_X1 U304 ( .A(N1842), .Z(n2285) );
  BUF_X1 U305 ( .A(N1906), .Z(n2282) );
  BUF_X1 U306 ( .A(N1970), .Z(n2279) );
  BUF_X1 U307 ( .A(N2034), .Z(n2276) );
  BUF_X1 U308 ( .A(N2098), .Z(n2273) );
  BUF_X1 U309 ( .A(N2162), .Z(n2270) );
  BUF_X1 U310 ( .A(N2226), .Z(n2267) );
  BUF_X1 U311 ( .A(N2290), .Z(n2264) );
  BUF_X1 U312 ( .A(N2354), .Z(n2261) );
  BUF_X1 U313 ( .A(N2418), .Z(n2258) );
  BUF_X1 U314 ( .A(N2482), .Z(n2255) );
  BUF_X1 U315 ( .A(N2546), .Z(n2252) );
  BUF_X1 U316 ( .A(N2610), .Z(n2249) );
  BUF_X1 U317 ( .A(N2674), .Z(n2246) );
  BUF_X1 U318 ( .A(N2738), .Z(n2243) );
  BUF_X1 U319 ( .A(N2802), .Z(n2240) );
  BUF_X1 U320 ( .A(N2866), .Z(n2237) );
  NOR4_X1 U321 ( .A1(n1275), .A2(n1276), .A3(n1277), .A4(n1278), .ZN(n1274) );
  OAI221_X1 U322 ( .B1(n25), .B2(n2085), .C1(n27), .C2(n2082), .A(n1291), .ZN(
        n1276) );
  OAI221_X1 U323 ( .B1(n18), .B2(n2097), .C1(n20), .C2(n2094), .A(n1286), .ZN(
        n1277) );
  OAI221_X1 U324 ( .B1(n11), .B2(n2109), .C1(n13), .C2(n2106), .A(n1281), .ZN(
        n1278) );
  NOR4_X1 U325 ( .A1(n1326), .A2(n1327), .A3(n1328), .A4(n1329), .ZN(n1325) );
  OAI221_X1 U326 ( .B1(n87), .B2(n2085), .C1(n88), .C2(n2082), .A(n1332), .ZN(
        n1327) );
  OAI221_X1 U327 ( .B1(n84), .B2(n2097), .C1(n85), .C2(n2094), .A(n1331), .ZN(
        n1328) );
  OAI221_X1 U328 ( .B1(n81), .B2(n2109), .C1(n82), .C2(n2106), .A(n1330), .ZN(
        n1329) );
  NOR4_X1 U329 ( .A1(n1344), .A2(n1345), .A3(n1346), .A4(n1347), .ZN(n1343) );
  OAI221_X1 U330 ( .B1(n125), .B2(n2085), .C1(n126), .C2(n2082), .A(n1350), 
        .ZN(n1345) );
  OAI221_X1 U331 ( .B1(n122), .B2(n2097), .C1(n123), .C2(n2094), .A(n1349), 
        .ZN(n1346) );
  OAI221_X1 U332 ( .B1(n119), .B2(n2109), .C1(n120), .C2(n2106), .A(n1348), 
        .ZN(n1347) );
  NOR4_X1 U333 ( .A1(n1362), .A2(n1363), .A3(n1364), .A4(n1365), .ZN(n1361) );
  OAI221_X1 U334 ( .B1(n163), .B2(n2085), .C1(n164), .C2(n2082), .A(n1368), 
        .ZN(n1363) );
  OAI221_X1 U335 ( .B1(n160), .B2(n2097), .C1(n161), .C2(n2094), .A(n1367), 
        .ZN(n1364) );
  OAI221_X1 U336 ( .B1(n157), .B2(n2109), .C1(n158), .C2(n2106), .A(n1366), 
        .ZN(n1365) );
  NOR4_X1 U337 ( .A1(n1380), .A2(n1381), .A3(n1382), .A4(n1383), .ZN(n1379) );
  OAI221_X1 U338 ( .B1(n201), .B2(n2085), .C1(n202), .C2(n2082), .A(n1386), 
        .ZN(n1381) );
  OAI221_X1 U339 ( .B1(n198), .B2(n2097), .C1(n199), .C2(n2094), .A(n1385), 
        .ZN(n1382) );
  OAI221_X1 U340 ( .B1(n195), .B2(n2109), .C1(n196), .C2(n2106), .A(n1384), 
        .ZN(n1383) );
  NOR4_X1 U341 ( .A1(n1398), .A2(n1399), .A3(n1400), .A4(n1401), .ZN(n1397) );
  OAI221_X1 U342 ( .B1(n239), .B2(n2085), .C1(n240), .C2(n2082), .A(n1404), 
        .ZN(n1399) );
  OAI221_X1 U343 ( .B1(n236), .B2(n2097), .C1(n237), .C2(n2094), .A(n1403), 
        .ZN(n1400) );
  OAI221_X1 U344 ( .B1(n233), .B2(n2109), .C1(n234), .C2(n2106), .A(n1402), 
        .ZN(n1401) );
  NOR4_X1 U345 ( .A1(n1416), .A2(n1417), .A3(n1418), .A4(n1419), .ZN(n1415) );
  OAI221_X1 U346 ( .B1(n277), .B2(n2085), .C1(n278), .C2(n2082), .A(n1422), 
        .ZN(n1417) );
  OAI221_X1 U347 ( .B1(n274), .B2(n2097), .C1(n275), .C2(n2094), .A(n1421), 
        .ZN(n1418) );
  OAI221_X1 U348 ( .B1(n271), .B2(n2109), .C1(n272), .C2(n2106), .A(n1420), 
        .ZN(n1419) );
  NOR4_X1 U349 ( .A1(n1434), .A2(n1435), .A3(n1436), .A4(n1437), .ZN(n1433) );
  OAI221_X1 U350 ( .B1(n315), .B2(n2085), .C1(n316), .C2(n2082), .A(n1440), 
        .ZN(n1435) );
  OAI221_X1 U351 ( .B1(n312), .B2(n2097), .C1(n313), .C2(n2094), .A(n1439), 
        .ZN(n1436) );
  OAI221_X1 U352 ( .B1(n309), .B2(n2109), .C1(n310), .C2(n2106), .A(n1438), 
        .ZN(n1437) );
  NOR4_X1 U353 ( .A1(n1452), .A2(n1453), .A3(n1454), .A4(n1455), .ZN(n1451) );
  OAI221_X1 U354 ( .B1(n353), .B2(n2085), .C1(n354), .C2(n2082), .A(n1458), 
        .ZN(n1453) );
  OAI221_X1 U355 ( .B1(n350), .B2(n2097), .C1(n351), .C2(n2094), .A(n1457), 
        .ZN(n1454) );
  OAI221_X1 U356 ( .B1(n347), .B2(n2109), .C1(n348), .C2(n2106), .A(n1456), 
        .ZN(n1455) );
  NOR4_X1 U357 ( .A1(n1470), .A2(n1471), .A3(n1472), .A4(n1473), .ZN(n1469) );
  OAI221_X1 U358 ( .B1(n391), .B2(n2085), .C1(n392), .C2(n2082), .A(n1476), 
        .ZN(n1471) );
  OAI221_X1 U359 ( .B1(n388), .B2(n2097), .C1(n389), .C2(n2094), .A(n1475), 
        .ZN(n1472) );
  OAI221_X1 U360 ( .B1(n385), .B2(n2109), .C1(n386), .C2(n2106), .A(n1474), 
        .ZN(n1473) );
  NOR4_X1 U361 ( .A1(n1488), .A2(n1489), .A3(n1490), .A4(n1491), .ZN(n1487) );
  OAI221_X1 U362 ( .B1(n429), .B2(n2085), .C1(n430), .C2(n2082), .A(n1494), 
        .ZN(n1489) );
  OAI221_X1 U363 ( .B1(n426), .B2(n2097), .C1(n427), .C2(n2094), .A(n1493), 
        .ZN(n1490) );
  OAI221_X1 U364 ( .B1(n423), .B2(n2109), .C1(n424), .C2(n2106), .A(n1492), 
        .ZN(n1491) );
  NOR4_X1 U365 ( .A1(n1506), .A2(n1507), .A3(n1508), .A4(n1509), .ZN(n1505) );
  OAI221_X1 U366 ( .B1(n467), .B2(n2085), .C1(n468), .C2(n2082), .A(n1512), 
        .ZN(n1507) );
  OAI221_X1 U367 ( .B1(n464), .B2(n2097), .C1(n465), .C2(n2094), .A(n1511), 
        .ZN(n1508) );
  OAI221_X1 U368 ( .B1(n461), .B2(n2109), .C1(n462), .C2(n2106), .A(n1510), 
        .ZN(n1509) );
  NOR4_X1 U369 ( .A1(n1524), .A2(n1525), .A3(n1526), .A4(n1527), .ZN(n1523) );
  OAI221_X1 U370 ( .B1(n505), .B2(n2085), .C1(n506), .C2(n2082), .A(n1530), 
        .ZN(n1525) );
  OAI221_X1 U371 ( .B1(n502), .B2(n2097), .C1(n503), .C2(n2094), .A(n1529), 
        .ZN(n1526) );
  OAI221_X1 U372 ( .B1(n499), .B2(n2109), .C1(n500), .C2(n2106), .A(n1528), 
        .ZN(n1527) );
  NOR4_X1 U373 ( .A1(n1542), .A2(n1543), .A3(n1544), .A4(n1545), .ZN(n1541) );
  OAI221_X1 U374 ( .B1(n543), .B2(n2086), .C1(n544), .C2(n2083), .A(n1548), 
        .ZN(n1543) );
  OAI221_X1 U375 ( .B1(n540), .B2(n2098), .C1(n541), .C2(n2095), .A(n1547), 
        .ZN(n1544) );
  OAI221_X1 U376 ( .B1(n537), .B2(n2110), .C1(n538), .C2(n2107), .A(n1546), 
        .ZN(n1545) );
  NOR4_X1 U377 ( .A1(n1560), .A2(n1561), .A3(n1562), .A4(n1563), .ZN(n1559) );
  OAI221_X1 U378 ( .B1(n581), .B2(n2086), .C1(n582), .C2(n2083), .A(n1566), 
        .ZN(n1561) );
  OAI221_X1 U379 ( .B1(n578), .B2(n2098), .C1(n579), .C2(n2095), .A(n1565), 
        .ZN(n1562) );
  OAI221_X1 U380 ( .B1(n575), .B2(n2110), .C1(n576), .C2(n2107), .A(n1564), 
        .ZN(n1563) );
  NOR4_X1 U381 ( .A1(n1578), .A2(n1579), .A3(n1580), .A4(n1581), .ZN(n1577) );
  OAI221_X1 U382 ( .B1(n619), .B2(n2086), .C1(n620), .C2(n2083), .A(n1584), 
        .ZN(n1579) );
  OAI221_X1 U383 ( .B1(n616), .B2(n2098), .C1(n617), .C2(n2095), .A(n1583), 
        .ZN(n1580) );
  OAI221_X1 U384 ( .B1(n613), .B2(n2110), .C1(n614), .C2(n2107), .A(n1582), 
        .ZN(n1581) );
  NOR4_X1 U385 ( .A1(n1596), .A2(n1597), .A3(n1598), .A4(n1599), .ZN(n1595) );
  OAI221_X1 U386 ( .B1(n657), .B2(n2086), .C1(n658), .C2(n2083), .A(n1602), 
        .ZN(n1597) );
  OAI221_X1 U387 ( .B1(n654), .B2(n2098), .C1(n655), .C2(n2095), .A(n1601), 
        .ZN(n1598) );
  OAI221_X1 U388 ( .B1(n651), .B2(n2110), .C1(n652), .C2(n2107), .A(n1600), 
        .ZN(n1599) );
  NOR4_X1 U389 ( .A1(n1614), .A2(n1615), .A3(n1616), .A4(n1617), .ZN(n1613) );
  OAI221_X1 U390 ( .B1(n695), .B2(n2086), .C1(n696), .C2(n2083), .A(n1620), 
        .ZN(n1615) );
  OAI221_X1 U391 ( .B1(n692), .B2(n2098), .C1(n693), .C2(n2095), .A(n1619), 
        .ZN(n1616) );
  OAI221_X1 U392 ( .B1(n689), .B2(n2110), .C1(n690), .C2(n2107), .A(n1618), 
        .ZN(n1617) );
  NOR4_X1 U393 ( .A1(n1632), .A2(n1633), .A3(n1634), .A4(n1635), .ZN(n1631) );
  OAI221_X1 U394 ( .B1(n733), .B2(n2086), .C1(n734), .C2(n2083), .A(n1638), 
        .ZN(n1633) );
  OAI221_X1 U395 ( .B1(n730), .B2(n2098), .C1(n731), .C2(n2095), .A(n1637), 
        .ZN(n1634) );
  OAI221_X1 U396 ( .B1(n727), .B2(n2110), .C1(n728), .C2(n2107), .A(n1636), 
        .ZN(n1635) );
  NOR4_X1 U397 ( .A1(n1650), .A2(n1651), .A3(n1652), .A4(n1653), .ZN(n1649) );
  OAI221_X1 U398 ( .B1(n771), .B2(n2086), .C1(n772), .C2(n2083), .A(n1656), 
        .ZN(n1651) );
  OAI221_X1 U399 ( .B1(n768), .B2(n2098), .C1(n769), .C2(n2095), .A(n1655), 
        .ZN(n1652) );
  OAI221_X1 U400 ( .B1(n765), .B2(n2110), .C1(n766), .C2(n2107), .A(n1654), 
        .ZN(n1653) );
  NOR4_X1 U401 ( .A1(n1668), .A2(n1669), .A3(n1670), .A4(n1671), .ZN(n1667) );
  OAI221_X1 U402 ( .B1(n809), .B2(n2086), .C1(n810), .C2(n2083), .A(n1674), 
        .ZN(n1669) );
  OAI221_X1 U403 ( .B1(n806), .B2(n2098), .C1(n807), .C2(n2095), .A(n1673), 
        .ZN(n1670) );
  OAI221_X1 U404 ( .B1(n803), .B2(n2110), .C1(n804), .C2(n2107), .A(n1672), 
        .ZN(n1671) );
  NOR4_X1 U405 ( .A1(n1686), .A2(n1687), .A3(n1688), .A4(n1689), .ZN(n1685) );
  OAI221_X1 U406 ( .B1(n847), .B2(n2086), .C1(n848), .C2(n2083), .A(n1692), 
        .ZN(n1687) );
  OAI221_X1 U407 ( .B1(n844), .B2(n2098), .C1(n845), .C2(n2095), .A(n1691), 
        .ZN(n1688) );
  OAI221_X1 U408 ( .B1(n841), .B2(n2110), .C1(n842), .C2(n2107), .A(n1690), 
        .ZN(n1689) );
  NOR4_X1 U409 ( .A1(n1704), .A2(n1705), .A3(n1706), .A4(n1707), .ZN(n1703) );
  OAI221_X1 U410 ( .B1(n885), .B2(n2086), .C1(n886), .C2(n2083), .A(n1710), 
        .ZN(n1705) );
  OAI221_X1 U411 ( .B1(n882), .B2(n2098), .C1(n883), .C2(n2095), .A(n1709), 
        .ZN(n1706) );
  OAI221_X1 U412 ( .B1(n879), .B2(n2110), .C1(n880), .C2(n2107), .A(n1708), 
        .ZN(n1707) );
  NOR4_X1 U413 ( .A1(n1722), .A2(n1723), .A3(n1724), .A4(n1725), .ZN(n1721) );
  OAI221_X1 U414 ( .B1(n923), .B2(n2086), .C1(n924), .C2(n2083), .A(n1728), 
        .ZN(n1723) );
  OAI221_X1 U415 ( .B1(n920), .B2(n2098), .C1(n921), .C2(n2095), .A(n1727), 
        .ZN(n1724) );
  OAI221_X1 U416 ( .B1(n917), .B2(n2110), .C1(n918), .C2(n2107), .A(n1726), 
        .ZN(n1725) );
  NOR4_X1 U417 ( .A1(n1740), .A2(n1741), .A3(n1742), .A4(n1743), .ZN(n1739) );
  OAI221_X1 U418 ( .B1(n961), .B2(n2086), .C1(n962), .C2(n2083), .A(n1746), 
        .ZN(n1741) );
  OAI221_X1 U419 ( .B1(n958), .B2(n2098), .C1(n959), .C2(n2095), .A(n1745), 
        .ZN(n1742) );
  OAI221_X1 U420 ( .B1(n955), .B2(n2110), .C1(n956), .C2(n2107), .A(n1744), 
        .ZN(n1743) );
  NOR4_X1 U421 ( .A1(n1758), .A2(n1759), .A3(n1760), .A4(n1761), .ZN(n1757) );
  OAI221_X1 U422 ( .B1(n999), .B2(n2086), .C1(n1000), .C2(n2083), .A(n1764), 
        .ZN(n1759) );
  OAI221_X1 U423 ( .B1(n996), .B2(n2098), .C1(n997), .C2(n2095), .A(n1763), 
        .ZN(n1760) );
  OAI221_X1 U424 ( .B1(n993), .B2(n2110), .C1(n994), .C2(n2107), .A(n1762), 
        .ZN(n1761) );
  NOR4_X1 U425 ( .A1(n77), .A2(n78), .A3(n79), .A4(n80), .ZN(n76) );
  OAI221_X1 U426 ( .B1(n2184), .B2(n87), .C1(n2181), .C2(n88), .A(n89), .ZN(
        n78) );
  OAI221_X1 U427 ( .B1(n2196), .B2(n84), .C1(n2193), .C2(n85), .A(n86), .ZN(
        n79) );
  OAI221_X1 U428 ( .B1(n2208), .B2(n81), .C1(n2205), .C2(n82), .A(n83), .ZN(
        n80) );
  NOR4_X1 U429 ( .A1(n115), .A2(n116), .A3(n117), .A4(n118), .ZN(n114) );
  OAI221_X1 U430 ( .B1(n2184), .B2(n125), .C1(n2181), .C2(n126), .A(n127), 
        .ZN(n116) );
  OAI221_X1 U431 ( .B1(n2196), .B2(n122), .C1(n2193), .C2(n123), .A(n124), 
        .ZN(n117) );
  OAI221_X1 U432 ( .B1(n2208), .B2(n119), .C1(n2205), .C2(n120), .A(n121), 
        .ZN(n118) );
  NOR4_X1 U433 ( .A1(n153), .A2(n154), .A3(n155), .A4(n156), .ZN(n152) );
  OAI221_X1 U434 ( .B1(n2184), .B2(n163), .C1(n2181), .C2(n164), .A(n165), 
        .ZN(n154) );
  OAI221_X1 U435 ( .B1(n2196), .B2(n160), .C1(n2193), .C2(n161), .A(n162), 
        .ZN(n155) );
  OAI221_X1 U436 ( .B1(n2208), .B2(n157), .C1(n2205), .C2(n158), .A(n159), 
        .ZN(n156) );
  NOR4_X1 U437 ( .A1(n191), .A2(n192), .A3(n193), .A4(n194), .ZN(n190) );
  OAI221_X1 U438 ( .B1(n2184), .B2(n201), .C1(n2181), .C2(n202), .A(n203), 
        .ZN(n192) );
  OAI221_X1 U439 ( .B1(n2196), .B2(n198), .C1(n2193), .C2(n199), .A(n200), 
        .ZN(n193) );
  OAI221_X1 U440 ( .B1(n2208), .B2(n195), .C1(n2205), .C2(n196), .A(n197), 
        .ZN(n194) );
  NOR4_X1 U441 ( .A1(n229), .A2(n230), .A3(n231), .A4(n232), .ZN(n228) );
  OAI221_X1 U442 ( .B1(n2184), .B2(n239), .C1(n2181), .C2(n240), .A(n241), 
        .ZN(n230) );
  OAI221_X1 U443 ( .B1(n2196), .B2(n236), .C1(n2193), .C2(n237), .A(n238), 
        .ZN(n231) );
  OAI221_X1 U444 ( .B1(n2208), .B2(n233), .C1(n2205), .C2(n234), .A(n235), 
        .ZN(n232) );
  OAI221_X1 U445 ( .B1(n2184), .B2(n277), .C1(n2181), .C2(n278), .A(n279), 
        .ZN(n268) );
  OAI221_X1 U446 ( .B1(n2196), .B2(n274), .C1(n2193), .C2(n275), .A(n276), 
        .ZN(n269) );
  OAI221_X1 U447 ( .B1(n2208), .B2(n271), .C1(n2205), .C2(n272), .A(n273), 
        .ZN(n270) );
  OAI221_X1 U448 ( .B1(n2184), .B2(n315), .C1(n2181), .C2(n316), .A(n317), 
        .ZN(n306) );
  OAI221_X1 U449 ( .B1(n2196), .B2(n312), .C1(n2193), .C2(n313), .A(n314), 
        .ZN(n307) );
  OAI221_X1 U450 ( .B1(n2208), .B2(n309), .C1(n2205), .C2(n310), .A(n311), 
        .ZN(n308) );
  OAI221_X1 U451 ( .B1(n2184), .B2(n353), .C1(n2181), .C2(n354), .A(n355), 
        .ZN(n344) );
  OAI221_X1 U452 ( .B1(n2196), .B2(n350), .C1(n2193), .C2(n351), .A(n352), 
        .ZN(n345) );
  OAI221_X1 U453 ( .B1(n2208), .B2(n347), .C1(n2205), .C2(n348), .A(n349), 
        .ZN(n346) );
  OAI221_X1 U454 ( .B1(n2184), .B2(n391), .C1(n2181), .C2(n392), .A(n393), 
        .ZN(n382) );
  OAI221_X1 U455 ( .B1(n2196), .B2(n388), .C1(n2193), .C2(n389), .A(n390), 
        .ZN(n383) );
  OAI221_X1 U456 ( .B1(n2208), .B2(n385), .C1(n2205), .C2(n386), .A(n387), 
        .ZN(n384) );
  OAI221_X1 U457 ( .B1(n2184), .B2(n429), .C1(n2181), .C2(n430), .A(n431), 
        .ZN(n420) );
  OAI221_X1 U458 ( .B1(n2196), .B2(n426), .C1(n2193), .C2(n427), .A(n428), 
        .ZN(n421) );
  OAI221_X1 U459 ( .B1(n2208), .B2(n423), .C1(n2205), .C2(n424), .A(n425), 
        .ZN(n422) );
  OAI221_X1 U460 ( .B1(n2184), .B2(n467), .C1(n2181), .C2(n468), .A(n469), 
        .ZN(n458) );
  OAI221_X1 U461 ( .B1(n2196), .B2(n464), .C1(n2193), .C2(n465), .A(n466), 
        .ZN(n459) );
  OAI221_X1 U462 ( .B1(n2208), .B2(n461), .C1(n2205), .C2(n462), .A(n463), 
        .ZN(n460) );
  OAI221_X1 U463 ( .B1(n2184), .B2(n505), .C1(n2181), .C2(n506), .A(n507), 
        .ZN(n496) );
  OAI221_X1 U464 ( .B1(n2196), .B2(n502), .C1(n2193), .C2(n503), .A(n504), 
        .ZN(n497) );
  OAI221_X1 U465 ( .B1(n2208), .B2(n499), .C1(n2205), .C2(n500), .A(n501), 
        .ZN(n498) );
  OAI221_X1 U466 ( .B1(n2185), .B2(n543), .C1(n2182), .C2(n544), .A(n545), 
        .ZN(n534) );
  OAI221_X1 U467 ( .B1(n2197), .B2(n540), .C1(n2194), .C2(n541), .A(n542), 
        .ZN(n535) );
  OAI221_X1 U468 ( .B1(n2209), .B2(n537), .C1(n2206), .C2(n538), .A(n539), 
        .ZN(n536) );
  OAI221_X1 U469 ( .B1(n2185), .B2(n581), .C1(n2182), .C2(n582), .A(n583), 
        .ZN(n572) );
  OAI221_X1 U470 ( .B1(n2197), .B2(n578), .C1(n2194), .C2(n579), .A(n580), 
        .ZN(n573) );
  OAI221_X1 U471 ( .B1(n2209), .B2(n575), .C1(n2206), .C2(n576), .A(n577), 
        .ZN(n574) );
  OAI221_X1 U472 ( .B1(n2185), .B2(n619), .C1(n2182), .C2(n620), .A(n621), 
        .ZN(n610) );
  OAI221_X1 U473 ( .B1(n2197), .B2(n616), .C1(n2194), .C2(n617), .A(n618), 
        .ZN(n611) );
  OAI221_X1 U474 ( .B1(n2209), .B2(n613), .C1(n2206), .C2(n614), .A(n615), 
        .ZN(n612) );
  OAI221_X1 U475 ( .B1(n2185), .B2(n657), .C1(n2182), .C2(n658), .A(n659), 
        .ZN(n648) );
  OAI221_X1 U476 ( .B1(n2197), .B2(n654), .C1(n2194), .C2(n655), .A(n656), 
        .ZN(n649) );
  OAI221_X1 U477 ( .B1(n2209), .B2(n651), .C1(n2206), .C2(n652), .A(n653), 
        .ZN(n650) );
  OAI221_X1 U478 ( .B1(n2185), .B2(n695), .C1(n2182), .C2(n696), .A(n697), 
        .ZN(n686) );
  OAI221_X1 U479 ( .B1(n2197), .B2(n692), .C1(n2194), .C2(n693), .A(n694), 
        .ZN(n687) );
  OAI221_X1 U480 ( .B1(n2209), .B2(n689), .C1(n2206), .C2(n690), .A(n691), 
        .ZN(n688) );
  OAI221_X1 U481 ( .B1(n2185), .B2(n733), .C1(n2182), .C2(n734), .A(n735), 
        .ZN(n724) );
  OAI221_X1 U482 ( .B1(n2197), .B2(n730), .C1(n2194), .C2(n731), .A(n732), 
        .ZN(n725) );
  OAI221_X1 U483 ( .B1(n2209), .B2(n727), .C1(n2206), .C2(n728), .A(n729), 
        .ZN(n726) );
  OAI221_X1 U484 ( .B1(n2185), .B2(n771), .C1(n2182), .C2(n772), .A(n773), 
        .ZN(n762) );
  OAI221_X1 U485 ( .B1(n2197), .B2(n768), .C1(n2194), .C2(n769), .A(n770), 
        .ZN(n763) );
  OAI221_X1 U486 ( .B1(n2209), .B2(n765), .C1(n2206), .C2(n766), .A(n767), 
        .ZN(n764) );
  NOR4_X1 U487 ( .A1(n799), .A2(n800), .A3(n801), .A4(n802), .ZN(n798) );
  OAI221_X1 U488 ( .B1(n2185), .B2(n809), .C1(n2182), .C2(n810), .A(n811), 
        .ZN(n800) );
  OAI221_X1 U489 ( .B1(n2197), .B2(n806), .C1(n2194), .C2(n807), .A(n808), 
        .ZN(n801) );
  OAI221_X1 U490 ( .B1(n2209), .B2(n803), .C1(n2206), .C2(n804), .A(n805), 
        .ZN(n802) );
  NOR4_X1 U491 ( .A1(n837), .A2(n838), .A3(n839), .A4(n840), .ZN(n836) );
  OAI221_X1 U492 ( .B1(n2185), .B2(n847), .C1(n2182), .C2(n848), .A(n849), 
        .ZN(n838) );
  OAI221_X1 U493 ( .B1(n2197), .B2(n844), .C1(n2194), .C2(n845), .A(n846), 
        .ZN(n839) );
  OAI221_X1 U494 ( .B1(n2209), .B2(n841), .C1(n2206), .C2(n842), .A(n843), 
        .ZN(n840) );
  NOR4_X1 U495 ( .A1(n875), .A2(n876), .A3(n877), .A4(n878), .ZN(n874) );
  OAI221_X1 U496 ( .B1(n2185), .B2(n885), .C1(n2182), .C2(n886), .A(n887), 
        .ZN(n876) );
  OAI221_X1 U497 ( .B1(n2197), .B2(n882), .C1(n2194), .C2(n883), .A(n884), 
        .ZN(n877) );
  OAI221_X1 U498 ( .B1(n2209), .B2(n879), .C1(n2206), .C2(n880), .A(n881), 
        .ZN(n878) );
  NOR4_X1 U499 ( .A1(n913), .A2(n914), .A3(n915), .A4(n916), .ZN(n912) );
  OAI221_X1 U500 ( .B1(n2185), .B2(n923), .C1(n2182), .C2(n924), .A(n925), 
        .ZN(n914) );
  OAI221_X1 U501 ( .B1(n2197), .B2(n920), .C1(n2194), .C2(n921), .A(n922), 
        .ZN(n915) );
  OAI221_X1 U502 ( .B1(n2209), .B2(n917), .C1(n2206), .C2(n918), .A(n919), 
        .ZN(n916) );
  NOR4_X1 U503 ( .A1(n951), .A2(n952), .A3(n953), .A4(n954), .ZN(n950) );
  OAI221_X1 U504 ( .B1(n2185), .B2(n961), .C1(n2182), .C2(n962), .A(n963), 
        .ZN(n952) );
  OAI221_X1 U505 ( .B1(n2197), .B2(n958), .C1(n2194), .C2(n959), .A(n960), 
        .ZN(n953) );
  OAI221_X1 U506 ( .B1(n2209), .B2(n955), .C1(n2206), .C2(n956), .A(n957), 
        .ZN(n954) );
  NOR4_X1 U507 ( .A1(n989), .A2(n990), .A3(n991), .A4(n992), .ZN(n988) );
  OAI221_X1 U508 ( .B1(n2185), .B2(n999), .C1(n2182), .C2(n1000), .A(n1001), 
        .ZN(n990) );
  OAI221_X1 U509 ( .B1(n2197), .B2(n996), .C1(n2194), .C2(n997), .A(n998), 
        .ZN(n991) );
  OAI221_X1 U510 ( .B1(n2209), .B2(n993), .C1(n2206), .C2(n994), .A(n995), 
        .ZN(n992) );
  NOR4_X1 U511 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1026) );
  OAI221_X1 U512 ( .B1(n2186), .B2(n1037), .C1(n2183), .C2(n1038), .A(n1039), 
        .ZN(n1028) );
  OAI221_X1 U513 ( .B1(n2198), .B2(n1034), .C1(n2195), .C2(n1035), .A(n1036), 
        .ZN(n1029) );
  OAI221_X1 U514 ( .B1(n2210), .B2(n1031), .C1(n2207), .C2(n1032), .A(n1033), 
        .ZN(n1030) );
  NOR4_X1 U515 ( .A1(n1065), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1064) );
  OAI221_X1 U516 ( .B1(n2186), .B2(n1075), .C1(n2183), .C2(n1076), .A(n1077), 
        .ZN(n1066) );
  OAI221_X1 U517 ( .B1(n2198), .B2(n1072), .C1(n2195), .C2(n1073), .A(n1074), 
        .ZN(n1067) );
  OAI221_X1 U518 ( .B1(n2210), .B2(n1069), .C1(n2207), .C2(n1070), .A(n1071), 
        .ZN(n1068) );
  NOR4_X1 U519 ( .A1(n1103), .A2(n1104), .A3(n1105), .A4(n1106), .ZN(n1102) );
  OAI221_X1 U520 ( .B1(n2186), .B2(n1113), .C1(n2183), .C2(n1114), .A(n1115), 
        .ZN(n1104) );
  OAI221_X1 U521 ( .B1(n2198), .B2(n1110), .C1(n2195), .C2(n1111), .A(n1112), 
        .ZN(n1105) );
  OAI221_X1 U522 ( .B1(n2210), .B2(n1107), .C1(n2207), .C2(n1108), .A(n1109), 
        .ZN(n1106) );
  NOR4_X1 U523 ( .A1(n1141), .A2(n1142), .A3(n1143), .A4(n1144), .ZN(n1140) );
  OAI221_X1 U524 ( .B1(n2186), .B2(n1151), .C1(n2183), .C2(n1152), .A(n1153), 
        .ZN(n1142) );
  OAI221_X1 U525 ( .B1(n2198), .B2(n1148), .C1(n2195), .C2(n1149), .A(n1150), 
        .ZN(n1143) );
  OAI221_X1 U526 ( .B1(n2210), .B2(n1145), .C1(n2207), .C2(n1146), .A(n1147), 
        .ZN(n1144) );
  NOR4_X1 U527 ( .A1(n1179), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1178) );
  OAI221_X1 U528 ( .B1(n2186), .B2(n1189), .C1(n2183), .C2(n1190), .A(n1191), 
        .ZN(n1180) );
  OAI221_X1 U529 ( .B1(n2198), .B2(n1186), .C1(n2195), .C2(n1187), .A(n1188), 
        .ZN(n1181) );
  OAI221_X1 U530 ( .B1(n2210), .B2(n1183), .C1(n2207), .C2(n1184), .A(n1185), 
        .ZN(n1182) );
  NOR4_X1 U531 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1216) );
  OAI221_X1 U532 ( .B1(n2186), .B2(n1236), .C1(n2183), .C2(n1237), .A(n1238), 
        .ZN(n1218) );
  OAI221_X1 U533 ( .B1(n2198), .B2(n1231), .C1(n2195), .C2(n1232), .A(n1233), 
        .ZN(n1219) );
  OAI221_X1 U534 ( .B1(n2210), .B2(n1221), .C1(n2207), .C2(n1222), .A(n1223), 
        .ZN(n1220) );
  NOR4_X1 U535 ( .A1(n1776), .A2(n1777), .A3(n1778), .A4(n1779), .ZN(n1775) );
  OAI221_X1 U536 ( .B1(n1037), .B2(n2087), .C1(n1038), .C2(n2084), .A(n1782), 
        .ZN(n1777) );
  OAI221_X1 U537 ( .B1(n1034), .B2(n2099), .C1(n1035), .C2(n2096), .A(n1781), 
        .ZN(n1778) );
  OAI221_X1 U538 ( .B1(n1031), .B2(n2111), .C1(n1032), .C2(n2108), .A(n1780), 
        .ZN(n1779) );
  NOR4_X1 U539 ( .A1(n1794), .A2(n1795), .A3(n1796), .A4(n1797), .ZN(n1793) );
  OAI221_X1 U540 ( .B1(n1075), .B2(n2087), .C1(n1076), .C2(n2084), .A(n1800), 
        .ZN(n1795) );
  OAI221_X1 U541 ( .B1(n1072), .B2(n2099), .C1(n1073), .C2(n2096), .A(n1799), 
        .ZN(n1796) );
  OAI221_X1 U542 ( .B1(n1069), .B2(n2111), .C1(n1070), .C2(n2108), .A(n1798), 
        .ZN(n1797) );
  NOR4_X1 U543 ( .A1(n1812), .A2(n1813), .A3(n1814), .A4(n1815), .ZN(n1811) );
  OAI221_X1 U544 ( .B1(n1113), .B2(n2087), .C1(n1114), .C2(n2084), .A(n1818), 
        .ZN(n1813) );
  OAI221_X1 U545 ( .B1(n1110), .B2(n2099), .C1(n1111), .C2(n2096), .A(n1817), 
        .ZN(n1814) );
  OAI221_X1 U546 ( .B1(n1107), .B2(n2111), .C1(n1108), .C2(n2108), .A(n1816), 
        .ZN(n1815) );
  NOR4_X1 U547 ( .A1(n1830), .A2(n1831), .A3(n1832), .A4(n1833), .ZN(n1829) );
  OAI221_X1 U548 ( .B1(n1151), .B2(n2087), .C1(n1152), .C2(n2084), .A(n1836), 
        .ZN(n1831) );
  OAI221_X1 U549 ( .B1(n1148), .B2(n2099), .C1(n1149), .C2(n2096), .A(n1835), 
        .ZN(n1832) );
  OAI221_X1 U550 ( .B1(n1145), .B2(n2111), .C1(n1146), .C2(n2108), .A(n1834), 
        .ZN(n1833) );
  NOR4_X1 U551 ( .A1(n1848), .A2(n1849), .A3(n1850), .A4(n1851), .ZN(n1847) );
  OAI221_X1 U552 ( .B1(n1189), .B2(n2087), .C1(n1190), .C2(n2084), .A(n1854), 
        .ZN(n1849) );
  OAI221_X1 U553 ( .B1(n1186), .B2(n2099), .C1(n1187), .C2(n2096), .A(n1853), 
        .ZN(n1850) );
  OAI221_X1 U554 ( .B1(n1183), .B2(n2111), .C1(n1184), .C2(n2108), .A(n1852), 
        .ZN(n1851) );
  NOR4_X1 U555 ( .A1(n1866), .A2(n1867), .A3(n1868), .A4(n1869), .ZN(n1865) );
  OAI221_X1 U556 ( .B1(n1236), .B2(n2087), .C1(n1237), .C2(n2084), .A(n1881), 
        .ZN(n1867) );
  OAI221_X1 U557 ( .B1(n1231), .B2(n2099), .C1(n1232), .C2(n2096), .A(n1878), 
        .ZN(n1868) );
  OAI221_X1 U558 ( .B1(n1221), .B2(n2111), .C1(n1222), .C2(n2108), .A(n1870), 
        .ZN(n1869) );
  OAI221_X1 U559 ( .B1(n2184), .B2(n25), .C1(n2181), .C2(n27), .A(n28), .ZN(n7) );
  OAI221_X1 U560 ( .B1(n2196), .B2(n18), .C1(n2193), .C2(n20), .A(n21), .ZN(n8) );
  OAI221_X1 U561 ( .B1(n2208), .B2(n11), .C1(n2205), .C2(n13), .A(n14), .ZN(n9) );
  NOR2_X1 U562 ( .A1(n1269), .A2(n1256), .ZN(n1247) );
  NOR2_X1 U563 ( .A1(n1898), .A2(n1893), .ZN(n1888) );
  OAI22_X1 U564 ( .A1(n1047), .A2(n2062), .B1(n1048), .B2(n2059), .ZN(n1787)
         );
  OAI22_X1 U565 ( .A1(n1085), .A2(n2062), .B1(n1086), .B2(n2059), .ZN(n1805)
         );
  OAI22_X1 U566 ( .A1(n1123), .A2(n2062), .B1(n1124), .B2(n2059), .ZN(n1823)
         );
  OAI22_X1 U567 ( .A1(n1161), .A2(n2062), .B1(n1162), .B2(n2059), .ZN(n1841)
         );
  OAI22_X1 U568 ( .A1(n1199), .A2(n2062), .B1(n1200), .B2(n2059), .ZN(n1859)
         );
  OAI22_X1 U569 ( .A1(n1252), .A2(n2062), .B1(n1253), .B2(n2059), .ZN(n1892)
         );
  OAI22_X1 U570 ( .A1(n2161), .A2(n1047), .B1(n2158), .B2(n1048), .ZN(n1046)
         );
  OAI22_X1 U571 ( .A1(n2161), .A2(n1085), .B1(n2158), .B2(n1086), .ZN(n1084)
         );
  OAI22_X1 U572 ( .A1(n2161), .A2(n1123), .B1(n2158), .B2(n1124), .ZN(n1122)
         );
  OAI22_X1 U573 ( .A1(n2161), .A2(n1161), .B1(n2158), .B2(n1162), .ZN(n1160)
         );
  OAI22_X1 U574 ( .A1(n2161), .A2(n1199), .B1(n2158), .B2(n1200), .ZN(n1198)
         );
  OAI22_X1 U575 ( .A1(n2161), .A2(n1252), .B1(n2158), .B2(n1253), .ZN(n1251)
         );
  OAI22_X1 U576 ( .A1(n2159), .A2(n44), .B1(n2156), .B2(n46), .ZN(n42) );
  OAI22_X1 U577 ( .A1(n2159), .A2(n97), .B1(n2156), .B2(n98), .ZN(n96) );
  OAI22_X1 U578 ( .A1(n2159), .A2(n135), .B1(n2156), .B2(n136), .ZN(n134) );
  OAI22_X1 U579 ( .A1(n2159), .A2(n173), .B1(n2156), .B2(n174), .ZN(n172) );
  OAI22_X1 U580 ( .A1(n2159), .A2(n211), .B1(n2156), .B2(n212), .ZN(n210) );
  OAI22_X1 U581 ( .A1(n2159), .A2(n249), .B1(n2156), .B2(n250), .ZN(n248) );
  OAI22_X1 U582 ( .A1(n2159), .A2(n287), .B1(n2156), .B2(n288), .ZN(n286) );
  OAI22_X1 U583 ( .A1(n2159), .A2(n325), .B1(n2156), .B2(n326), .ZN(n324) );
  OAI22_X1 U584 ( .A1(n2159), .A2(n363), .B1(n2156), .B2(n364), .ZN(n362) );
  OAI22_X1 U585 ( .A1(n2159), .A2(n401), .B1(n2156), .B2(n402), .ZN(n400) );
  OAI22_X1 U586 ( .A1(n2159), .A2(n439), .B1(n2156), .B2(n440), .ZN(n438) );
  OAI22_X1 U587 ( .A1(n2159), .A2(n477), .B1(n2156), .B2(n478), .ZN(n476) );
  OAI22_X1 U588 ( .A1(n2159), .A2(n515), .B1(n2156), .B2(n516), .ZN(n514) );
  OAI22_X1 U589 ( .A1(n2160), .A2(n553), .B1(n2157), .B2(n554), .ZN(n552) );
  OAI22_X1 U590 ( .A1(n2160), .A2(n591), .B1(n2157), .B2(n592), .ZN(n590) );
  OAI22_X1 U591 ( .A1(n2160), .A2(n629), .B1(n2157), .B2(n630), .ZN(n628) );
  OAI22_X1 U592 ( .A1(n2160), .A2(n667), .B1(n2157), .B2(n668), .ZN(n666) );
  OAI22_X1 U593 ( .A1(n2160), .A2(n705), .B1(n2157), .B2(n706), .ZN(n704) );
  OAI22_X1 U594 ( .A1(n2160), .A2(n743), .B1(n2157), .B2(n744), .ZN(n742) );
  OAI22_X1 U595 ( .A1(n2160), .A2(n781), .B1(n2157), .B2(n782), .ZN(n780) );
  OAI22_X1 U596 ( .A1(n2160), .A2(n819), .B1(n2157), .B2(n820), .ZN(n818) );
  OAI22_X1 U597 ( .A1(n2160), .A2(n857), .B1(n2157), .B2(n858), .ZN(n856) );
  OAI22_X1 U600 ( .A1(n2160), .A2(n895), .B1(n2157), .B2(n896), .ZN(n894) );
  OAI22_X1 U601 ( .A1(n2160), .A2(n933), .B1(n2157), .B2(n934), .ZN(n932) );
  OAI22_X1 U602 ( .A1(n2160), .A2(n971), .B1(n2157), .B2(n972), .ZN(n970) );
  OAI22_X1 U603 ( .A1(n2160), .A2(n1009), .B1(n2157), .B2(n1010), .ZN(n1008)
         );
  OAI22_X1 U606 ( .A1(n44), .A2(n2060), .B1(n46), .B2(n2057), .ZN(n1303) );
  OAI22_X1 U607 ( .A1(n97), .A2(n2060), .B1(n98), .B2(n2057), .ZN(n1337) );
  OAI22_X1 U608 ( .A1(n135), .A2(n2060), .B1(n136), .B2(n2057), .ZN(n1355) );
  OAI22_X1 U609 ( .A1(n173), .A2(n2060), .B1(n174), .B2(n2057), .ZN(n1373) );
  OAI22_X1 U612 ( .A1(n211), .A2(n2060), .B1(n212), .B2(n2057), .ZN(n1391) );
  OAI22_X1 U613 ( .A1(n249), .A2(n2060), .B1(n250), .B2(n2057), .ZN(n1409) );
  OAI22_X1 U614 ( .A1(n287), .A2(n2060), .B1(n288), .B2(n2057), .ZN(n1427) );
  OAI22_X1 U615 ( .A1(n325), .A2(n2060), .B1(n326), .B2(n2057), .ZN(n1445) );
  OAI22_X1 U616 ( .A1(n363), .A2(n2060), .B1(n364), .B2(n2057), .ZN(n1463) );
  OAI22_X1 U617 ( .A1(n401), .A2(n2060), .B1(n402), .B2(n2057), .ZN(n1481) );
  OAI22_X1 U619 ( .A1(n439), .A2(n2060), .B1(n440), .B2(n2057), .ZN(n1499) );
  OAI22_X1 U621 ( .A1(n477), .A2(n2060), .B1(n478), .B2(n2057), .ZN(n1517) );
  OAI22_X1 U622 ( .A1(n515), .A2(n2060), .B1(n516), .B2(n2057), .ZN(n1535) );
  OAI22_X1 U623 ( .A1(n553), .A2(n2061), .B1(n554), .B2(n2058), .ZN(n1553) );
  OAI22_X1 U626 ( .A1(n591), .A2(n2061), .B1(n592), .B2(n2058), .ZN(n1571) );
  OAI22_X1 U628 ( .A1(n629), .A2(n2061), .B1(n630), .B2(n2058), .ZN(n1589) );
  OAI22_X1 U630 ( .A1(n667), .A2(n2061), .B1(n668), .B2(n2058), .ZN(n1607) );
  OAI22_X1 U631 ( .A1(n705), .A2(n2061), .B1(n706), .B2(n2058), .ZN(n1625) );
  OAI22_X1 U634 ( .A1(n743), .A2(n2061), .B1(n744), .B2(n2058), .ZN(n1643) );
  OAI22_X1 U635 ( .A1(n781), .A2(n2061), .B1(n782), .B2(n2058), .ZN(n1661) );
  OAI22_X1 U637 ( .A1(n819), .A2(n2061), .B1(n820), .B2(n2058), .ZN(n1679) );
  OAI22_X1 U639 ( .A1(n857), .A2(n2061), .B1(n858), .B2(n2058), .ZN(n1697) );
  OAI22_X1 U640 ( .A1(n895), .A2(n2061), .B1(n896), .B2(n2058), .ZN(n1715) );
  OAI22_X1 U641 ( .A1(n933), .A2(n2061), .B1(n934), .B2(n2058), .ZN(n1733) );
  OAI22_X1 U644 ( .A1(n971), .A2(n2061), .B1(n972), .B2(n2058), .ZN(n1751) );
  OAI22_X1 U645 ( .A1(n1009), .A2(n2061), .B1(n1010), .B2(n2058), .ZN(n1769)
         );
  OAI22_X1 U646 ( .A1(n1049), .A2(n2056), .B1(n1050), .B2(n2053), .ZN(n1786)
         );
  OAI22_X1 U647 ( .A1(n1087), .A2(n2056), .B1(n1088), .B2(n2053), .ZN(n1804)
         );
  OAI22_X1 U648 ( .A1(n1125), .A2(n2056), .B1(n1126), .B2(n2053), .ZN(n1822)
         );
  OAI22_X1 U649 ( .A1(n1163), .A2(n2056), .B1(n1164), .B2(n2053), .ZN(n1840)
         );
  OAI22_X1 U651 ( .A1(n1201), .A2(n2056), .B1(n1202), .B2(n2053), .ZN(n1858)
         );
  OAI22_X1 U653 ( .A1(n1254), .A2(n2056), .B1(n1255), .B2(n2053), .ZN(n1891)
         );
  OAI22_X1 U654 ( .A1(n2155), .A2(n1049), .B1(n2152), .B2(n1050), .ZN(n1045)
         );
  OAI22_X1 U655 ( .A1(n2155), .A2(n1087), .B1(n2152), .B2(n1088), .ZN(n1083)
         );
  OAI22_X1 U656 ( .A1(n2155), .A2(n1125), .B1(n2152), .B2(n1126), .ZN(n1121)
         );
  OAI22_X1 U657 ( .A1(n2155), .A2(n1163), .B1(n2152), .B2(n1164), .ZN(n1159)
         );
  OAI22_X1 U658 ( .A1(n2155), .A2(n1201), .B1(n2152), .B2(n1202), .ZN(n1197)
         );
  OAI22_X1 U659 ( .A1(n2155), .A2(n1254), .B1(n2152), .B2(n1255), .ZN(n1250)
         );
  OAI22_X1 U660 ( .A1(n1056), .A2(n1968), .B1(n1057), .B2(n1965), .ZN(n1788)
         );
  OAI22_X1 U661 ( .A1(n1059), .A2(n1954), .B1(n1060), .B2(n1951), .ZN(n1789)
         );
  OAI22_X1 U662 ( .A1(n1094), .A2(n1968), .B1(n1095), .B2(n1965), .ZN(n1806)
         );
  OAI22_X1 U663 ( .A1(n1097), .A2(n1954), .B1(n1098), .B2(n1951), .ZN(n1807)
         );
  OAI22_X1 U664 ( .A1(n1132), .A2(n1968), .B1(n1133), .B2(n1965), .ZN(n1824)
         );
  OAI22_X1 U665 ( .A1(n1135), .A2(n1954), .B1(n1136), .B2(n1951), .ZN(n1825)
         );
  OAI22_X1 U666 ( .A1(n1170), .A2(n1968), .B1(n1171), .B2(n1965), .ZN(n1842)
         );
  OAI22_X1 U667 ( .A1(n1173), .A2(n1954), .B1(n1174), .B2(n1951), .ZN(n1843)
         );
  OAI22_X1 U668 ( .A1(n1208), .A2(n1968), .B1(n1209), .B2(n1965), .ZN(n1860)
         );
  OAI22_X1 U669 ( .A1(n1211), .A2(n1954), .B1(n1212), .B2(n1951), .ZN(n1861)
         );
  OAI22_X1 U670 ( .A1(n1264), .A2(n1968), .B1(n1265), .B2(n1965), .ZN(n1896)
         );
  OAI22_X1 U671 ( .A1(n1267), .A2(n1954), .B1(n1268), .B2(n1951), .ZN(n1897)
         );
  OAI22_X1 U672 ( .A1(n2131), .A2(n1056), .B1(n2128), .B2(n1057), .ZN(n1055)
         );
  OAI22_X1 U673 ( .A1(n2117), .A2(n1059), .B1(n2114), .B2(n1060), .ZN(n1058)
         );
  OAI22_X1 U674 ( .A1(n2131), .A2(n1094), .B1(n2128), .B2(n1095), .ZN(n1093)
         );
  OAI22_X1 U675 ( .A1(n2117), .A2(n1097), .B1(n2114), .B2(n1098), .ZN(n1096)
         );
  OAI22_X1 U676 ( .A1(n2131), .A2(n1132), .B1(n2128), .B2(n1133), .ZN(n1131)
         );
  OAI22_X1 U677 ( .A1(n2117), .A2(n1135), .B1(n2114), .B2(n1136), .ZN(n1134)
         );
  OAI22_X1 U678 ( .A1(n2131), .A2(n1170), .B1(n2128), .B2(n1171), .ZN(n1169)
         );
  OAI22_X1 U679 ( .A1(n2117), .A2(n1173), .B1(n2114), .B2(n1174), .ZN(n1172)
         );
  OAI22_X1 U680 ( .A1(n2131), .A2(n1208), .B1(n2128), .B2(n1209), .ZN(n1207)
         );
  OAI22_X1 U681 ( .A1(n2117), .A2(n1211), .B1(n2114), .B2(n1212), .ZN(n1210)
         );
  OAI22_X1 U682 ( .A1(n2131), .A2(n1264), .B1(n2128), .B2(n1265), .ZN(n1263)
         );
  OAI22_X1 U683 ( .A1(n2117), .A2(n1267), .B1(n2114), .B2(n1268), .ZN(n1266)
         );
  OAI22_X1 U684 ( .A1(n2153), .A2(n48), .B1(n2150), .B2(n50), .ZN(n41) );
  OAI22_X1 U685 ( .A1(n2153), .A2(n99), .B1(n2150), .B2(n100), .ZN(n95) );
  OAI22_X1 U686 ( .A1(n2153), .A2(n137), .B1(n2150), .B2(n138), .ZN(n133) );
  OAI22_X1 U687 ( .A1(n2153), .A2(n175), .B1(n2150), .B2(n176), .ZN(n171) );
  OAI22_X1 U688 ( .A1(n2153), .A2(n213), .B1(n2150), .B2(n214), .ZN(n209) );
  OAI22_X1 U689 ( .A1(n2153), .A2(n251), .B1(n2150), .B2(n252), .ZN(n247) );
  OAI22_X1 U690 ( .A1(n2153), .A2(n289), .B1(n2150), .B2(n290), .ZN(n285) );
  OAI22_X1 U691 ( .A1(n2153), .A2(n327), .B1(n2150), .B2(n328), .ZN(n323) );
  OAI22_X1 U692 ( .A1(n2153), .A2(n365), .B1(n2150), .B2(n366), .ZN(n361) );
  OAI22_X1 U693 ( .A1(n2153), .A2(n403), .B1(n2150), .B2(n404), .ZN(n399) );
  OAI22_X1 U694 ( .A1(n2153), .A2(n441), .B1(n2150), .B2(n442), .ZN(n437) );
  OAI22_X1 U695 ( .A1(n2153), .A2(n479), .B1(n2150), .B2(n480), .ZN(n475) );
  OAI22_X1 U696 ( .A1(n2153), .A2(n517), .B1(n2150), .B2(n518), .ZN(n513) );
  OAI22_X1 U697 ( .A1(n2154), .A2(n555), .B1(n2151), .B2(n556), .ZN(n551) );
  OAI22_X1 U698 ( .A1(n2154), .A2(n593), .B1(n2151), .B2(n594), .ZN(n589) );
  OAI22_X1 U699 ( .A1(n2154), .A2(n631), .B1(n2151), .B2(n632), .ZN(n627) );
  OAI22_X1 U700 ( .A1(n2154), .A2(n669), .B1(n2151), .B2(n670), .ZN(n665) );
  OAI22_X1 U701 ( .A1(n2154), .A2(n707), .B1(n2151), .B2(n708), .ZN(n703) );
  OAI22_X1 U702 ( .A1(n2154), .A2(n745), .B1(n2151), .B2(n746), .ZN(n741) );
  OAI22_X1 U703 ( .A1(n2154), .A2(n783), .B1(n2151), .B2(n784), .ZN(n779) );
  OAI22_X1 U704 ( .A1(n2154), .A2(n821), .B1(n2151), .B2(n822), .ZN(n817) );
  OAI22_X1 U705 ( .A1(n2154), .A2(n859), .B1(n2151), .B2(n860), .ZN(n855) );
  OAI22_X1 U706 ( .A1(n2154), .A2(n897), .B1(n2151), .B2(n898), .ZN(n893) );
  OAI22_X1 U707 ( .A1(n2154), .A2(n935), .B1(n2151), .B2(n936), .ZN(n931) );
  OAI22_X1 U708 ( .A1(n2154), .A2(n973), .B1(n2151), .B2(n974), .ZN(n969) );
  OAI22_X1 U709 ( .A1(n2154), .A2(n1011), .B1(n2151), .B2(n1012), .ZN(n1007)
         );
  OAI22_X1 U710 ( .A1(n48), .A2(n2054), .B1(n50), .B2(n2051), .ZN(n1302) );
  OAI22_X1 U711 ( .A1(n99), .A2(n2054), .B1(n100), .B2(n2051), .ZN(n1336) );
  OAI22_X1 U712 ( .A1(n137), .A2(n2054), .B1(n138), .B2(n2051), .ZN(n1354) );
  OAI22_X1 U713 ( .A1(n175), .A2(n2054), .B1(n176), .B2(n2051), .ZN(n1372) );
  OAI22_X1 U714 ( .A1(n213), .A2(n2054), .B1(n214), .B2(n2051), .ZN(n1390) );
  OAI22_X1 U715 ( .A1(n251), .A2(n2054), .B1(n252), .B2(n2051), .ZN(n1408) );
  OAI22_X1 U716 ( .A1(n289), .A2(n2054), .B1(n290), .B2(n2051), .ZN(n1426) );
  OAI22_X1 U717 ( .A1(n327), .A2(n2054), .B1(n328), .B2(n2051), .ZN(n1444) );
  OAI22_X1 U718 ( .A1(n365), .A2(n2054), .B1(n366), .B2(n2051), .ZN(n1462) );
  OAI22_X1 U719 ( .A1(n403), .A2(n2054), .B1(n404), .B2(n2051), .ZN(n1480) );
  OAI22_X1 U720 ( .A1(n441), .A2(n2054), .B1(n442), .B2(n2051), .ZN(n1498) );
  OAI22_X1 U721 ( .A1(n479), .A2(n2054), .B1(n480), .B2(n2051), .ZN(n1516) );
  OAI22_X1 U722 ( .A1(n517), .A2(n2054), .B1(n518), .B2(n2051), .ZN(n1534) );
  OAI22_X1 U723 ( .A1(n555), .A2(n2055), .B1(n556), .B2(n2052), .ZN(n1552) );
  OAI22_X1 U724 ( .A1(n593), .A2(n2055), .B1(n594), .B2(n2052), .ZN(n1570) );
  OAI22_X1 U725 ( .A1(n631), .A2(n2055), .B1(n632), .B2(n2052), .ZN(n1588) );
  OAI22_X1 U726 ( .A1(n669), .A2(n2055), .B1(n670), .B2(n2052), .ZN(n1606) );
  OAI22_X1 U727 ( .A1(n707), .A2(n2055), .B1(n708), .B2(n2052), .ZN(n1624) );
  OAI22_X1 U728 ( .A1(n745), .A2(n2055), .B1(n746), .B2(n2052), .ZN(n1642) );
  OAI22_X1 U729 ( .A1(n783), .A2(n2055), .B1(n784), .B2(n2052), .ZN(n1660) );
  OAI22_X1 U730 ( .A1(n821), .A2(n2055), .B1(n822), .B2(n2052), .ZN(n1678) );
  OAI22_X1 U731 ( .A1(n859), .A2(n2055), .B1(n860), .B2(n2052), .ZN(n1696) );
  OAI22_X1 U732 ( .A1(n897), .A2(n2055), .B1(n898), .B2(n2052), .ZN(n1714) );
  OAI22_X1 U733 ( .A1(n935), .A2(n2055), .B1(n936), .B2(n2052), .ZN(n1732) );
  OAI22_X1 U734 ( .A1(n973), .A2(n2055), .B1(n974), .B2(n2052), .ZN(n1750) );
  OAI22_X1 U735 ( .A1(n1011), .A2(n2055), .B1(n1012), .B2(n2052), .ZN(n1768)
         );
  OAI22_X1 U736 ( .A1(n2129), .A2(n63), .B1(n2126), .B2(n65), .ZN(n61) );
  OAI22_X1 U737 ( .A1(n2115), .A2(n70), .B1(n2112), .B2(n72), .ZN(n68) );
  OAI22_X1 U738 ( .A1(n2129), .A2(n106), .B1(n2126), .B2(n107), .ZN(n105) );
  OAI22_X1 U739 ( .A1(n2115), .A2(n109), .B1(n2112), .B2(n110), .ZN(n108) );
  OAI22_X1 U740 ( .A1(n2129), .A2(n144), .B1(n2126), .B2(n145), .ZN(n143) );
  OAI22_X1 U741 ( .A1(n2115), .A2(n147), .B1(n2112), .B2(n148), .ZN(n146) );
  OAI22_X1 U742 ( .A1(n2129), .A2(n182), .B1(n2126), .B2(n183), .ZN(n181) );
  OAI22_X1 U743 ( .A1(n2115), .A2(n185), .B1(n2112), .B2(n186), .ZN(n184) );
  OAI22_X1 U744 ( .A1(n2129), .A2(n220), .B1(n2126), .B2(n221), .ZN(n219) );
  OAI22_X1 U745 ( .A1(n2115), .A2(n223), .B1(n2112), .B2(n224), .ZN(n222) );
  OAI22_X1 U746 ( .A1(n2129), .A2(n258), .B1(n2126), .B2(n259), .ZN(n257) );
  OAI22_X1 U747 ( .A1(n2115), .A2(n261), .B1(n2112), .B2(n262), .ZN(n260) );
  OAI22_X1 U748 ( .A1(n2129), .A2(n296), .B1(n2126), .B2(n297), .ZN(n295) );
  OAI22_X1 U749 ( .A1(n2115), .A2(n299), .B1(n2112), .B2(n300), .ZN(n298) );
  OAI22_X1 U750 ( .A1(n2129), .A2(n334), .B1(n2126), .B2(n335), .ZN(n333) );
  OAI22_X1 U751 ( .A1(n2115), .A2(n337), .B1(n2112), .B2(n338), .ZN(n336) );
  OAI22_X1 U752 ( .A1(n2129), .A2(n372), .B1(n2126), .B2(n373), .ZN(n371) );
  OAI22_X1 U753 ( .A1(n2115), .A2(n375), .B1(n2112), .B2(n376), .ZN(n374) );
  OAI22_X1 U754 ( .A1(n2129), .A2(n410), .B1(n2126), .B2(n411), .ZN(n409) );
  OAI22_X1 U755 ( .A1(n2115), .A2(n413), .B1(n2112), .B2(n414), .ZN(n412) );
  OAI22_X1 U756 ( .A1(n2129), .A2(n448), .B1(n2126), .B2(n449), .ZN(n447) );
  OAI22_X1 U757 ( .A1(n2115), .A2(n451), .B1(n2112), .B2(n452), .ZN(n450) );
  OAI22_X1 U758 ( .A1(n2129), .A2(n486), .B1(n2126), .B2(n487), .ZN(n485) );
  OAI22_X1 U759 ( .A1(n2115), .A2(n489), .B1(n2112), .B2(n490), .ZN(n488) );
  OAI22_X1 U760 ( .A1(n2129), .A2(n524), .B1(n2126), .B2(n525), .ZN(n523) );
  OAI22_X1 U761 ( .A1(n2115), .A2(n527), .B1(n2112), .B2(n528), .ZN(n526) );
  OAI22_X1 U762 ( .A1(n2130), .A2(n562), .B1(n2127), .B2(n563), .ZN(n561) );
  OAI22_X1 U763 ( .A1(n2116), .A2(n565), .B1(n2113), .B2(n566), .ZN(n564) );
  OAI22_X1 U764 ( .A1(n2130), .A2(n600), .B1(n2127), .B2(n601), .ZN(n599) );
  OAI22_X1 U765 ( .A1(n2116), .A2(n603), .B1(n2113), .B2(n604), .ZN(n602) );
  OAI22_X1 U766 ( .A1(n2130), .A2(n638), .B1(n2127), .B2(n639), .ZN(n637) );
  OAI22_X1 U767 ( .A1(n2116), .A2(n641), .B1(n2113), .B2(n642), .ZN(n640) );
  OAI22_X1 U768 ( .A1(n2130), .A2(n676), .B1(n2127), .B2(n677), .ZN(n675) );
  OAI22_X1 U769 ( .A1(n2116), .A2(n679), .B1(n2113), .B2(n680), .ZN(n678) );
  OAI22_X1 U770 ( .A1(n2130), .A2(n714), .B1(n2127), .B2(n715), .ZN(n713) );
  OAI22_X1 U771 ( .A1(n2116), .A2(n717), .B1(n2113), .B2(n718), .ZN(n716) );
  OAI22_X1 U772 ( .A1(n2130), .A2(n752), .B1(n2127), .B2(n753), .ZN(n751) );
  OAI22_X1 U773 ( .A1(n2116), .A2(n755), .B1(n2113), .B2(n756), .ZN(n754) );
  OAI22_X1 U774 ( .A1(n2130), .A2(n790), .B1(n2127), .B2(n791), .ZN(n789) );
  OAI22_X1 U775 ( .A1(n2116), .A2(n793), .B1(n2113), .B2(n794), .ZN(n792) );
  OAI22_X1 U776 ( .A1(n2130), .A2(n828), .B1(n2127), .B2(n829), .ZN(n827) );
  OAI22_X1 U777 ( .A1(n2116), .A2(n831), .B1(n2113), .B2(n832), .ZN(n830) );
  OAI22_X1 U778 ( .A1(n2130), .A2(n866), .B1(n2127), .B2(n867), .ZN(n865) );
  OAI22_X1 U779 ( .A1(n2116), .A2(n869), .B1(n2113), .B2(n870), .ZN(n868) );
  OAI22_X1 U780 ( .A1(n2130), .A2(n904), .B1(n2127), .B2(n905), .ZN(n903) );
  OAI22_X1 U781 ( .A1(n2116), .A2(n907), .B1(n2113), .B2(n908), .ZN(n906) );
  OAI22_X1 U782 ( .A1(n2130), .A2(n942), .B1(n2127), .B2(n943), .ZN(n941) );
  OAI22_X1 U783 ( .A1(n2116), .A2(n945), .B1(n2113), .B2(n946), .ZN(n944) );
  OAI22_X1 U784 ( .A1(n2130), .A2(n980), .B1(n2127), .B2(n981), .ZN(n979) );
  OAI22_X1 U785 ( .A1(n2116), .A2(n983), .B1(n2113), .B2(n984), .ZN(n982) );
  OAI22_X1 U786 ( .A1(n2130), .A2(n1018), .B1(n2127), .B2(n1019), .ZN(n1017)
         );
  OAI22_X1 U787 ( .A1(n2116), .A2(n1021), .B1(n2113), .B2(n1022), .ZN(n1020)
         );
  OAI22_X1 U788 ( .A1(n63), .A2(n1966), .B1(n65), .B2(n1963), .ZN(n1314) );
  OAI22_X1 U789 ( .A1(n70), .A2(n1952), .B1(n72), .B2(n1949), .ZN(n1319) );
  OAI22_X1 U790 ( .A1(n106), .A2(n1966), .B1(n107), .B2(n1963), .ZN(n1338) );
  OAI22_X1 U791 ( .A1(n109), .A2(n1952), .B1(n110), .B2(n1949), .ZN(n1339) );
  OAI22_X1 U792 ( .A1(n144), .A2(n1966), .B1(n145), .B2(n1963), .ZN(n1356) );
  OAI22_X1 U793 ( .A1(n147), .A2(n1952), .B1(n148), .B2(n1949), .ZN(n1357) );
  OAI22_X1 U794 ( .A1(n182), .A2(n1966), .B1(n183), .B2(n1963), .ZN(n1374) );
  OAI22_X1 U795 ( .A1(n185), .A2(n1952), .B1(n186), .B2(n1949), .ZN(n1375) );
  OAI22_X1 U796 ( .A1(n220), .A2(n1966), .B1(n221), .B2(n1963), .ZN(n1392) );
  OAI22_X1 U797 ( .A1(n223), .A2(n1952), .B1(n224), .B2(n1949), .ZN(n1393) );
  OAI22_X1 U798 ( .A1(n258), .A2(n1966), .B1(n259), .B2(n1963), .ZN(n1410) );
  OAI22_X1 U799 ( .A1(n261), .A2(n1952), .B1(n262), .B2(n1949), .ZN(n1411) );
  OAI22_X1 U800 ( .A1(n296), .A2(n1966), .B1(n297), .B2(n1963), .ZN(n1428) );
  OAI22_X1 U801 ( .A1(n299), .A2(n1952), .B1(n300), .B2(n1949), .ZN(n1429) );
  OAI22_X1 U802 ( .A1(n334), .A2(n1966), .B1(n335), .B2(n1963), .ZN(n1446) );
  OAI22_X1 U803 ( .A1(n337), .A2(n1952), .B1(n338), .B2(n1949), .ZN(n1447) );
  OAI22_X1 U804 ( .A1(n372), .A2(n1966), .B1(n373), .B2(n1963), .ZN(n1464) );
  OAI22_X1 U805 ( .A1(n375), .A2(n1952), .B1(n376), .B2(n1949), .ZN(n1465) );
  OAI22_X1 U806 ( .A1(n410), .A2(n1966), .B1(n411), .B2(n1963), .ZN(n1482) );
  OAI22_X1 U807 ( .A1(n413), .A2(n1952), .B1(n414), .B2(n1949), .ZN(n1483) );
  OAI22_X1 U808 ( .A1(n448), .A2(n1966), .B1(n449), .B2(n1963), .ZN(n1500) );
  OAI22_X1 U809 ( .A1(n451), .A2(n1952), .B1(n452), .B2(n1949), .ZN(n1501) );
  OAI22_X1 U810 ( .A1(n486), .A2(n1966), .B1(n487), .B2(n1963), .ZN(n1518) );
  OAI22_X1 U811 ( .A1(n489), .A2(n1952), .B1(n490), .B2(n1949), .ZN(n1519) );
  OAI22_X1 U812 ( .A1(n524), .A2(n1966), .B1(n525), .B2(n1963), .ZN(n1536) );
  OAI22_X1 U813 ( .A1(n527), .A2(n1952), .B1(n528), .B2(n1949), .ZN(n1537) );
  OAI22_X1 U814 ( .A1(n562), .A2(n1967), .B1(n563), .B2(n1964), .ZN(n1554) );
  OAI22_X1 U815 ( .A1(n565), .A2(n1953), .B1(n566), .B2(n1950), .ZN(n1555) );
  OAI22_X1 U816 ( .A1(n600), .A2(n1967), .B1(n601), .B2(n1964), .ZN(n1572) );
  OAI22_X1 U817 ( .A1(n603), .A2(n1953), .B1(n604), .B2(n1950), .ZN(n1573) );
  OAI22_X1 U818 ( .A1(n638), .A2(n1967), .B1(n639), .B2(n1964), .ZN(n1590) );
  OAI22_X1 U819 ( .A1(n641), .A2(n1953), .B1(n642), .B2(n1950), .ZN(n1591) );
  OAI22_X1 U820 ( .A1(n676), .A2(n1967), .B1(n677), .B2(n1964), .ZN(n1608) );
  OAI22_X1 U821 ( .A1(n679), .A2(n1953), .B1(n680), .B2(n1950), .ZN(n1609) );
  OAI22_X1 U822 ( .A1(n714), .A2(n1967), .B1(n715), .B2(n1964), .ZN(n1626) );
  OAI22_X1 U823 ( .A1(n717), .A2(n1953), .B1(n718), .B2(n1950), .ZN(n1627) );
  OAI22_X1 U824 ( .A1(n752), .A2(n1967), .B1(n753), .B2(n1964), .ZN(n1644) );
  OAI22_X1 U825 ( .A1(n755), .A2(n1953), .B1(n756), .B2(n1950), .ZN(n1645) );
  OAI22_X1 U826 ( .A1(n790), .A2(n1967), .B1(n791), .B2(n1964), .ZN(n1662) );
  OAI22_X1 U827 ( .A1(n793), .A2(n1953), .B1(n794), .B2(n1950), .ZN(n1663) );
  OAI22_X1 U828 ( .A1(n828), .A2(n1967), .B1(n829), .B2(n1964), .ZN(n1680) );
  OAI22_X1 U829 ( .A1(n831), .A2(n1953), .B1(n832), .B2(n1950), .ZN(n1681) );
  OAI22_X1 U830 ( .A1(n866), .A2(n1967), .B1(n867), .B2(n1964), .ZN(n1698) );
  OAI22_X1 U831 ( .A1(n869), .A2(n1953), .B1(n870), .B2(n1950), .ZN(n1699) );
  OAI22_X1 U832 ( .A1(n904), .A2(n1967), .B1(n905), .B2(n1964), .ZN(n1716) );
  OAI22_X1 U833 ( .A1(n907), .A2(n1953), .B1(n908), .B2(n1950), .ZN(n1717) );
  OAI22_X1 U834 ( .A1(n942), .A2(n1967), .B1(n943), .B2(n1964), .ZN(n1734) );
  OAI22_X1 U835 ( .A1(n945), .A2(n1953), .B1(n946), .B2(n1950), .ZN(n1735) );
  OAI22_X1 U836 ( .A1(n980), .A2(n1967), .B1(n981), .B2(n1964), .ZN(n1752) );
  OAI22_X1 U837 ( .A1(n983), .A2(n1953), .B1(n984), .B2(n1950), .ZN(n1753) );
  OAI22_X1 U838 ( .A1(n1018), .A2(n1967), .B1(n1019), .B2(n1964), .ZN(n1770)
         );
  OAI22_X1 U839 ( .A1(n1021), .A2(n1953), .B1(n1022), .B2(n1950), .ZN(n1771)
         );
  OAI22_X1 U840 ( .A1(n1051), .A2(n2050), .B1(n1052), .B2(n2047), .ZN(n1785)
         );
  OAI22_X1 U841 ( .A1(n1089), .A2(n2050), .B1(n1090), .B2(n2047), .ZN(n1803)
         );
  OAI22_X1 U842 ( .A1(n1127), .A2(n2050), .B1(n1128), .B2(n2047), .ZN(n1821)
         );
  OAI22_X1 U843 ( .A1(n1165), .A2(n2050), .B1(n1166), .B2(n2047), .ZN(n1839)
         );
  OAI22_X1 U844 ( .A1(n1203), .A2(n2050), .B1(n1204), .B2(n2047), .ZN(n1857)
         );
  OAI22_X1 U845 ( .A1(n1257), .A2(n2050), .B1(n1258), .B2(n2047), .ZN(n1890)
         );
  OAI22_X1 U846 ( .A1(n2149), .A2(n1051), .B1(n2146), .B2(n1052), .ZN(n1044)
         );
  OAI22_X1 U847 ( .A1(n2149), .A2(n1089), .B1(n2146), .B2(n1090), .ZN(n1082)
         );
  OAI22_X1 U848 ( .A1(n2149), .A2(n1127), .B1(n2146), .B2(n1128), .ZN(n1120)
         );
  OAI22_X1 U849 ( .A1(n2149), .A2(n1165), .B1(n2146), .B2(n1166), .ZN(n1158)
         );
  OAI22_X1 U850 ( .A1(n2149), .A2(n1203), .B1(n2146), .B2(n1204), .ZN(n1196)
         );
  OAI22_X1 U851 ( .A1(n2149), .A2(n1257), .B1(n2146), .B2(n1258), .ZN(n1249)
         );
  OAI22_X1 U852 ( .A1(n1053), .A2(n2044), .B1(n1054), .B2(n1977), .ZN(n1784)
         );
  OAI22_X1 U853 ( .A1(n1091), .A2(n2044), .B1(n1092), .B2(n1977), .ZN(n1802)
         );
  OAI22_X1 U854 ( .A1(n1129), .A2(n2044), .B1(n1130), .B2(n1977), .ZN(n1820)
         );
  OAI22_X1 U855 ( .A1(n1167), .A2(n2044), .B1(n1168), .B2(n1977), .ZN(n1838)
         );
  OAI22_X1 U856 ( .A1(n1205), .A2(n2044), .B1(n1206), .B2(n1977), .ZN(n1856)
         );
  OAI22_X1 U857 ( .A1(n1260), .A2(n2044), .B1(n1261), .B2(n1977), .ZN(n1889)
         );
  OAI22_X1 U858 ( .A1(n2143), .A2(n1053), .B1(n2140), .B2(n1054), .ZN(n1043)
         );
  OAI22_X1 U859 ( .A1(n2143), .A2(n1091), .B1(n2140), .B2(n1092), .ZN(n1081)
         );
  OAI22_X1 U860 ( .A1(n2143), .A2(n1129), .B1(n2140), .B2(n1130), .ZN(n1119)
         );
  OAI22_X1 U861 ( .A1(n2143), .A2(n1167), .B1(n2140), .B2(n1168), .ZN(n1157)
         );
  OAI22_X1 U862 ( .A1(n2143), .A2(n1205), .B1(n2140), .B2(n1206), .ZN(n1195)
         );
  OAI22_X1 U863 ( .A1(n2143), .A2(n1260), .B1(n2140), .B2(n1261), .ZN(n1248)
         );
  OAI22_X1 U864 ( .A1(n2147), .A2(n52), .B1(n2144), .B2(n54), .ZN(n40) );
  OAI22_X1 U865 ( .A1(n2147), .A2(n101), .B1(n2144), .B2(n102), .ZN(n94) );
  OAI22_X1 U866 ( .A1(n2147), .A2(n139), .B1(n2144), .B2(n140), .ZN(n132) );
  OAI22_X1 U867 ( .A1(n2147), .A2(n177), .B1(n2144), .B2(n178), .ZN(n170) );
  OAI22_X1 U868 ( .A1(n2147), .A2(n215), .B1(n2144), .B2(n216), .ZN(n208) );
  OAI22_X1 U869 ( .A1(n2147), .A2(n253), .B1(n2144), .B2(n254), .ZN(n246) );
  OAI22_X1 U870 ( .A1(n2147), .A2(n291), .B1(n2144), .B2(n292), .ZN(n284) );
  OAI22_X1 U871 ( .A1(n2147), .A2(n329), .B1(n2144), .B2(n330), .ZN(n322) );
  OAI22_X1 U872 ( .A1(n2147), .A2(n367), .B1(n2144), .B2(n368), .ZN(n360) );
  OAI22_X1 U873 ( .A1(n2147), .A2(n405), .B1(n2144), .B2(n406), .ZN(n398) );
  OAI22_X1 U874 ( .A1(n2147), .A2(n443), .B1(n2144), .B2(n444), .ZN(n436) );
  OAI22_X1 U875 ( .A1(n2147), .A2(n481), .B1(n2144), .B2(n482), .ZN(n474) );
  OAI22_X1 U876 ( .A1(n2147), .A2(n519), .B1(n2144), .B2(n520), .ZN(n512) );
  OAI22_X1 U877 ( .A1(n2148), .A2(n557), .B1(n2145), .B2(n558), .ZN(n550) );
  OAI22_X1 U878 ( .A1(n2148), .A2(n595), .B1(n2145), .B2(n596), .ZN(n588) );
  OAI22_X1 U879 ( .A1(n2148), .A2(n633), .B1(n2145), .B2(n634), .ZN(n626) );
  OAI22_X1 U880 ( .A1(n2148), .A2(n671), .B1(n2145), .B2(n672), .ZN(n664) );
  OAI22_X1 U881 ( .A1(n2148), .A2(n709), .B1(n2145), .B2(n710), .ZN(n702) );
  OAI22_X1 U882 ( .A1(n2148), .A2(n747), .B1(n2145), .B2(n748), .ZN(n740) );
  OAI22_X1 U883 ( .A1(n2148), .A2(n785), .B1(n2145), .B2(n786), .ZN(n778) );
  OAI22_X1 U884 ( .A1(n2148), .A2(n823), .B1(n2145), .B2(n824), .ZN(n816) );
  OAI22_X1 U885 ( .A1(n2148), .A2(n861), .B1(n2145), .B2(n862), .ZN(n854) );
  OAI22_X1 U886 ( .A1(n2148), .A2(n899), .B1(n2145), .B2(n900), .ZN(n892) );
  OAI22_X1 U887 ( .A1(n2148), .A2(n937), .B1(n2145), .B2(n938), .ZN(n930) );
  OAI22_X1 U888 ( .A1(n2148), .A2(n975), .B1(n2145), .B2(n976), .ZN(n968) );
  OAI22_X1 U889 ( .A1(n2148), .A2(n1013), .B1(n2145), .B2(n1014), .ZN(n1006)
         );
  OAI22_X1 U890 ( .A1(n52), .A2(n2048), .B1(n54), .B2(n2045), .ZN(n1301) );
  OAI22_X1 U891 ( .A1(n101), .A2(n2048), .B1(n102), .B2(n2045), .ZN(n1335) );
  OAI22_X1 U892 ( .A1(n139), .A2(n2048), .B1(n140), .B2(n2045), .ZN(n1353) );
  OAI22_X1 U893 ( .A1(n177), .A2(n2048), .B1(n178), .B2(n2045), .ZN(n1371) );
  OAI22_X1 U894 ( .A1(n215), .A2(n2048), .B1(n216), .B2(n2045), .ZN(n1389) );
  OAI22_X1 U895 ( .A1(n253), .A2(n2048), .B1(n254), .B2(n2045), .ZN(n1407) );
  OAI22_X1 U896 ( .A1(n291), .A2(n2048), .B1(n292), .B2(n2045), .ZN(n1425) );
  OAI22_X1 U897 ( .A1(n329), .A2(n2048), .B1(n330), .B2(n2045), .ZN(n1443) );
  OAI22_X1 U898 ( .A1(n367), .A2(n2048), .B1(n368), .B2(n2045), .ZN(n1461) );
  OAI22_X1 U899 ( .A1(n405), .A2(n2048), .B1(n406), .B2(n2045), .ZN(n1479) );
  OAI22_X1 U900 ( .A1(n443), .A2(n2048), .B1(n444), .B2(n2045), .ZN(n1497) );
  OAI22_X1 U901 ( .A1(n481), .A2(n2048), .B1(n482), .B2(n2045), .ZN(n1515) );
  OAI22_X1 U902 ( .A1(n519), .A2(n2048), .B1(n520), .B2(n2045), .ZN(n1533) );
  OAI22_X1 U903 ( .A1(n557), .A2(n2049), .B1(n558), .B2(n2046), .ZN(n1551) );
  OAI22_X1 U904 ( .A1(n595), .A2(n2049), .B1(n596), .B2(n2046), .ZN(n1569) );
  OAI22_X1 U905 ( .A1(n633), .A2(n2049), .B1(n634), .B2(n2046), .ZN(n1587) );
  OAI22_X1 U906 ( .A1(n671), .A2(n2049), .B1(n672), .B2(n2046), .ZN(n1605) );
  OAI22_X1 U907 ( .A1(n709), .A2(n2049), .B1(n710), .B2(n2046), .ZN(n1623) );
  OAI22_X1 U908 ( .A1(n747), .A2(n2049), .B1(n748), .B2(n2046), .ZN(n1641) );
  OAI22_X1 U909 ( .A1(n785), .A2(n2049), .B1(n786), .B2(n2046), .ZN(n1659) );
  OAI22_X1 U910 ( .A1(n823), .A2(n2049), .B1(n824), .B2(n2046), .ZN(n1677) );
  OAI22_X1 U911 ( .A1(n861), .A2(n2049), .B1(n862), .B2(n2046), .ZN(n1695) );
  OAI22_X1 U912 ( .A1(n899), .A2(n2049), .B1(n900), .B2(n2046), .ZN(n1713) );
  OAI22_X1 U913 ( .A1(n937), .A2(n2049), .B1(n938), .B2(n2046), .ZN(n1731) );
  OAI22_X1 U914 ( .A1(n975), .A2(n2049), .B1(n976), .B2(n2046), .ZN(n1749) );
  OAI22_X1 U915 ( .A1(n1013), .A2(n2049), .B1(n1014), .B2(n2046), .ZN(n1767)
         );
  OAI22_X1 U916 ( .A1(n2141), .A2(n103), .B1(n2138), .B2(n104), .ZN(n93) );
  OAI22_X1 U917 ( .A1(n2141), .A2(n141), .B1(n2138), .B2(n142), .ZN(n131) );
  OAI22_X1 U918 ( .A1(n2141), .A2(n179), .B1(n2138), .B2(n180), .ZN(n169) );
  OAI22_X1 U919 ( .A1(n2141), .A2(n217), .B1(n2138), .B2(n218), .ZN(n207) );
  OAI22_X1 U920 ( .A1(n2141), .A2(n255), .B1(n2138), .B2(n256), .ZN(n245) );
  OAI22_X1 U921 ( .A1(n2141), .A2(n293), .B1(n2138), .B2(n294), .ZN(n283) );
  OAI22_X1 U922 ( .A1(n2141), .A2(n331), .B1(n2138), .B2(n332), .ZN(n321) );
  OAI22_X1 U923 ( .A1(n2141), .A2(n369), .B1(n2138), .B2(n370), .ZN(n359) );
  OAI22_X1 U924 ( .A1(n2141), .A2(n407), .B1(n2138), .B2(n408), .ZN(n397) );
  OAI22_X1 U925 ( .A1(n2141), .A2(n445), .B1(n2138), .B2(n446), .ZN(n435) );
  OAI22_X1 U926 ( .A1(n2141), .A2(n483), .B1(n2138), .B2(n484), .ZN(n473) );
  OAI22_X1 U927 ( .A1(n2141), .A2(n521), .B1(n2138), .B2(n522), .ZN(n511) );
  OAI22_X1 U928 ( .A1(n2142), .A2(n559), .B1(n2139), .B2(n560), .ZN(n549) );
  OAI22_X1 U929 ( .A1(n2142), .A2(n597), .B1(n2139), .B2(n598), .ZN(n587) );
  OAI22_X1 U930 ( .A1(n2142), .A2(n635), .B1(n2139), .B2(n636), .ZN(n625) );
  OAI22_X1 U931 ( .A1(n2142), .A2(n673), .B1(n2139), .B2(n674), .ZN(n663) );
  OAI22_X1 U932 ( .A1(n2142), .A2(n711), .B1(n2139), .B2(n712), .ZN(n701) );
  OAI22_X1 U933 ( .A1(n2142), .A2(n749), .B1(n2139), .B2(n750), .ZN(n739) );
  OAI22_X1 U934 ( .A1(n2142), .A2(n787), .B1(n2139), .B2(n788), .ZN(n777) );
  OAI22_X1 U935 ( .A1(n2142), .A2(n825), .B1(n2139), .B2(n826), .ZN(n815) );
  OAI22_X1 U936 ( .A1(n2142), .A2(n863), .B1(n2139), .B2(n864), .ZN(n853) );
  OAI22_X1 U937 ( .A1(n2142), .A2(n901), .B1(n2139), .B2(n902), .ZN(n891) );
  OAI22_X1 U938 ( .A1(n2142), .A2(n939), .B1(n2139), .B2(n940), .ZN(n929) );
  OAI22_X1 U939 ( .A1(n2142), .A2(n977), .B1(n2139), .B2(n978), .ZN(n967) );
  OAI22_X1 U940 ( .A1(n2142), .A2(n1015), .B1(n2139), .B2(n1016), .ZN(n1005)
         );
  OAI22_X1 U941 ( .A1(n56), .A2(n1978), .B1(n58), .B2(n1975), .ZN(n1300) );
  OAI22_X1 U942 ( .A1(n103), .A2(n1978), .B1(n104), .B2(n1975), .ZN(n1334) );
  OAI22_X1 U943 ( .A1(n141), .A2(n1978), .B1(n142), .B2(n1975), .ZN(n1352) );
  OAI22_X1 U944 ( .A1(n179), .A2(n1978), .B1(n180), .B2(n1975), .ZN(n1370) );
  OAI22_X1 U945 ( .A1(n217), .A2(n1978), .B1(n218), .B2(n1975), .ZN(n1388) );
  OAI22_X1 U946 ( .A1(n255), .A2(n1978), .B1(n256), .B2(n1975), .ZN(n1406) );
  OAI22_X1 U947 ( .A1(n293), .A2(n1978), .B1(n294), .B2(n1975), .ZN(n1424) );
  OAI22_X1 U948 ( .A1(n331), .A2(n1978), .B1(n332), .B2(n1975), .ZN(n1442) );
  OAI22_X1 U949 ( .A1(n369), .A2(n1978), .B1(n370), .B2(n1975), .ZN(n1460) );
  OAI22_X1 U950 ( .A1(n407), .A2(n1978), .B1(n408), .B2(n1975), .ZN(n1478) );
  OAI22_X1 U951 ( .A1(n445), .A2(n1978), .B1(n446), .B2(n1975), .ZN(n1496) );
  OAI22_X1 U952 ( .A1(n483), .A2(n1978), .B1(n484), .B2(n1975), .ZN(n1514) );
  OAI22_X1 U953 ( .A1(n521), .A2(n1978), .B1(n522), .B2(n1975), .ZN(n1532) );
  OAI22_X1 U954 ( .A1(n559), .A2(n1979), .B1(n560), .B2(n1976), .ZN(n1550) );
  OAI22_X1 U955 ( .A1(n597), .A2(n1979), .B1(n598), .B2(n1976), .ZN(n1568) );
  OAI22_X1 U956 ( .A1(n635), .A2(n1979), .B1(n636), .B2(n1976), .ZN(n1586) );
  OAI22_X1 U957 ( .A1(n673), .A2(n1979), .B1(n674), .B2(n1976), .ZN(n1604) );
  OAI22_X1 U958 ( .A1(n711), .A2(n1979), .B1(n712), .B2(n1976), .ZN(n1622) );
  OAI22_X1 U959 ( .A1(n749), .A2(n1979), .B1(n750), .B2(n1976), .ZN(n1640) );
  OAI22_X1 U960 ( .A1(n787), .A2(n1979), .B1(n788), .B2(n1976), .ZN(n1658) );
  OAI22_X1 U961 ( .A1(n825), .A2(n1979), .B1(n826), .B2(n1976), .ZN(n1676) );
  OAI22_X1 U962 ( .A1(n863), .A2(n1979), .B1(n864), .B2(n1976), .ZN(n1694) );
  OAI22_X1 U963 ( .A1(n901), .A2(n1979), .B1(n902), .B2(n1976), .ZN(n1712) );
  OAI22_X1 U964 ( .A1(n939), .A2(n1979), .B1(n940), .B2(n1976), .ZN(n1730) );
  OAI22_X1 U965 ( .A1(n977), .A2(n1979), .B1(n978), .B2(n1976), .ZN(n1748) );
  OAI22_X1 U966 ( .A1(n1015), .A2(n1979), .B1(n1016), .B2(n1976), .ZN(n1766)
         );
  OAI22_X1 U967 ( .A1(n2141), .A2(n56), .B1(n2138), .B2(n58), .ZN(n39) );
  AND2_X1 U968 ( .A1(n1874), .A2(n1875), .ZN(n1299) );
  AND3_X1 U969 ( .A1(n1226), .A2(n2121), .A3(n1230), .ZN(n60) );
  AND3_X1 U970 ( .A1(n1873), .A2(n1958), .A3(n1877), .ZN(n1313) );
  AND3_X1 U971 ( .A1(n1247), .A2(n2121), .A3(n1234), .ZN(n59) );
  AND3_X1 U972 ( .A1(n1247), .A2(n2121), .A3(n1224), .ZN(n66) );
  AND3_X1 U973 ( .A1(n1888), .A2(n1958), .A3(n1879), .ZN(n1312) );
  AND3_X1 U974 ( .A1(n1888), .A2(n1958), .A3(n1871), .ZN(n1317) );
  AND2_X1 U975 ( .A1(n1234), .A2(n1225), .ZN(n23) );
  AND2_X1 U976 ( .A1(n1871), .A2(n1872), .ZN(n1283) );
  AND2_X1 U977 ( .A1(n1879), .A2(n1872), .ZN(n1288) );
  AND2_X1 U978 ( .A1(n1226), .A2(n1227), .ZN(n15) );
  AND2_X1 U979 ( .A1(n1235), .A2(n1227), .ZN(n22) );
  AND2_X1 U980 ( .A1(n1873), .A2(n1874), .ZN(n1282) );
  AND2_X1 U981 ( .A1(n1880), .A2(n1874), .ZN(n1287) );
  AND2_X1 U982 ( .A1(n1241), .A2(n1227), .ZN(n29) );
  AND2_X1 U983 ( .A1(n1884), .A2(n1874), .ZN(n1292) );
  AND2_X1 U984 ( .A1(n1245), .A2(n1225), .ZN(n36) );
  AND2_X1 U985 ( .A1(n1239), .A2(n1240), .ZN(n30) );
  AND2_X1 U986 ( .A1(n1886), .A2(n1872), .ZN(n1297) );
  AND2_X1 U987 ( .A1(n1882), .A2(n1883), .ZN(n1293) );
  INV_X1 U988 ( .A(RST), .ZN(n1916) );
  OAI21_X1 U989 ( .B1(n1899), .B2(n1907), .A(n1876), .ZN(N2930) );
  OAI21_X1 U990 ( .B1(n1899), .B2(n1906), .A(n1270), .ZN(N2994) );
  OAI21_X1 U991 ( .B1(n1899), .B2(n1905), .A(n1270), .ZN(N3058) );
  OAI21_X1 U992 ( .B1(n1899), .B2(n1904), .A(n1270), .ZN(N3122) );
  OAI21_X1 U993 ( .B1(n1899), .B2(n1903), .A(n1270), .ZN(N3186) );
  OAI21_X1 U994 ( .B1(n1899), .B2(n1902), .A(n1270), .ZN(N3250) );
  OAI21_X1 U995 ( .B1(n1899), .B2(n1901), .A(n1270), .ZN(N3314) );
  OAI21_X1 U996 ( .B1(n1899), .B2(n1900), .A(n1876), .ZN(N3378) );
  OAI21_X1 U997 ( .B1(n1906), .B2(n1912), .A(n1876), .ZN(N1458) );
  OAI21_X1 U998 ( .B1(n1905), .B2(n1912), .A(n1876), .ZN(N1522) );
  OAI21_X1 U999 ( .B1(n1904), .B2(n1912), .A(n1876), .ZN(N1586) );
  OAI21_X1 U1000 ( .B1(n1903), .B2(n1912), .A(n1876), .ZN(N1650) );
  OAI21_X1 U1001 ( .B1(n1902), .B2(n1912), .A(n1876), .ZN(N1714) );
  OAI21_X1 U1002 ( .B1(n1901), .B2(n1912), .A(n1876), .ZN(N1778) );
  OAI21_X1 U1003 ( .B1(n1900), .B2(n1912), .A(n1876), .ZN(N1842) );
  OAI21_X1 U1004 ( .B1(n1907), .B2(n1910), .A(n1876), .ZN(N1906) );
  OAI21_X1 U1005 ( .B1(n1906), .B2(n1910), .A(n1876), .ZN(N1970) );
  OAI21_X1 U1006 ( .B1(n1905), .B2(n1910), .A(n1876), .ZN(N2034) );
  OAI21_X1 U1007 ( .B1(n1904), .B2(n1910), .A(n1876), .ZN(N2098) );
  OAI21_X1 U1008 ( .B1(n1903), .B2(n1910), .A(n1270), .ZN(N2162) );
  OAI21_X1 U1009 ( .B1(n1902), .B2(n1910), .A(n1876), .ZN(N2226) );
  OAI21_X1 U1010 ( .B1(n1901), .B2(n1910), .A(n1876), .ZN(N2290) );
  OAI21_X1 U1011 ( .B1(n1900), .B2(n1910), .A(n1876), .ZN(N2354) );
  OAI21_X1 U1012 ( .B1(n1907), .B2(n1908), .A(n1876), .ZN(N2418) );
  OAI21_X1 U1013 ( .B1(n1906), .B2(n1908), .A(n1876), .ZN(N2482) );
  OAI21_X1 U1014 ( .B1(n1905), .B2(n1908), .A(n1876), .ZN(N2546) );
  OAI21_X1 U1015 ( .B1(n1904), .B2(n1908), .A(n1876), .ZN(N2610) );
  OAI21_X1 U1016 ( .B1(n1903), .B2(n1908), .A(n1876), .ZN(N2674) );
  OAI21_X1 U1017 ( .B1(n1902), .B2(n1908), .A(n1876), .ZN(N2738) );
  OAI21_X1 U1018 ( .B1(n1901), .B2(n1908), .A(n1876), .ZN(N2802) );
  OAI21_X1 U1019 ( .B1(n1900), .B2(n1908), .A(n1876), .ZN(N2866) );
  AND2_X1 U1020 ( .A1(DATA_IN[0]), .A2(n1270), .ZN(n1917) );
  AND2_X1 U1021 ( .A1(DATA_IN[1]), .A2(n1270), .ZN(n1918) );
  AND2_X1 U1022 ( .A1(DATA_IN[2]), .A2(n1270), .ZN(n1919) );
  AND2_X1 U1023 ( .A1(DATA_IN[3]), .A2(n1270), .ZN(n1920) );
  AND2_X1 U1024 ( .A1(DATA_IN[4]), .A2(n1270), .ZN(n1921) );
  AND2_X1 U1025 ( .A1(DATA_IN[5]), .A2(n1270), .ZN(n1922) );
  AND2_X1 U1026 ( .A1(DATA_IN[6]), .A2(n1270), .ZN(n1923) );
  AND2_X1 U1027 ( .A1(DATA_IN[7]), .A2(n1270), .ZN(n1924) );
  AND2_X1 U1028 ( .A1(DATA_IN[8]), .A2(n1270), .ZN(n1925) );
  AND2_X1 U1029 ( .A1(DATA_IN[0]), .A2(n1270), .ZN(N3317) );
  AND2_X1 U1030 ( .A1(DATA_IN[1]), .A2(n1270), .ZN(N3319) );
  AND2_X1 U1031 ( .A1(DATA_IN[2]), .A2(n1270), .ZN(N3321) );
  AND2_X1 U1032 ( .A1(DATA_IN[3]), .A2(n1270), .ZN(N3323) );
  AND2_X1 U1033 ( .A1(DATA_IN[4]), .A2(n1270), .ZN(N3325) );
  AND2_X1 U1034 ( .A1(DATA_IN[5]), .A2(n1270), .ZN(N3327) );
  AND2_X1 U1035 ( .A1(DATA_IN[6]), .A2(n1270), .ZN(N3329) );
  AND2_X1 U1036 ( .A1(DATA_IN[7]), .A2(n1270), .ZN(N3331) );
  AND2_X1 U1037 ( .A1(DATA_IN[8]), .A2(n1270), .ZN(N3333) );
  AND2_X1 U1038 ( .A1(DATA_IN[9]), .A2(n1229), .ZN(n1926) );
  AND2_X1 U1039 ( .A1(DATA_IN[10]), .A2(n1229), .ZN(n1927) );
  AND2_X1 U1040 ( .A1(DATA_IN[11]), .A2(n1229), .ZN(n1928) );
  AND2_X1 U1041 ( .A1(DATA_IN[12]), .A2(n1229), .ZN(n1929) );
  AND2_X1 U1042 ( .A1(DATA_IN[13]), .A2(n1229), .ZN(n1930) );
  AND2_X1 U1043 ( .A1(DATA_IN[14]), .A2(n1229), .ZN(n1931) );
  AND2_X1 U1044 ( .A1(DATA_IN[15]), .A2(n1229), .ZN(n1932) );
  AND2_X1 U1045 ( .A1(DATA_IN[16]), .A2(n1229), .ZN(n1933) );
  AND2_X1 U1046 ( .A1(DATA_IN[17]), .A2(n1229), .ZN(n1934) );
  AND2_X1 U1047 ( .A1(DATA_IN[18]), .A2(n1229), .ZN(n1935) );
  AND2_X1 U1048 ( .A1(DATA_IN[19]), .A2(n1229), .ZN(n1936) );
  AND2_X1 U1049 ( .A1(DATA_IN[31]), .A2(n1229), .ZN(n1948) );
  AND2_X1 U1050 ( .A1(DATA_IN[9]), .A2(n1229), .ZN(N3335) );
  AND2_X1 U1051 ( .A1(DATA_IN[10]), .A2(n1229), .ZN(N3337) );
  AND2_X1 U1052 ( .A1(DATA_IN[11]), .A2(n1229), .ZN(N3339) );
  AND2_X1 U1053 ( .A1(DATA_IN[12]), .A2(n1229), .ZN(N3341) );
  AND2_X1 U1054 ( .A1(DATA_IN[13]), .A2(n1229), .ZN(N3343) );
  AND2_X1 U1055 ( .A1(DATA_IN[14]), .A2(n1229), .ZN(N3345) );
  AND2_X1 U1056 ( .A1(DATA_IN[15]), .A2(n1229), .ZN(N3347) );
  AND2_X1 U1057 ( .A1(DATA_IN[16]), .A2(n1229), .ZN(N3349) );
  AND2_X1 U1058 ( .A1(DATA_IN[17]), .A2(n1229), .ZN(N3351) );
  AND2_X1 U1059 ( .A1(DATA_IN[18]), .A2(n1229), .ZN(N3353) );
  AND2_X1 U1060 ( .A1(DATA_IN[20]), .A2(n1229), .ZN(N3357) );
  AND2_X1 U1061 ( .A1(DATA_IN[31]), .A2(n1229), .ZN(N3379) );
  AND2_X1 U1062 ( .A1(DATA_IN[20]), .A2(n1), .ZN(n1937) );
  AND2_X1 U1063 ( .A1(DATA_IN[21]), .A2(n1), .ZN(n1938) );
  AND2_X1 U1064 ( .A1(DATA_IN[22]), .A2(n1), .ZN(n1939) );
  AND2_X1 U1065 ( .A1(DATA_IN[23]), .A2(n1), .ZN(n1940) );
  AND2_X1 U1066 ( .A1(DATA_IN[24]), .A2(n1), .ZN(n1941) );
  AND2_X1 U1067 ( .A1(DATA_IN[25]), .A2(n1), .ZN(n1942) );
  AND2_X1 U1068 ( .A1(DATA_IN[26]), .A2(n1), .ZN(n1943) );
  AND2_X1 U1069 ( .A1(DATA_IN[27]), .A2(n1), .ZN(n1944) );
  AND2_X1 U1070 ( .A1(DATA_IN[28]), .A2(n1), .ZN(n1945) );
  AND2_X1 U1071 ( .A1(DATA_IN[29]), .A2(n1), .ZN(n1946) );
  AND2_X1 U1072 ( .A1(DATA_IN[30]), .A2(n1), .ZN(n1947) );
  AND2_X1 U1073 ( .A1(DATA_IN[19]), .A2(n1), .ZN(N3355) );
  AND2_X1 U1074 ( .A1(DATA_IN[21]), .A2(n1), .ZN(N3359) );
  AND2_X1 U1075 ( .A1(DATA_IN[22]), .A2(n1), .ZN(N3361) );
  AND2_X1 U1076 ( .A1(DATA_IN[23]), .A2(n1), .ZN(N3363) );
  AND2_X1 U1077 ( .A1(DATA_IN[24]), .A2(n1), .ZN(N3365) );
  AND2_X1 U1078 ( .A1(DATA_IN[25]), .A2(n1), .ZN(N3367) );
  AND2_X1 U1079 ( .A1(DATA_IN[26]), .A2(n1), .ZN(N3369) );
  AND2_X1 U1080 ( .A1(DATA_IN[27]), .A2(n1), .ZN(N3371) );
  AND2_X1 U1081 ( .A1(DATA_IN[28]), .A2(n1), .ZN(N3373) );
  AND2_X1 U1082 ( .A1(DATA_IN[29]), .A2(n1), .ZN(N3375) );
  AND2_X1 U1083 ( .A1(DATA_IN[30]), .A2(n1), .ZN(N3377) );
  OAI221_X1 U1084 ( .B1(n2172), .B2(n90), .C1(n2169), .C2(n91), .A(n92), .ZN(
        n77) );
  AOI222_X1 U1085 ( .A1(\REGISTERS[21][1] ), .A2(n2168), .B1(
        \REGISTERS[20][1] ), .B2(n2165), .C1(\REGISTERS[16][1] ), .C2(n2164), 
        .ZN(n92) );
  OAI221_X1 U1086 ( .B1(n2172), .B2(n128), .C1(n2169), .C2(n129), .A(n130), 
        .ZN(n115) );
  AOI222_X1 U1087 ( .A1(\REGISTERS[21][2] ), .A2(n2168), .B1(
        \REGISTERS[20][2] ), .B2(n2165), .C1(\REGISTERS[16][2] ), .C2(n2164), 
        .ZN(n130) );
  OAI221_X1 U1088 ( .B1(n2172), .B2(n166), .C1(n2169), .C2(n167), .A(n168), 
        .ZN(n153) );
  AOI222_X1 U1089 ( .A1(\REGISTERS[21][3] ), .A2(n2168), .B1(
        \REGISTERS[20][3] ), .B2(n2165), .C1(\REGISTERS[16][3] ), .C2(n2164), 
        .ZN(n168) );
  OAI221_X1 U1090 ( .B1(n2172), .B2(n204), .C1(n2169), .C2(n205), .A(n206), 
        .ZN(n191) );
  AOI222_X1 U1091 ( .A1(\REGISTERS[21][4] ), .A2(n2168), .B1(
        \REGISTERS[20][4] ), .B2(n2165), .C1(\REGISTERS[16][4] ), .C2(n2164), 
        .ZN(n206) );
  OAI221_X1 U1092 ( .B1(n2172), .B2(n242), .C1(n2169), .C2(n243), .A(n244), 
        .ZN(n229) );
  AOI222_X1 U1093 ( .A1(\REGISTERS[21][5] ), .A2(n2168), .B1(
        \REGISTERS[20][5] ), .B2(n2165), .C1(\REGISTERS[16][5] ), .C2(n2164), 
        .ZN(n244) );
  AOI222_X1 U1094 ( .A1(n2069), .A2(\REGISTERS[21][1] ), .B1(n2066), .B2(
        \REGISTERS[20][1] ), .C1(n2065), .C2(\REGISTERS[16][1] ), .ZN(n1333)
         );
  NOR3_X1 U1095 ( .A1(ADDR_RD2[1]), .A2(ADDR_RD2[2]), .A3(n67), .ZN(n1227) );
  NOR3_X1 U1096 ( .A1(n1259), .A2(ADDR_RD2[4]), .A3(n1262), .ZN(n1224) );
  NOR3_X1 U1097 ( .A1(ADDR_RD2[3]), .A2(ADDR_RD2[4]), .A3(n1259), .ZN(n1234)
         );
  NOR3_X1 U1098 ( .A1(n1894), .A2(ADDR_RD1[4]), .A3(n1895), .ZN(n1871) );
  NOR3_X1 U1099 ( .A1(ADDR_RD1[3]), .A2(ADDR_RD1[4]), .A3(n1894), .ZN(n1879)
         );
  NOR3_X1 U1100 ( .A1(ADDR_RD2[0]), .A2(ADDR_RD2[4]), .A3(n1262), .ZN(n1226)
         );
  NOR3_X1 U1101 ( .A1(ADDR_RD2[3]), .A2(ADDR_RD2[4]), .A3(ADDR_RD2[0]), .ZN(
        n1235) );
  NOR3_X1 U1102 ( .A1(ADDR_RD1[0]), .A2(ADDR_RD1[4]), .A3(n1895), .ZN(n1873)
         );
  NOR3_X1 U1103 ( .A1(ADDR_RD1[3]), .A2(ADDR_RD1[4]), .A3(ADDR_RD1[0]), .ZN(
        n1880) );
  NOR2_X1 U1104 ( .A1(n1269), .A2(ADDR_RD2[2]), .ZN(n1230) );
  NOR2_X1 U1105 ( .A1(n1898), .A2(ADDR_RD1[2]), .ZN(n1877) );
  OAI221_X1 U1106 ( .B1(n2174), .B2(n1040), .C1(n2171), .C2(n1041), .A(n1042), 
        .ZN(n1027) );
  AOI222_X1 U1107 ( .A1(\REGISTERS[21][26] ), .A2(n2166), .B1(
        \REGISTERS[20][26] ), .B2(n2165), .C1(\REGISTERS[16][26] ), .C2(n2162), 
        .ZN(n1042) );
  OAI221_X1 U1108 ( .B1(n2174), .B2(n1078), .C1(n2171), .C2(n1079), .A(n1080), 
        .ZN(n1065) );
  AOI222_X1 U1109 ( .A1(\REGISTERS[21][27] ), .A2(n2166), .B1(
        \REGISTERS[20][27] ), .B2(n2165), .C1(\REGISTERS[16][27] ), .C2(n2162), 
        .ZN(n1080) );
  OAI221_X1 U1110 ( .B1(n2174), .B2(n1116), .C1(n2171), .C2(n1117), .A(n1118), 
        .ZN(n1103) );
  AOI222_X1 U1111 ( .A1(\REGISTERS[21][28] ), .A2(n2166), .B1(
        \REGISTERS[20][28] ), .B2(n2165), .C1(\REGISTERS[16][28] ), .C2(n2162), 
        .ZN(n1118) );
  OAI221_X1 U1112 ( .B1(n2174), .B2(n1154), .C1(n2171), .C2(n1155), .A(n1156), 
        .ZN(n1141) );
  AOI222_X1 U1113 ( .A1(\REGISTERS[21][29] ), .A2(n2166), .B1(
        \REGISTERS[20][29] ), .B2(n2165), .C1(\REGISTERS[16][29] ), .C2(n2162), 
        .ZN(n1156) );
  OAI221_X1 U1114 ( .B1(n2174), .B2(n1192), .C1(n2171), .C2(n1193), .A(n1194), 
        .ZN(n1179) );
  AOI222_X1 U1115 ( .A1(\REGISTERS[21][30] ), .A2(n2166), .B1(
        \REGISTERS[20][30] ), .B2(n2165), .C1(\REGISTERS[16][30] ), .C2(n2162), 
        .ZN(n1194) );
  OAI221_X1 U1116 ( .B1(n2174), .B2(n1242), .C1(n2171), .C2(n1243), .A(n1244), 
        .ZN(n1217) );
  AOI222_X1 U1117 ( .A1(\REGISTERS[21][31] ), .A2(n2166), .B1(
        \REGISTERS[20][31] ), .B2(n2165), .C1(\REGISTERS[16][31] ), .C2(n2162), 
        .ZN(n1244) );
  OAI221_X1 U1118 ( .B1(n1040), .B2(n2075), .C1(n1041), .C2(n2072), .A(n1783), 
        .ZN(n1776) );
  AOI222_X1 U1119 ( .A1(n2067), .A2(\REGISTERS[21][26] ), .B1(n2066), .B2(
        \REGISTERS[20][26] ), .C1(n2063), .C2(\REGISTERS[16][26] ), .ZN(n1783)
         );
  OAI221_X1 U1120 ( .B1(n1078), .B2(n2075), .C1(n1079), .C2(n2072), .A(n1801), 
        .ZN(n1794) );
  AOI222_X1 U1121 ( .A1(n2067), .A2(\REGISTERS[21][27] ), .B1(n2066), .B2(
        \REGISTERS[20][27] ), .C1(n2063), .C2(\REGISTERS[16][27] ), .ZN(n1801)
         );
  OAI221_X1 U1122 ( .B1(n1116), .B2(n2075), .C1(n1117), .C2(n2072), .A(n1819), 
        .ZN(n1812) );
  AOI222_X1 U1123 ( .A1(n2067), .A2(\REGISTERS[21][28] ), .B1(n2066), .B2(
        \REGISTERS[20][28] ), .C1(n2063), .C2(\REGISTERS[16][28] ), .ZN(n1819)
         );
  OAI221_X1 U1124 ( .B1(n1154), .B2(n2075), .C1(n1155), .C2(n2072), .A(n1837), 
        .ZN(n1830) );
  AOI222_X1 U1125 ( .A1(n2067), .A2(\REGISTERS[21][29] ), .B1(n2066), .B2(
        \REGISTERS[20][29] ), .C1(n2063), .C2(\REGISTERS[16][29] ), .ZN(n1837)
         );
  OAI221_X1 U1126 ( .B1(n1192), .B2(n2075), .C1(n1193), .C2(n2072), .A(n1855), 
        .ZN(n1848) );
  AOI222_X1 U1127 ( .A1(n2067), .A2(\REGISTERS[21][30] ), .B1(n2066), .B2(
        \REGISTERS[20][30] ), .C1(n2063), .C2(\REGISTERS[16][30] ), .ZN(n1855)
         );
  OAI221_X1 U1128 ( .B1(n1242), .B2(n2075), .C1(n1243), .C2(n2072), .A(n1885), 
        .ZN(n1866) );
  AOI222_X1 U1129 ( .A1(n2067), .A2(\REGISTERS[21][31] ), .B1(n2066), .B2(
        \REGISTERS[20][31] ), .C1(n2063), .C2(\REGISTERS[16][31] ), .ZN(n1885)
         );
  OAI221_X1 U1130 ( .B1(n2172), .B2(n280), .C1(n2169), .C2(n281), .A(n282), 
        .ZN(n267) );
  AOI222_X1 U1131 ( .A1(\REGISTERS[21][6] ), .A2(n2167), .B1(
        \REGISTERS[20][6] ), .B2(n2165), .C1(\REGISTERS[16][6] ), .C2(n2163), 
        .ZN(n282) );
  OAI221_X1 U1132 ( .B1(n2172), .B2(n318), .C1(n2169), .C2(n319), .A(n320), 
        .ZN(n305) );
  AOI222_X1 U1133 ( .A1(\REGISTERS[21][7] ), .A2(n2167), .B1(
        \REGISTERS[20][7] ), .B2(n2165), .C1(\REGISTERS[16][7] ), .C2(n2163), 
        .ZN(n320) );
  OAI221_X1 U1134 ( .B1(n2172), .B2(n356), .C1(n2169), .C2(n357), .A(n358), 
        .ZN(n343) );
  AOI222_X1 U1135 ( .A1(\REGISTERS[21][8] ), .A2(n2167), .B1(
        \REGISTERS[20][8] ), .B2(n2165), .C1(\REGISTERS[16][8] ), .C2(n2163), 
        .ZN(n358) );
  OAI221_X1 U1136 ( .B1(n2172), .B2(n394), .C1(n2169), .C2(n395), .A(n396), 
        .ZN(n381) );
  AOI222_X1 U1137 ( .A1(\REGISTERS[21][9] ), .A2(n2167), .B1(
        \REGISTERS[20][9] ), .B2(n2165), .C1(\REGISTERS[16][9] ), .C2(n2163), 
        .ZN(n396) );
  OAI221_X1 U1138 ( .B1(n2172), .B2(n432), .C1(n2169), .C2(n433), .A(n434), 
        .ZN(n419) );
  AOI222_X1 U1139 ( .A1(\REGISTERS[21][10] ), .A2(n2167), .B1(
        \REGISTERS[20][10] ), .B2(n2165), .C1(\REGISTERS[16][10] ), .C2(n2163), 
        .ZN(n434) );
  OAI221_X1 U1140 ( .B1(n2172), .B2(n470), .C1(n2169), .C2(n471), .A(n472), 
        .ZN(n457) );
  AOI222_X1 U1141 ( .A1(\REGISTERS[21][11] ), .A2(n2167), .B1(
        \REGISTERS[20][11] ), .B2(n2165), .C1(\REGISTERS[16][11] ), .C2(n2163), 
        .ZN(n472) );
  OAI221_X1 U1142 ( .B1(n2172), .B2(n508), .C1(n2169), .C2(n509), .A(n510), 
        .ZN(n495) );
  AOI222_X1 U1143 ( .A1(\REGISTERS[21][12] ), .A2(n2167), .B1(
        \REGISTERS[20][12] ), .B2(n2165), .C1(\REGISTERS[16][12] ), .C2(n2163), 
        .ZN(n510) );
  OAI221_X1 U1144 ( .B1(n2173), .B2(n546), .C1(n2170), .C2(n547), .A(n548), 
        .ZN(n533) );
  AOI222_X1 U1145 ( .A1(\REGISTERS[21][13] ), .A2(n2167), .B1(
        \REGISTERS[20][13] ), .B2(n2165), .C1(\REGISTERS[16][13] ), .C2(n2163), 
        .ZN(n548) );
  OAI221_X1 U1146 ( .B1(n2173), .B2(n584), .C1(n2170), .C2(n585), .A(n586), 
        .ZN(n571) );
  AOI222_X1 U1147 ( .A1(\REGISTERS[21][14] ), .A2(n2167), .B1(
        \REGISTERS[20][14] ), .B2(n2165), .C1(\REGISTERS[16][14] ), .C2(n2163), 
        .ZN(n586) );
  OAI221_X1 U1148 ( .B1(n2173), .B2(n622), .C1(n2170), .C2(n623), .A(n624), 
        .ZN(n609) );
  AOI222_X1 U1149 ( .A1(\REGISTERS[21][15] ), .A2(n2167), .B1(
        \REGISTERS[20][15] ), .B2(n2165), .C1(\REGISTERS[16][15] ), .C2(n2163), 
        .ZN(n624) );
  OAI221_X1 U1150 ( .B1(n2173), .B2(n660), .C1(n2170), .C2(n661), .A(n662), 
        .ZN(n647) );
  AOI222_X1 U1151 ( .A1(\REGISTERS[21][16] ), .A2(n2167), .B1(
        \REGISTERS[20][16] ), .B2(n2165), .C1(\REGISTERS[16][16] ), .C2(n2163), 
        .ZN(n662) );
  OAI221_X1 U1152 ( .B1(n2173), .B2(n698), .C1(n2170), .C2(n699), .A(n700), 
        .ZN(n685) );
  AOI222_X1 U1153 ( .A1(\REGISTERS[21][17] ), .A2(n2167), .B1(
        \REGISTERS[20][17] ), .B2(n2165), .C1(\REGISTERS[16][17] ), .C2(n2163), 
        .ZN(n700) );
  OAI221_X1 U1154 ( .B1(n2173), .B2(n736), .C1(n2170), .C2(n737), .A(n738), 
        .ZN(n723) );
  AOI222_X1 U1155 ( .A1(\REGISTERS[21][18] ), .A2(n2167), .B1(
        \REGISTERS[20][18] ), .B2(n2165), .C1(\REGISTERS[16][18] ), .C2(n2163), 
        .ZN(n738) );
  OAI221_X1 U1156 ( .B1(n2173), .B2(n774), .C1(n2170), .C2(n775), .A(n776), 
        .ZN(n761) );
  AOI222_X1 U1157 ( .A1(\REGISTERS[21][19] ), .A2(n2166), .B1(
        \REGISTERS[20][19] ), .B2(n2165), .C1(\REGISTERS[16][19] ), .C2(n2162), 
        .ZN(n776) );
  OAI221_X1 U1158 ( .B1(n2173), .B2(n812), .C1(n2170), .C2(n813), .A(n814), 
        .ZN(n799) );
  AOI222_X1 U1159 ( .A1(\REGISTERS[21][20] ), .A2(n2166), .B1(
        \REGISTERS[20][20] ), .B2(n2165), .C1(\REGISTERS[16][20] ), .C2(n2162), 
        .ZN(n814) );
  OAI221_X1 U1160 ( .B1(n2173), .B2(n850), .C1(n2170), .C2(n851), .A(n852), 
        .ZN(n837) );
  AOI222_X1 U1161 ( .A1(\REGISTERS[21][21] ), .A2(n2166), .B1(
        \REGISTERS[20][21] ), .B2(n2165), .C1(\REGISTERS[16][21] ), .C2(n2162), 
        .ZN(n852) );
  OAI221_X1 U1162 ( .B1(n2173), .B2(n888), .C1(n2170), .C2(n889), .A(n890), 
        .ZN(n875) );
  AOI222_X1 U1163 ( .A1(\REGISTERS[21][22] ), .A2(n2166), .B1(
        \REGISTERS[20][22] ), .B2(n2165), .C1(\REGISTERS[16][22] ), .C2(n2162), 
        .ZN(n890) );
  OAI221_X1 U1164 ( .B1(n2173), .B2(n926), .C1(n2170), .C2(n927), .A(n928), 
        .ZN(n913) );
  AOI222_X1 U1165 ( .A1(\REGISTERS[21][23] ), .A2(n2166), .B1(
        \REGISTERS[20][23] ), .B2(n2165), .C1(\REGISTERS[16][23] ), .C2(n2162), 
        .ZN(n928) );
  OAI221_X1 U1166 ( .B1(n2173), .B2(n964), .C1(n2170), .C2(n965), .A(n966), 
        .ZN(n951) );
  AOI222_X1 U1167 ( .A1(\REGISTERS[21][24] ), .A2(n2166), .B1(
        \REGISTERS[20][24] ), .B2(n2165), .C1(\REGISTERS[16][24] ), .C2(n2162), 
        .ZN(n966) );
  OAI221_X1 U1168 ( .B1(n2173), .B2(n1002), .C1(n2170), .C2(n1003), .A(n1004), 
        .ZN(n989) );
  AOI222_X1 U1169 ( .A1(\REGISTERS[21][25] ), .A2(n2166), .B1(
        \REGISTERS[20][25] ), .B2(n2165), .C1(\REGISTERS[16][25] ), .C2(n2162), 
        .ZN(n1004) );
  OAI221_X1 U1170 ( .B1(n32), .B2(n2073), .C1(n34), .C2(n2070), .A(n1296), 
        .ZN(n1275) );
  AOI222_X1 U1171 ( .A1(n2069), .A2(\REGISTERS[21][0] ), .B1(n2066), .B2(
        \REGISTERS[20][0] ), .C1(n2065), .C2(\REGISTERS[16][0] ), .ZN(n1296)
         );
  OAI221_X1 U1172 ( .B1(n128), .B2(n2073), .C1(n129), .C2(n2070), .A(n1351), 
        .ZN(n1344) );
  AOI222_X1 U1173 ( .A1(n2069), .A2(\REGISTERS[21][2] ), .B1(n2066), .B2(
        \REGISTERS[20][2] ), .C1(n2065), .C2(\REGISTERS[16][2] ), .ZN(n1351)
         );
  OAI221_X1 U1174 ( .B1(n166), .B2(n2073), .C1(n167), .C2(n2070), .A(n1369), 
        .ZN(n1362) );
  AOI222_X1 U1175 ( .A1(n2069), .A2(\REGISTERS[21][3] ), .B1(n2066), .B2(
        \REGISTERS[20][3] ), .C1(n2065), .C2(\REGISTERS[16][3] ), .ZN(n1369)
         );
  OAI221_X1 U1176 ( .B1(n204), .B2(n2073), .C1(n205), .C2(n2070), .A(n1387), 
        .ZN(n1380) );
  AOI222_X1 U1177 ( .A1(n2069), .A2(\REGISTERS[21][4] ), .B1(n2066), .B2(
        \REGISTERS[20][4] ), .C1(n2065), .C2(\REGISTERS[16][4] ), .ZN(n1387)
         );
  OAI221_X1 U1178 ( .B1(n242), .B2(n2073), .C1(n243), .C2(n2070), .A(n1405), 
        .ZN(n1398) );
  AOI222_X1 U1179 ( .A1(n2069), .A2(\REGISTERS[21][5] ), .B1(n2066), .B2(
        \REGISTERS[20][5] ), .C1(n2065), .C2(\REGISTERS[16][5] ), .ZN(n1405)
         );
  OAI221_X1 U1180 ( .B1(n280), .B2(n2073), .C1(n281), .C2(n2070), .A(n1423), 
        .ZN(n1416) );
  AOI222_X1 U1181 ( .A1(n2068), .A2(\REGISTERS[21][6] ), .B1(n2066), .B2(
        \REGISTERS[20][6] ), .C1(n2064), .C2(\REGISTERS[16][6] ), .ZN(n1423)
         );
  OAI221_X1 U1182 ( .B1(n318), .B2(n2073), .C1(n319), .C2(n2070), .A(n1441), 
        .ZN(n1434) );
  AOI222_X1 U1183 ( .A1(n2068), .A2(\REGISTERS[21][7] ), .B1(n2066), .B2(
        \REGISTERS[20][7] ), .C1(n2064), .C2(\REGISTERS[16][7] ), .ZN(n1441)
         );
  OAI221_X1 U1184 ( .B1(n356), .B2(n2073), .C1(n357), .C2(n2070), .A(n1459), 
        .ZN(n1452) );
  AOI222_X1 U1185 ( .A1(n2068), .A2(\REGISTERS[21][8] ), .B1(n2066), .B2(
        \REGISTERS[20][8] ), .C1(n2064), .C2(\REGISTERS[16][8] ), .ZN(n1459)
         );
  OAI221_X1 U1186 ( .B1(n394), .B2(n2073), .C1(n395), .C2(n2070), .A(n1477), 
        .ZN(n1470) );
  AOI222_X1 U1187 ( .A1(n2068), .A2(\REGISTERS[21][9] ), .B1(n2066), .B2(
        \REGISTERS[20][9] ), .C1(n2064), .C2(\REGISTERS[16][9] ), .ZN(n1477)
         );
  OAI221_X1 U1188 ( .B1(n432), .B2(n2073), .C1(n433), .C2(n2070), .A(n1495), 
        .ZN(n1488) );
  AOI222_X1 U1189 ( .A1(n2068), .A2(\REGISTERS[21][10] ), .B1(n2066), .B2(
        \REGISTERS[20][10] ), .C1(n2064), .C2(\REGISTERS[16][10] ), .ZN(n1495)
         );
  OAI221_X1 U1190 ( .B1(n470), .B2(n2073), .C1(n471), .C2(n2070), .A(n1513), 
        .ZN(n1506) );
  AOI222_X1 U1191 ( .A1(n2068), .A2(\REGISTERS[21][11] ), .B1(n2066), .B2(
        \REGISTERS[20][11] ), .C1(n2064), .C2(\REGISTERS[16][11] ), .ZN(n1513)
         );
  OAI221_X1 U1192 ( .B1(n508), .B2(n2073), .C1(n509), .C2(n2070), .A(n1531), 
        .ZN(n1524) );
  AOI222_X1 U1193 ( .A1(n2068), .A2(\REGISTERS[21][12] ), .B1(n2066), .B2(
        \REGISTERS[20][12] ), .C1(n2064), .C2(\REGISTERS[16][12] ), .ZN(n1531)
         );
  OAI221_X1 U1194 ( .B1(n546), .B2(n2074), .C1(n547), .C2(n2071), .A(n1549), 
        .ZN(n1542) );
  AOI222_X1 U1195 ( .A1(n2068), .A2(\REGISTERS[21][13] ), .B1(n2066), .B2(
        \REGISTERS[20][13] ), .C1(n2064), .C2(\REGISTERS[16][13] ), .ZN(n1549)
         );
  OAI221_X1 U1196 ( .B1(n584), .B2(n2074), .C1(n585), .C2(n2071), .A(n1567), 
        .ZN(n1560) );
  AOI222_X1 U1197 ( .A1(n2068), .A2(\REGISTERS[21][14] ), .B1(n2066), .B2(
        \REGISTERS[20][14] ), .C1(n2064), .C2(\REGISTERS[16][14] ), .ZN(n1567)
         );
  OAI221_X1 U1198 ( .B1(n622), .B2(n2074), .C1(n623), .C2(n2071), .A(n1585), 
        .ZN(n1578) );
  AOI222_X1 U1199 ( .A1(n2068), .A2(\REGISTERS[21][15] ), .B1(n2066), .B2(
        \REGISTERS[20][15] ), .C1(n2064), .C2(\REGISTERS[16][15] ), .ZN(n1585)
         );
  OAI221_X1 U1200 ( .B1(n660), .B2(n2074), .C1(n661), .C2(n2071), .A(n1603), 
        .ZN(n1596) );
  AOI222_X1 U1201 ( .A1(n2068), .A2(\REGISTERS[21][16] ), .B1(n2066), .B2(
        \REGISTERS[20][16] ), .C1(n2064), .C2(\REGISTERS[16][16] ), .ZN(n1603)
         );
  OAI221_X1 U1202 ( .B1(n698), .B2(n2074), .C1(n699), .C2(n2071), .A(n1621), 
        .ZN(n1614) );
  AOI222_X1 U1203 ( .A1(n2068), .A2(\REGISTERS[21][17] ), .B1(n2066), .B2(
        \REGISTERS[20][17] ), .C1(n2064), .C2(\REGISTERS[16][17] ), .ZN(n1621)
         );
  OAI221_X1 U1204 ( .B1(n736), .B2(n2074), .C1(n737), .C2(n2071), .A(n1639), 
        .ZN(n1632) );
  AOI222_X1 U1205 ( .A1(n2068), .A2(\REGISTERS[21][18] ), .B1(n2066), .B2(
        \REGISTERS[20][18] ), .C1(n2064), .C2(\REGISTERS[16][18] ), .ZN(n1639)
         );
  OAI221_X1 U1206 ( .B1(n774), .B2(n2074), .C1(n775), .C2(n2071), .A(n1657), 
        .ZN(n1650) );
  AOI222_X1 U1207 ( .A1(n2067), .A2(\REGISTERS[21][19] ), .B1(n2066), .B2(
        \REGISTERS[20][19] ), .C1(n2063), .C2(\REGISTERS[16][19] ), .ZN(n1657)
         );
  OAI221_X1 U1208 ( .B1(n812), .B2(n2074), .C1(n813), .C2(n2071), .A(n1675), 
        .ZN(n1668) );
  AOI222_X1 U1209 ( .A1(n2067), .A2(\REGISTERS[21][20] ), .B1(n2066), .B2(
        \REGISTERS[20][20] ), .C1(n2063), .C2(\REGISTERS[16][20] ), .ZN(n1675)
         );
  OAI221_X1 U1210 ( .B1(n850), .B2(n2074), .C1(n851), .C2(n2071), .A(n1693), 
        .ZN(n1686) );
  AOI222_X1 U1211 ( .A1(n2067), .A2(\REGISTERS[21][21] ), .B1(n2066), .B2(
        \REGISTERS[20][21] ), .C1(n2063), .C2(\REGISTERS[16][21] ), .ZN(n1693)
         );
  OAI221_X1 U1212 ( .B1(n888), .B2(n2074), .C1(n889), .C2(n2071), .A(n1711), 
        .ZN(n1704) );
  AOI222_X1 U1213 ( .A1(n2067), .A2(\REGISTERS[21][22] ), .B1(n2066), .B2(
        \REGISTERS[20][22] ), .C1(n2063), .C2(\REGISTERS[16][22] ), .ZN(n1711)
         );
  OAI221_X1 U1214 ( .B1(n926), .B2(n2074), .C1(n927), .C2(n2071), .A(n1729), 
        .ZN(n1722) );
  AOI222_X1 U1215 ( .A1(n2067), .A2(\REGISTERS[21][23] ), .B1(n2066), .B2(
        \REGISTERS[20][23] ), .C1(n2063), .C2(\REGISTERS[16][23] ), .ZN(n1729)
         );
  OAI221_X1 U1216 ( .B1(n964), .B2(n2074), .C1(n965), .C2(n2071), .A(n1747), 
        .ZN(n1740) );
  AOI222_X1 U1217 ( .A1(n2067), .A2(\REGISTERS[21][24] ), .B1(n2066), .B2(
        \REGISTERS[20][24] ), .C1(n2063), .C2(\REGISTERS[16][24] ), .ZN(n1747)
         );
  OAI221_X1 U1218 ( .B1(n1002), .B2(n2074), .C1(n1003), .C2(n2071), .A(n1765), 
        .ZN(n1758) );
  AOI222_X1 U1219 ( .A1(n2067), .A2(\REGISTERS[21][25] ), .B1(n2066), .B2(
        \REGISTERS[20][25] ), .C1(n2063), .C2(\REGISTERS[16][25] ), .ZN(n1765)
         );
  AOI22_X1 U1220 ( .A1(\REGISTERS[8][0] ), .A2(n2204), .B1(\REGISTERS[13][0] ), 
        .B2(n2201), .ZN(n14) );
  AOI22_X1 U1221 ( .A1(\REGISTERS[0][0] ), .A2(n2192), .B1(\REGISTERS[5][0] ), 
        .B2(n2189), .ZN(n21) );
  AOI22_X1 U1222 ( .A1(\REGISTERS[24][0] ), .A2(n2180), .B1(\REGISTERS[31][0] ), .B2(n2177), .ZN(n28) );
  AOI22_X1 U1223 ( .A1(\REGISTERS[8][1] ), .A2(n2204), .B1(\REGISTERS[13][1] ), 
        .B2(n2201), .ZN(n83) );
  AOI22_X1 U1224 ( .A1(\REGISTERS[0][1] ), .A2(n2192), .B1(\REGISTERS[5][1] ), 
        .B2(n2189), .ZN(n86) );
  AOI22_X1 U1225 ( .A1(\REGISTERS[24][1] ), .A2(n2180), .B1(\REGISTERS[31][1] ), .B2(n2177), .ZN(n89) );
  AOI22_X1 U1226 ( .A1(\REGISTERS[8][2] ), .A2(n2204), .B1(\REGISTERS[13][2] ), 
        .B2(n2201), .ZN(n121) );
  AOI22_X1 U1227 ( .A1(\REGISTERS[0][2] ), .A2(n2192), .B1(\REGISTERS[5][2] ), 
        .B2(n2189), .ZN(n124) );
  AOI22_X1 U1228 ( .A1(\REGISTERS[24][2] ), .A2(n2180), .B1(\REGISTERS[31][2] ), .B2(n2177), .ZN(n127) );
  AOI22_X1 U1229 ( .A1(\REGISTERS[8][3] ), .A2(n2204), .B1(\REGISTERS[13][3] ), 
        .B2(n2201), .ZN(n159) );
  AOI22_X1 U1230 ( .A1(\REGISTERS[0][3] ), .A2(n2192), .B1(\REGISTERS[5][3] ), 
        .B2(n2189), .ZN(n162) );
  AOI22_X1 U1231 ( .A1(\REGISTERS[24][3] ), .A2(n2180), .B1(\REGISTERS[31][3] ), .B2(n2177), .ZN(n165) );
  AOI22_X1 U1232 ( .A1(\REGISTERS[8][4] ), .A2(n2204), .B1(\REGISTERS[13][4] ), 
        .B2(n2201), .ZN(n197) );
  AOI22_X1 U1233 ( .A1(\REGISTERS[0][4] ), .A2(n2192), .B1(\REGISTERS[5][4] ), 
        .B2(n2189), .ZN(n200) );
  AOI22_X1 U1234 ( .A1(\REGISTERS[24][4] ), .A2(n2180), .B1(\REGISTERS[31][4] ), .B2(n2177), .ZN(n203) );
  AOI22_X1 U1235 ( .A1(\REGISTERS[8][5] ), .A2(n2204), .B1(\REGISTERS[13][5] ), 
        .B2(n2201), .ZN(n235) );
  AOI22_X1 U1236 ( .A1(\REGISTERS[0][5] ), .A2(n2192), .B1(\REGISTERS[5][5] ), 
        .B2(n2189), .ZN(n238) );
  AOI22_X1 U1237 ( .A1(\REGISTERS[24][5] ), .A2(n2180), .B1(\REGISTERS[31][5] ), .B2(n2177), .ZN(n241) );
  AOI22_X1 U1238 ( .A1(\REGISTERS[8][6] ), .A2(n2203), .B1(\REGISTERS[13][6] ), 
        .B2(n2200), .ZN(n273) );
  AOI22_X1 U1239 ( .A1(\REGISTERS[0][6] ), .A2(n2191), .B1(\REGISTERS[5][6] ), 
        .B2(n2188), .ZN(n276) );
  AOI22_X1 U1240 ( .A1(\REGISTERS[24][6] ), .A2(n2179), .B1(\REGISTERS[31][6] ), .B2(n2176), .ZN(n279) );
  AOI22_X1 U1241 ( .A1(\REGISTERS[8][7] ), .A2(n2203), .B1(\REGISTERS[13][7] ), 
        .B2(n2200), .ZN(n311) );
  AOI22_X1 U1242 ( .A1(\REGISTERS[0][7] ), .A2(n2191), .B1(\REGISTERS[5][7] ), 
        .B2(n2188), .ZN(n314) );
  AOI22_X1 U1243 ( .A1(\REGISTERS[24][7] ), .A2(n2179), .B1(\REGISTERS[31][7] ), .B2(n2176), .ZN(n317) );
  AOI22_X1 U1244 ( .A1(\REGISTERS[8][8] ), .A2(n2203), .B1(\REGISTERS[13][8] ), 
        .B2(n2200), .ZN(n349) );
  AOI22_X1 U1245 ( .A1(\REGISTERS[0][8] ), .A2(n2191), .B1(\REGISTERS[5][8] ), 
        .B2(n2188), .ZN(n352) );
  AOI22_X1 U1246 ( .A1(\REGISTERS[24][8] ), .A2(n2179), .B1(\REGISTERS[31][8] ), .B2(n2176), .ZN(n355) );
  AOI22_X1 U1247 ( .A1(\REGISTERS[8][9] ), .A2(n2203), .B1(\REGISTERS[13][9] ), 
        .B2(n2200), .ZN(n387) );
  AOI22_X1 U1248 ( .A1(\REGISTERS[0][9] ), .A2(n2191), .B1(\REGISTERS[5][9] ), 
        .B2(n2188), .ZN(n390) );
  AOI22_X1 U1249 ( .A1(\REGISTERS[24][9] ), .A2(n2179), .B1(\REGISTERS[31][9] ), .B2(n2176), .ZN(n393) );
  AOI22_X1 U1250 ( .A1(\REGISTERS[8][10] ), .A2(n2203), .B1(
        \REGISTERS[13][10] ), .B2(n2200), .ZN(n425) );
  AOI22_X1 U1251 ( .A1(\REGISTERS[0][10] ), .A2(n2191), .B1(\REGISTERS[5][10] ), .B2(n2188), .ZN(n428) );
  AOI22_X1 U1252 ( .A1(\REGISTERS[24][10] ), .A2(n2179), .B1(
        \REGISTERS[31][10] ), .B2(n2176), .ZN(n431) );
  AOI22_X1 U1253 ( .A1(\REGISTERS[8][11] ), .A2(n2203), .B1(
        \REGISTERS[13][11] ), .B2(n2200), .ZN(n463) );
  AOI22_X1 U1254 ( .A1(\REGISTERS[0][11] ), .A2(n2191), .B1(\REGISTERS[5][11] ), .B2(n2188), .ZN(n466) );
  AOI22_X1 U1255 ( .A1(\REGISTERS[24][11] ), .A2(n2179), .B1(
        \REGISTERS[31][11] ), .B2(n2176), .ZN(n469) );
  AOI22_X1 U1256 ( .A1(\REGISTERS[8][12] ), .A2(n2203), .B1(
        \REGISTERS[13][12] ), .B2(n2200), .ZN(n501) );
  AOI22_X1 U1257 ( .A1(\REGISTERS[0][12] ), .A2(n2191), .B1(\REGISTERS[5][12] ), .B2(n2188), .ZN(n504) );
  AOI22_X1 U1258 ( .A1(\REGISTERS[24][12] ), .A2(n2179), .B1(
        \REGISTERS[31][12] ), .B2(n2176), .ZN(n507) );
  AOI22_X1 U1259 ( .A1(\REGISTERS[8][13] ), .A2(n2203), .B1(
        \REGISTERS[13][13] ), .B2(n2200), .ZN(n539) );
  AOI22_X1 U1260 ( .A1(\REGISTERS[0][13] ), .A2(n2191), .B1(\REGISTERS[5][13] ), .B2(n2188), .ZN(n542) );
  AOI22_X1 U1261 ( .A1(\REGISTERS[24][13] ), .A2(n2179), .B1(
        \REGISTERS[31][13] ), .B2(n2176), .ZN(n545) );
  AOI22_X1 U1262 ( .A1(\REGISTERS[8][14] ), .A2(n2203), .B1(
        \REGISTERS[13][14] ), .B2(n2200), .ZN(n577) );
  AOI22_X1 U1263 ( .A1(\REGISTERS[0][14] ), .A2(n2191), .B1(\REGISTERS[5][14] ), .B2(n2188), .ZN(n580) );
  AOI22_X1 U1264 ( .A1(\REGISTERS[24][14] ), .A2(n2179), .B1(
        \REGISTERS[31][14] ), .B2(n2176), .ZN(n583) );
  AOI22_X1 U1265 ( .A1(\REGISTERS[8][15] ), .A2(n2203), .B1(
        \REGISTERS[13][15] ), .B2(n2200), .ZN(n615) );
  AOI22_X1 U1266 ( .A1(\REGISTERS[0][15] ), .A2(n2191), .B1(\REGISTERS[5][15] ), .B2(n2188), .ZN(n618) );
  AOI22_X1 U1267 ( .A1(\REGISTERS[24][15] ), .A2(n2179), .B1(
        \REGISTERS[31][15] ), .B2(n2176), .ZN(n621) );
  AOI22_X1 U1268 ( .A1(\REGISTERS[8][16] ), .A2(n2203), .B1(
        \REGISTERS[13][16] ), .B2(n2200), .ZN(n653) );
  AOI22_X1 U1269 ( .A1(\REGISTERS[0][16] ), .A2(n2191), .B1(\REGISTERS[5][16] ), .B2(n2188), .ZN(n656) );
  AOI22_X1 U1270 ( .A1(\REGISTERS[24][16] ), .A2(n2179), .B1(
        \REGISTERS[31][16] ), .B2(n2176), .ZN(n659) );
  AOI22_X1 U1271 ( .A1(\REGISTERS[8][17] ), .A2(n2203), .B1(
        \REGISTERS[13][17] ), .B2(n2200), .ZN(n691) );
  AOI22_X1 U1272 ( .A1(\REGISTERS[0][17] ), .A2(n2191), .B1(\REGISTERS[5][17] ), .B2(n2188), .ZN(n694) );
  AOI22_X1 U1273 ( .A1(\REGISTERS[24][17] ), .A2(n2179), .B1(
        \REGISTERS[31][17] ), .B2(n2176), .ZN(n697) );
  AOI22_X1 U1274 ( .A1(\REGISTERS[8][18] ), .A2(n2203), .B1(
        \REGISTERS[13][18] ), .B2(n2200), .ZN(n729) );
  AOI22_X1 U1275 ( .A1(\REGISTERS[0][18] ), .A2(n2191), .B1(\REGISTERS[5][18] ), .B2(n2188), .ZN(n732) );
  AOI22_X1 U1276 ( .A1(\REGISTERS[24][18] ), .A2(n2179), .B1(
        \REGISTERS[31][18] ), .B2(n2176), .ZN(n735) );
  AOI22_X1 U1277 ( .A1(\REGISTERS[8][19] ), .A2(n2202), .B1(
        \REGISTERS[13][19] ), .B2(n2199), .ZN(n767) );
  AOI22_X1 U1278 ( .A1(\REGISTERS[0][19] ), .A2(n2190), .B1(\REGISTERS[5][19] ), .B2(n2187), .ZN(n770) );
  AOI22_X1 U1279 ( .A1(\REGISTERS[24][19] ), .A2(n2178), .B1(
        \REGISTERS[31][19] ), .B2(n2175), .ZN(n773) );
  AOI22_X1 U1280 ( .A1(\REGISTERS[8][20] ), .A2(n2202), .B1(
        \REGISTERS[13][20] ), .B2(n2199), .ZN(n805) );
  AOI22_X1 U1281 ( .A1(\REGISTERS[0][20] ), .A2(n2190), .B1(\REGISTERS[5][20] ), .B2(n2187), .ZN(n808) );
  AOI22_X1 U1282 ( .A1(\REGISTERS[24][20] ), .A2(n2178), .B1(
        \REGISTERS[31][20] ), .B2(n2175), .ZN(n811) );
  AOI22_X1 U1283 ( .A1(\REGISTERS[8][21] ), .A2(n2202), .B1(
        \REGISTERS[13][21] ), .B2(n2199), .ZN(n843) );
  AOI22_X1 U1284 ( .A1(\REGISTERS[0][21] ), .A2(n2190), .B1(\REGISTERS[5][21] ), .B2(n2187), .ZN(n846) );
  AOI22_X1 U1285 ( .A1(\REGISTERS[24][21] ), .A2(n2178), .B1(
        \REGISTERS[31][21] ), .B2(n2175), .ZN(n849) );
  AOI22_X1 U1286 ( .A1(\REGISTERS[8][22] ), .A2(n2202), .B1(
        \REGISTERS[13][22] ), .B2(n2199), .ZN(n881) );
  AOI22_X1 U1287 ( .A1(\REGISTERS[0][22] ), .A2(n2190), .B1(\REGISTERS[5][22] ), .B2(n2187), .ZN(n884) );
  AOI22_X1 U1288 ( .A1(\REGISTERS[24][22] ), .A2(n2178), .B1(
        \REGISTERS[31][22] ), .B2(n2175), .ZN(n887) );
  AOI22_X1 U1289 ( .A1(\REGISTERS[8][23] ), .A2(n2202), .B1(
        \REGISTERS[13][23] ), .B2(n2199), .ZN(n919) );
  AOI22_X1 U1290 ( .A1(\REGISTERS[0][23] ), .A2(n2190), .B1(\REGISTERS[5][23] ), .B2(n2187), .ZN(n922) );
  AOI22_X1 U1291 ( .A1(\REGISTERS[24][23] ), .A2(n2178), .B1(
        \REGISTERS[31][23] ), .B2(n2175), .ZN(n925) );
  AOI22_X1 U1292 ( .A1(\REGISTERS[8][24] ), .A2(n2202), .B1(
        \REGISTERS[13][24] ), .B2(n2199), .ZN(n957) );
  AOI22_X1 U1293 ( .A1(\REGISTERS[0][24] ), .A2(n2190), .B1(\REGISTERS[5][24] ), .B2(n2187), .ZN(n960) );
  AOI22_X1 U1294 ( .A1(\REGISTERS[24][24] ), .A2(n2178), .B1(
        \REGISTERS[31][24] ), .B2(n2175), .ZN(n963) );
  AOI22_X1 U1295 ( .A1(\REGISTERS[8][25] ), .A2(n2202), .B1(
        \REGISTERS[13][25] ), .B2(n2199), .ZN(n995) );
  AOI22_X1 U1296 ( .A1(\REGISTERS[0][25] ), .A2(n2190), .B1(\REGISTERS[5][25] ), .B2(n2187), .ZN(n998) );
  AOI22_X1 U1297 ( .A1(\REGISTERS[24][25] ), .A2(n2178), .B1(
        \REGISTERS[31][25] ), .B2(n2175), .ZN(n1001) );
  AOI22_X1 U1298 ( .A1(\REGISTERS[8][26] ), .A2(n2202), .B1(
        \REGISTERS[13][26] ), .B2(n2199), .ZN(n1033) );
  AOI22_X1 U1299 ( .A1(\REGISTERS[0][26] ), .A2(n2190), .B1(\REGISTERS[5][26] ), .B2(n2187), .ZN(n1036) );
  AOI22_X1 U1300 ( .A1(\REGISTERS[24][26] ), .A2(n2178), .B1(
        \REGISTERS[31][26] ), .B2(n2175), .ZN(n1039) );
  AOI22_X1 U1301 ( .A1(\REGISTERS[8][27] ), .A2(n2202), .B1(
        \REGISTERS[13][27] ), .B2(n2199), .ZN(n1071) );
  AOI22_X1 U1302 ( .A1(\REGISTERS[0][27] ), .A2(n2190), .B1(\REGISTERS[5][27] ), .B2(n2187), .ZN(n1074) );
  AOI22_X1 U1303 ( .A1(\REGISTERS[24][27] ), .A2(n2178), .B1(
        \REGISTERS[31][27] ), .B2(n2175), .ZN(n1077) );
  AOI22_X1 U1304 ( .A1(\REGISTERS[8][28] ), .A2(n2202), .B1(
        \REGISTERS[13][28] ), .B2(n2199), .ZN(n1109) );
  AOI22_X1 U1305 ( .A1(\REGISTERS[0][28] ), .A2(n2190), .B1(\REGISTERS[5][28] ), .B2(n2187), .ZN(n1112) );
  AOI22_X1 U1306 ( .A1(\REGISTERS[24][28] ), .A2(n2178), .B1(
        \REGISTERS[31][28] ), .B2(n2175), .ZN(n1115) );
  AOI22_X1 U1307 ( .A1(\REGISTERS[8][29] ), .A2(n2202), .B1(
        \REGISTERS[13][29] ), .B2(n2199), .ZN(n1147) );
  AOI22_X1 U1308 ( .A1(\REGISTERS[0][29] ), .A2(n2190), .B1(\REGISTERS[5][29] ), .B2(n2187), .ZN(n1150) );
  AOI22_X1 U1309 ( .A1(\REGISTERS[24][29] ), .A2(n2178), .B1(
        \REGISTERS[31][29] ), .B2(n2175), .ZN(n1153) );
  AOI22_X1 U1310 ( .A1(\REGISTERS[8][30] ), .A2(n2202), .B1(
        \REGISTERS[13][30] ), .B2(n2199), .ZN(n1185) );
  AOI22_X1 U1311 ( .A1(\REGISTERS[0][30] ), .A2(n2190), .B1(\REGISTERS[5][30] ), .B2(n2187), .ZN(n1188) );
  AOI22_X1 U1312 ( .A1(\REGISTERS[24][30] ), .A2(n2178), .B1(
        \REGISTERS[31][30] ), .B2(n2175), .ZN(n1191) );
  AOI22_X1 U1313 ( .A1(\REGISTERS[8][31] ), .A2(n2202), .B1(
        \REGISTERS[13][31] ), .B2(n2199), .ZN(n1223) );
  AOI22_X1 U1314 ( .A1(\REGISTERS[0][31] ), .A2(n2190), .B1(\REGISTERS[5][31] ), .B2(n2187), .ZN(n1233) );
  AOI22_X1 U1315 ( .A1(\REGISTERS[24][31] ), .A2(n2178), .B1(
        \REGISTERS[31][31] ), .B2(n2175), .ZN(n1238) );
  AOI22_X1 U1316 ( .A1(n2105), .A2(\REGISTERS[8][0] ), .B1(n2102), .B2(
        \REGISTERS[13][0] ), .ZN(n1281) );
  AOI22_X1 U1317 ( .A1(n2093), .A2(\REGISTERS[0][0] ), .B1(n2090), .B2(
        \REGISTERS[5][0] ), .ZN(n1286) );
  AOI22_X1 U1318 ( .A1(n2081), .A2(\REGISTERS[24][0] ), .B1(n2078), .B2(
        \REGISTERS[31][0] ), .ZN(n1291) );
  AOI22_X1 U1319 ( .A1(n2105), .A2(\REGISTERS[8][1] ), .B1(n2102), .B2(
        \REGISTERS[13][1] ), .ZN(n1330) );
  AOI22_X1 U1320 ( .A1(n2093), .A2(\REGISTERS[0][1] ), .B1(n2090), .B2(
        \REGISTERS[5][1] ), .ZN(n1331) );
  AOI22_X1 U1321 ( .A1(n2081), .A2(\REGISTERS[24][1] ), .B1(n2078), .B2(
        \REGISTERS[31][1] ), .ZN(n1332) );
  AOI22_X1 U1322 ( .A1(n2105), .A2(\REGISTERS[8][2] ), .B1(n2102), .B2(
        \REGISTERS[13][2] ), .ZN(n1348) );
  AOI22_X1 U1323 ( .A1(n2093), .A2(\REGISTERS[0][2] ), .B1(n2090), .B2(
        \REGISTERS[5][2] ), .ZN(n1349) );
  AOI22_X1 U1324 ( .A1(n2081), .A2(\REGISTERS[24][2] ), .B1(n2078), .B2(
        \REGISTERS[31][2] ), .ZN(n1350) );
  AOI22_X1 U1325 ( .A1(n2105), .A2(\REGISTERS[8][3] ), .B1(n2102), .B2(
        \REGISTERS[13][3] ), .ZN(n1366) );
  AOI22_X1 U1326 ( .A1(n2093), .A2(\REGISTERS[0][3] ), .B1(n2090), .B2(
        \REGISTERS[5][3] ), .ZN(n1367) );
  AOI22_X1 U1327 ( .A1(n2081), .A2(\REGISTERS[24][3] ), .B1(n2078), .B2(
        \REGISTERS[31][3] ), .ZN(n1368) );
  AOI22_X1 U1328 ( .A1(n2105), .A2(\REGISTERS[8][4] ), .B1(n2102), .B2(
        \REGISTERS[13][4] ), .ZN(n1384) );
  AOI22_X1 U1329 ( .A1(n2093), .A2(\REGISTERS[0][4] ), .B1(n2090), .B2(
        \REGISTERS[5][4] ), .ZN(n1385) );
  AOI22_X1 U1330 ( .A1(n2081), .A2(\REGISTERS[24][4] ), .B1(n2078), .B2(
        \REGISTERS[31][4] ), .ZN(n1386) );
  AOI22_X1 U1331 ( .A1(n2105), .A2(\REGISTERS[8][5] ), .B1(n2102), .B2(
        \REGISTERS[13][5] ), .ZN(n1402) );
  AOI22_X1 U1332 ( .A1(n2093), .A2(\REGISTERS[0][5] ), .B1(n2090), .B2(
        \REGISTERS[5][5] ), .ZN(n1403) );
  AOI22_X1 U1333 ( .A1(n2081), .A2(\REGISTERS[24][5] ), .B1(n2078), .B2(
        \REGISTERS[31][5] ), .ZN(n1404) );
  AOI22_X1 U1334 ( .A1(n2104), .A2(\REGISTERS[8][6] ), .B1(n2101), .B2(
        \REGISTERS[13][6] ), .ZN(n1420) );
  AOI22_X1 U1335 ( .A1(n2092), .A2(\REGISTERS[0][6] ), .B1(n2089), .B2(
        \REGISTERS[5][6] ), .ZN(n1421) );
  AOI22_X1 U1336 ( .A1(n2080), .A2(\REGISTERS[24][6] ), .B1(n2077), .B2(
        \REGISTERS[31][6] ), .ZN(n1422) );
  AOI22_X1 U1337 ( .A1(n2104), .A2(\REGISTERS[8][7] ), .B1(n2101), .B2(
        \REGISTERS[13][7] ), .ZN(n1438) );
  AOI22_X1 U1338 ( .A1(n2092), .A2(\REGISTERS[0][7] ), .B1(n2089), .B2(
        \REGISTERS[5][7] ), .ZN(n1439) );
  AOI22_X1 U1339 ( .A1(n2080), .A2(\REGISTERS[24][7] ), .B1(n2077), .B2(
        \REGISTERS[31][7] ), .ZN(n1440) );
  AOI22_X1 U1340 ( .A1(n2104), .A2(\REGISTERS[8][8] ), .B1(n2101), .B2(
        \REGISTERS[13][8] ), .ZN(n1456) );
  AOI22_X1 U1341 ( .A1(n2092), .A2(\REGISTERS[0][8] ), .B1(n2089), .B2(
        \REGISTERS[5][8] ), .ZN(n1457) );
  AOI22_X1 U1342 ( .A1(n2080), .A2(\REGISTERS[24][8] ), .B1(n2077), .B2(
        \REGISTERS[31][8] ), .ZN(n1458) );
  AOI22_X1 U1343 ( .A1(n2104), .A2(\REGISTERS[8][9] ), .B1(n2101), .B2(
        \REGISTERS[13][9] ), .ZN(n1474) );
  AOI22_X1 U1344 ( .A1(n2092), .A2(\REGISTERS[0][9] ), .B1(n2089), .B2(
        \REGISTERS[5][9] ), .ZN(n1475) );
  AOI22_X1 U1345 ( .A1(n2080), .A2(\REGISTERS[24][9] ), .B1(n2077), .B2(
        \REGISTERS[31][9] ), .ZN(n1476) );
  AOI22_X1 U1346 ( .A1(n2104), .A2(\REGISTERS[8][10] ), .B1(n2101), .B2(
        \REGISTERS[13][10] ), .ZN(n1492) );
  AOI22_X1 U1347 ( .A1(n2092), .A2(\REGISTERS[0][10] ), .B1(n2089), .B2(
        \REGISTERS[5][10] ), .ZN(n1493) );
  AOI22_X1 U1348 ( .A1(n2080), .A2(\REGISTERS[24][10] ), .B1(n2077), .B2(
        \REGISTERS[31][10] ), .ZN(n1494) );
  AOI22_X1 U1349 ( .A1(n2104), .A2(\REGISTERS[8][11] ), .B1(n2101), .B2(
        \REGISTERS[13][11] ), .ZN(n1510) );
  AOI22_X1 U1350 ( .A1(n2092), .A2(\REGISTERS[0][11] ), .B1(n2089), .B2(
        \REGISTERS[5][11] ), .ZN(n1511) );
  AOI22_X1 U1351 ( .A1(n2080), .A2(\REGISTERS[24][11] ), .B1(n2077), .B2(
        \REGISTERS[31][11] ), .ZN(n1512) );
  AOI22_X1 U1352 ( .A1(n2104), .A2(\REGISTERS[8][12] ), .B1(n2101), .B2(
        \REGISTERS[13][12] ), .ZN(n1528) );
  AOI22_X1 U1353 ( .A1(n2092), .A2(\REGISTERS[0][12] ), .B1(n2089), .B2(
        \REGISTERS[5][12] ), .ZN(n1529) );
  AOI22_X1 U1354 ( .A1(n2080), .A2(\REGISTERS[24][12] ), .B1(n2077), .B2(
        \REGISTERS[31][12] ), .ZN(n1530) );
  AOI22_X1 U1355 ( .A1(n2104), .A2(\REGISTERS[8][13] ), .B1(n2101), .B2(
        \REGISTERS[13][13] ), .ZN(n1546) );
  AOI22_X1 U1356 ( .A1(n2092), .A2(\REGISTERS[0][13] ), .B1(n2089), .B2(
        \REGISTERS[5][13] ), .ZN(n1547) );
  AOI22_X1 U1357 ( .A1(n2080), .A2(\REGISTERS[24][13] ), .B1(n2077), .B2(
        \REGISTERS[31][13] ), .ZN(n1548) );
  AOI22_X1 U1358 ( .A1(n2104), .A2(\REGISTERS[8][14] ), .B1(n2101), .B2(
        \REGISTERS[13][14] ), .ZN(n1564) );
  AOI22_X1 U1359 ( .A1(n2092), .A2(\REGISTERS[0][14] ), .B1(n2089), .B2(
        \REGISTERS[5][14] ), .ZN(n1565) );
  AOI22_X1 U1360 ( .A1(n2080), .A2(\REGISTERS[24][14] ), .B1(n2077), .B2(
        \REGISTERS[31][14] ), .ZN(n1566) );
  AOI22_X1 U1361 ( .A1(n2104), .A2(\REGISTERS[8][15] ), .B1(n2101), .B2(
        \REGISTERS[13][15] ), .ZN(n1582) );
  AOI22_X1 U1362 ( .A1(n2092), .A2(\REGISTERS[0][15] ), .B1(n2089), .B2(
        \REGISTERS[5][15] ), .ZN(n1583) );
  AOI22_X1 U1363 ( .A1(n2080), .A2(\REGISTERS[24][15] ), .B1(n2077), .B2(
        \REGISTERS[31][15] ), .ZN(n1584) );
  AOI22_X1 U1364 ( .A1(n2104), .A2(\REGISTERS[8][16] ), .B1(n2101), .B2(
        \REGISTERS[13][16] ), .ZN(n1600) );
  AOI22_X1 U1365 ( .A1(n2092), .A2(\REGISTERS[0][16] ), .B1(n2089), .B2(
        \REGISTERS[5][16] ), .ZN(n1601) );
  AOI22_X1 U1366 ( .A1(n2080), .A2(\REGISTERS[24][16] ), .B1(n2077), .B2(
        \REGISTERS[31][16] ), .ZN(n1602) );
  AOI22_X1 U1367 ( .A1(n2104), .A2(\REGISTERS[8][17] ), .B1(n2101), .B2(
        \REGISTERS[13][17] ), .ZN(n1618) );
  AOI22_X1 U1368 ( .A1(n2092), .A2(\REGISTERS[0][17] ), .B1(n2089), .B2(
        \REGISTERS[5][17] ), .ZN(n1619) );
  AOI22_X1 U1369 ( .A1(n2080), .A2(\REGISTERS[24][17] ), .B1(n2077), .B2(
        \REGISTERS[31][17] ), .ZN(n1620) );
  AOI22_X1 U1370 ( .A1(n2104), .A2(\REGISTERS[8][18] ), .B1(n2101), .B2(
        \REGISTERS[13][18] ), .ZN(n1636) );
  AOI22_X1 U1371 ( .A1(n2092), .A2(\REGISTERS[0][18] ), .B1(n2089), .B2(
        \REGISTERS[5][18] ), .ZN(n1637) );
  AOI22_X1 U1372 ( .A1(n2080), .A2(\REGISTERS[24][18] ), .B1(n2077), .B2(
        \REGISTERS[31][18] ), .ZN(n1638) );
  AOI22_X1 U1373 ( .A1(n2103), .A2(\REGISTERS[8][19] ), .B1(n2100), .B2(
        \REGISTERS[13][19] ), .ZN(n1654) );
  AOI22_X1 U1374 ( .A1(n2091), .A2(\REGISTERS[0][19] ), .B1(n2088), .B2(
        \REGISTERS[5][19] ), .ZN(n1655) );
  AOI22_X1 U1375 ( .A1(n2079), .A2(\REGISTERS[24][19] ), .B1(n2076), .B2(
        \REGISTERS[31][19] ), .ZN(n1656) );
  AOI22_X1 U1376 ( .A1(n2103), .A2(\REGISTERS[8][20] ), .B1(n2100), .B2(
        \REGISTERS[13][20] ), .ZN(n1672) );
  AOI22_X1 U1377 ( .A1(n2091), .A2(\REGISTERS[0][20] ), .B1(n2088), .B2(
        \REGISTERS[5][20] ), .ZN(n1673) );
  AOI22_X1 U1378 ( .A1(n2079), .A2(\REGISTERS[24][20] ), .B1(n2076), .B2(
        \REGISTERS[31][20] ), .ZN(n1674) );
  AOI22_X1 U1379 ( .A1(n2103), .A2(\REGISTERS[8][21] ), .B1(n2100), .B2(
        \REGISTERS[13][21] ), .ZN(n1690) );
  AOI22_X1 U1380 ( .A1(n2091), .A2(\REGISTERS[0][21] ), .B1(n2088), .B2(
        \REGISTERS[5][21] ), .ZN(n1691) );
  AOI22_X1 U1381 ( .A1(n2079), .A2(\REGISTERS[24][21] ), .B1(n2076), .B2(
        \REGISTERS[31][21] ), .ZN(n1692) );
  AOI22_X1 U1382 ( .A1(n2103), .A2(\REGISTERS[8][22] ), .B1(n2100), .B2(
        \REGISTERS[13][22] ), .ZN(n1708) );
  AOI22_X1 U1383 ( .A1(n2091), .A2(\REGISTERS[0][22] ), .B1(n2088), .B2(
        \REGISTERS[5][22] ), .ZN(n1709) );
  AOI22_X1 U1384 ( .A1(n2079), .A2(\REGISTERS[24][22] ), .B1(n2076), .B2(
        \REGISTERS[31][22] ), .ZN(n1710) );
  AOI22_X1 U1385 ( .A1(n2103), .A2(\REGISTERS[8][23] ), .B1(n2100), .B2(
        \REGISTERS[13][23] ), .ZN(n1726) );
  AOI22_X1 U1386 ( .A1(n2091), .A2(\REGISTERS[0][23] ), .B1(n2088), .B2(
        \REGISTERS[5][23] ), .ZN(n1727) );
  AOI22_X1 U1387 ( .A1(n2079), .A2(\REGISTERS[24][23] ), .B1(n2076), .B2(
        \REGISTERS[31][23] ), .ZN(n1728) );
  AOI22_X1 U1388 ( .A1(n2103), .A2(\REGISTERS[8][24] ), .B1(n2100), .B2(
        \REGISTERS[13][24] ), .ZN(n1744) );
  AOI22_X1 U1389 ( .A1(n2091), .A2(\REGISTERS[0][24] ), .B1(n2088), .B2(
        \REGISTERS[5][24] ), .ZN(n1745) );
  AOI22_X1 U1390 ( .A1(n2079), .A2(\REGISTERS[24][24] ), .B1(n2076), .B2(
        \REGISTERS[31][24] ), .ZN(n1746) );
  AOI22_X1 U1391 ( .A1(n2103), .A2(\REGISTERS[8][25] ), .B1(n2100), .B2(
        \REGISTERS[13][25] ), .ZN(n1762) );
  AOI22_X1 U1392 ( .A1(n2091), .A2(\REGISTERS[0][25] ), .B1(n2088), .B2(
        \REGISTERS[5][25] ), .ZN(n1763) );
  AOI22_X1 U1393 ( .A1(n2079), .A2(\REGISTERS[24][25] ), .B1(n2076), .B2(
        \REGISTERS[31][25] ), .ZN(n1764) );
  AOI22_X1 U1394 ( .A1(n2103), .A2(\REGISTERS[8][26] ), .B1(n2100), .B2(
        \REGISTERS[13][26] ), .ZN(n1780) );
  AOI22_X1 U1395 ( .A1(n2091), .A2(\REGISTERS[0][26] ), .B1(n2088), .B2(
        \REGISTERS[5][26] ), .ZN(n1781) );
  AOI22_X1 U1396 ( .A1(n2079), .A2(\REGISTERS[24][26] ), .B1(n2076), .B2(
        \REGISTERS[31][26] ), .ZN(n1782) );
  AOI22_X1 U1397 ( .A1(n2103), .A2(\REGISTERS[8][27] ), .B1(n2100), .B2(
        \REGISTERS[13][27] ), .ZN(n1798) );
  AOI22_X1 U1398 ( .A1(n2091), .A2(\REGISTERS[0][27] ), .B1(n2088), .B2(
        \REGISTERS[5][27] ), .ZN(n1799) );
  AOI22_X1 U1399 ( .A1(n2079), .A2(\REGISTERS[24][27] ), .B1(n2076), .B2(
        \REGISTERS[31][27] ), .ZN(n1800) );
  AOI22_X1 U1400 ( .A1(n2103), .A2(\REGISTERS[8][28] ), .B1(n2100), .B2(
        \REGISTERS[13][28] ), .ZN(n1816) );
  AOI22_X1 U1401 ( .A1(n2091), .A2(\REGISTERS[0][28] ), .B1(n2088), .B2(
        \REGISTERS[5][28] ), .ZN(n1817) );
  AOI22_X1 U1402 ( .A1(n2079), .A2(\REGISTERS[24][28] ), .B1(n2076), .B2(
        \REGISTERS[31][28] ), .ZN(n1818) );
  AOI22_X1 U1403 ( .A1(n2103), .A2(\REGISTERS[8][29] ), .B1(n2100), .B2(
        \REGISTERS[13][29] ), .ZN(n1834) );
  AOI22_X1 U1404 ( .A1(n2091), .A2(\REGISTERS[0][29] ), .B1(n2088), .B2(
        \REGISTERS[5][29] ), .ZN(n1835) );
  AOI22_X1 U1405 ( .A1(n2079), .A2(\REGISTERS[24][29] ), .B1(n2076), .B2(
        \REGISTERS[31][29] ), .ZN(n1836) );
  AOI22_X1 U1406 ( .A1(n2103), .A2(\REGISTERS[8][30] ), .B1(n2100), .B2(
        \REGISTERS[13][30] ), .ZN(n1852) );
  AOI22_X1 U1407 ( .A1(n2091), .A2(\REGISTERS[0][30] ), .B1(n2088), .B2(
        \REGISTERS[5][30] ), .ZN(n1853) );
  AOI22_X1 U1408 ( .A1(n2079), .A2(\REGISTERS[24][30] ), .B1(n2076), .B2(
        \REGISTERS[31][30] ), .ZN(n1854) );
  AOI22_X1 U1409 ( .A1(n2103), .A2(\REGISTERS[8][31] ), .B1(n2100), .B2(
        \REGISTERS[13][31] ), .ZN(n1870) );
  AOI22_X1 U1410 ( .A1(n2091), .A2(\REGISTERS[0][31] ), .B1(n2088), .B2(
        \REGISTERS[5][31] ), .ZN(n1878) );
  AOI22_X1 U1411 ( .A1(n2079), .A2(\REGISTERS[24][31] ), .B1(n2076), .B2(
        \REGISTERS[31][31] ), .ZN(n1881) );
  NOR2_X1 U1412 ( .A1(n1256), .A2(ADDR_RD2[1]), .ZN(n1246) );
  NOR2_X1 U1413 ( .A1(n1893), .A2(ADDR_RD1[1]), .ZN(n1887) );
  NAND4_X1 U1414 ( .A1(n73), .A2(n74), .A3(n75), .A4(n76), .ZN(n1981) );
  AOI221_X1 U1415 ( .B1(\REGISTERS[15][1] ), .B2(n2125), .C1(DATA_OUT_2[1]), 
        .C2(n2118), .A(n108), .ZN(n73) );
  AOI221_X1 U1416 ( .B1(\REGISTERS[7][1] ), .B2(n2137), .C1(\REGISTERS[10][1] ), .C2(n2134), .A(n105), .ZN(n74) );
  NOR4_X1 U1417 ( .A1(n93), .A2(n94), .A3(n95), .A4(n96), .ZN(n75) );
  NAND4_X1 U1418 ( .A1(n111), .A2(n112), .A3(n113), .A4(n114), .ZN(n1982) );
  AOI221_X1 U1419 ( .B1(\REGISTERS[15][2] ), .B2(n2125), .C1(DATA_OUT_2[2]), 
        .C2(n2119), .A(n146), .ZN(n111) );
  AOI221_X1 U1420 ( .B1(\REGISTERS[7][2] ), .B2(n2137), .C1(\REGISTERS[10][2] ), .C2(n2134), .A(n143), .ZN(n112) );
  NOR4_X1 U1421 ( .A1(n131), .A2(n132), .A3(n133), .A4(n134), .ZN(n113) );
  NAND4_X1 U1422 ( .A1(n149), .A2(n150), .A3(n151), .A4(n152), .ZN(n1983) );
  AOI221_X1 U1423 ( .B1(\REGISTERS[15][3] ), .B2(n2125), .C1(DATA_OUT_2[3]), 
        .C2(n2119), .A(n184), .ZN(n149) );
  AOI221_X1 U1424 ( .B1(\REGISTERS[7][3] ), .B2(n2137), .C1(\REGISTERS[10][3] ), .C2(n2134), .A(n181), .ZN(n150) );
  NOR4_X1 U1425 ( .A1(n169), .A2(n170), .A3(n171), .A4(n172), .ZN(n151) );
  NAND4_X1 U1426 ( .A1(n187), .A2(n188), .A3(n189), .A4(n190), .ZN(n1984) );
  AOI221_X1 U1427 ( .B1(\REGISTERS[15][4] ), .B2(n2125), .C1(DATA_OUT_2[4]), 
        .C2(n2118), .A(n222), .ZN(n187) );
  AOI221_X1 U1428 ( .B1(\REGISTERS[7][4] ), .B2(n2137), .C1(\REGISTERS[10][4] ), .C2(n2134), .A(n219), .ZN(n188) );
  NOR4_X1 U1429 ( .A1(n207), .A2(n208), .A3(n209), .A4(n210), .ZN(n189) );
  NAND4_X1 U1430 ( .A1(n225), .A2(n226), .A3(n227), .A4(n228), .ZN(n1985) );
  AOI221_X1 U1431 ( .B1(\REGISTERS[15][5] ), .B2(n2125), .C1(DATA_OUT_2[5]), 
        .C2(n2118), .A(n260), .ZN(n225) );
  AOI221_X1 U1432 ( .B1(\REGISTERS[7][5] ), .B2(n2137), .C1(\REGISTERS[10][5] ), .C2(n2134), .A(n257), .ZN(n226) );
  NOR4_X1 U1433 ( .A1(n245), .A2(n246), .A3(n247), .A4(n248), .ZN(n227) );
  NAND4_X1 U1434 ( .A1(n263), .A2(n264), .A3(n265), .A4(n266), .ZN(n1986) );
  AOI221_X1 U1435 ( .B1(\REGISTERS[15][6] ), .B2(n2124), .C1(DATA_OUT_2[6]), 
        .C2(n2119), .A(n298), .ZN(n263) );
  AOI221_X1 U1436 ( .B1(\REGISTERS[7][6] ), .B2(n2136), .C1(\REGISTERS[10][6] ), .C2(n2133), .A(n295), .ZN(n264) );
  NOR4_X1 U1437 ( .A1(n283), .A2(n284), .A3(n285), .A4(n286), .ZN(n265) );
  NAND4_X1 U1438 ( .A1(n301), .A2(n302), .A3(n303), .A4(n304), .ZN(n1987) );
  AOI221_X1 U1439 ( .B1(\REGISTERS[15][7] ), .B2(n2124), .C1(DATA_OUT_2[7]), 
        .C2(n2119), .A(n336), .ZN(n301) );
  AOI221_X1 U1440 ( .B1(\REGISTERS[7][7] ), .B2(n2136), .C1(\REGISTERS[10][7] ), .C2(n2133), .A(n333), .ZN(n302) );
  NOR4_X1 U1441 ( .A1(n321), .A2(n322), .A3(n323), .A4(n324), .ZN(n303) );
  NAND4_X1 U1442 ( .A1(n339), .A2(n340), .A3(n341), .A4(n342), .ZN(n1988) );
  AOI221_X1 U1443 ( .B1(\REGISTERS[15][8] ), .B2(n2124), .C1(DATA_OUT_2[8]), 
        .C2(n2119), .A(n374), .ZN(n339) );
  AOI221_X1 U1444 ( .B1(\REGISTERS[7][8] ), .B2(n2136), .C1(\REGISTERS[10][8] ), .C2(n2133), .A(n371), .ZN(n340) );
  NOR4_X1 U1445 ( .A1(n359), .A2(n360), .A3(n361), .A4(n362), .ZN(n341) );
  NAND4_X1 U1446 ( .A1(n377), .A2(n378), .A3(n379), .A4(n380), .ZN(n1989) );
  AOI221_X1 U1447 ( .B1(\REGISTERS[15][9] ), .B2(n2124), .C1(DATA_OUT_2[9]), 
        .C2(n2119), .A(n412), .ZN(n377) );
  AOI221_X1 U1448 ( .B1(\REGISTERS[7][9] ), .B2(n2136), .C1(\REGISTERS[10][9] ), .C2(n2133), .A(n409), .ZN(n378) );
  NOR4_X1 U1449 ( .A1(n397), .A2(n398), .A3(n399), .A4(n400), .ZN(n379) );
  NAND4_X1 U1450 ( .A1(n415), .A2(n416), .A3(n417), .A4(n418), .ZN(n1990) );
  AOI221_X1 U1451 ( .B1(\REGISTERS[15][10] ), .B2(n2124), .C1(DATA_OUT_2[10]), 
        .C2(n2119), .A(n450), .ZN(n415) );
  AOI221_X1 U1452 ( .B1(\REGISTERS[7][10] ), .B2(n2136), .C1(
        \REGISTERS[10][10] ), .C2(n2133), .A(n447), .ZN(n416) );
  NOR4_X1 U1453 ( .A1(n435), .A2(n436), .A3(n437), .A4(n438), .ZN(n417) );
  NAND4_X1 U1454 ( .A1(n453), .A2(n454), .A3(n455), .A4(n456), .ZN(n1991) );
  AOI221_X1 U1455 ( .B1(\REGISTERS[15][11] ), .B2(n2124), .C1(DATA_OUT_2[11]), 
        .C2(n2119), .A(n488), .ZN(n453) );
  AOI221_X1 U1456 ( .B1(\REGISTERS[7][11] ), .B2(n2136), .C1(
        \REGISTERS[10][11] ), .C2(n2133), .A(n485), .ZN(n454) );
  NOR4_X1 U1457 ( .A1(n473), .A2(n474), .A3(n475), .A4(n476), .ZN(n455) );
  NAND4_X1 U1458 ( .A1(n491), .A2(n492), .A3(n493), .A4(n494), .ZN(n1992) );
  AOI221_X1 U1459 ( .B1(\REGISTERS[15][12] ), .B2(n2124), .C1(DATA_OUT_2[12]), 
        .C2(n2119), .A(n526), .ZN(n491) );
  AOI221_X1 U1460 ( .B1(\REGISTERS[7][12] ), .B2(n2136), .C1(
        \REGISTERS[10][12] ), .C2(n2133), .A(n523), .ZN(n492) );
  NOR4_X1 U1461 ( .A1(n511), .A2(n512), .A3(n513), .A4(n514), .ZN(n493) );
  NAND4_X1 U1462 ( .A1(n529), .A2(n530), .A3(n531), .A4(n532), .ZN(n1993) );
  AOI221_X1 U1463 ( .B1(\REGISTERS[15][13] ), .B2(n2124), .C1(DATA_OUT_2[13]), 
        .C2(n2119), .A(n564), .ZN(n529) );
  AOI221_X1 U1464 ( .B1(\REGISTERS[7][13] ), .B2(n2136), .C1(
        \REGISTERS[10][13] ), .C2(n2133), .A(n561), .ZN(n530) );
  NOR4_X1 U1465 ( .A1(n549), .A2(n550), .A3(n551), .A4(n552), .ZN(n531) );
  NAND4_X1 U1466 ( .A1(n567), .A2(n568), .A3(n569), .A4(n570), .ZN(n1994) );
  AOI221_X1 U1467 ( .B1(\REGISTERS[15][14] ), .B2(n2124), .C1(DATA_OUT_2[14]), 
        .C2(n2119), .A(n602), .ZN(n567) );
  AOI221_X1 U1468 ( .B1(\REGISTERS[7][14] ), .B2(n2136), .C1(
        \REGISTERS[10][14] ), .C2(n2133), .A(n599), .ZN(n568) );
  NOR4_X1 U1469 ( .A1(n587), .A2(n588), .A3(n589), .A4(n590), .ZN(n569) );
  NAND4_X1 U1470 ( .A1(n605), .A2(n606), .A3(n607), .A4(n608), .ZN(n1995) );
  AOI221_X1 U1471 ( .B1(\REGISTERS[15][15] ), .B2(n2124), .C1(DATA_OUT_2[15]), 
        .C2(n2119), .A(n640), .ZN(n605) );
  AOI221_X1 U1472 ( .B1(\REGISTERS[7][15] ), .B2(n2136), .C1(
        \REGISTERS[10][15] ), .C2(n2133), .A(n637), .ZN(n606) );
  NOR4_X1 U1473 ( .A1(n625), .A2(n626), .A3(n627), .A4(n628), .ZN(n607) );
  NAND4_X1 U1474 ( .A1(n643), .A2(n644), .A3(n645), .A4(n646), .ZN(n1996) );
  AOI221_X1 U1475 ( .B1(\REGISTERS[15][16] ), .B2(n2124), .C1(DATA_OUT_2[16]), 
        .C2(n2119), .A(n678), .ZN(n643) );
  AOI221_X1 U1476 ( .B1(\REGISTERS[7][16] ), .B2(n2136), .C1(
        \REGISTERS[10][16] ), .C2(n2133), .A(n675), .ZN(n644) );
  NOR4_X1 U1477 ( .A1(n663), .A2(n664), .A3(n665), .A4(n666), .ZN(n645) );
  NAND4_X1 U1478 ( .A1(n681), .A2(n682), .A3(n683), .A4(n684), .ZN(n1997) );
  AOI221_X1 U1479 ( .B1(\REGISTERS[15][17] ), .B2(n2124), .C1(DATA_OUT_2[17]), 
        .C2(n2119), .A(n716), .ZN(n681) );
  AOI221_X1 U1480 ( .B1(\REGISTERS[7][17] ), .B2(n2136), .C1(
        \REGISTERS[10][17] ), .C2(n2133), .A(n713), .ZN(n682) );
  NOR4_X1 U1481 ( .A1(n701), .A2(n702), .A3(n703), .A4(n704), .ZN(n683) );
  NAND4_X1 U1482 ( .A1(n719), .A2(n720), .A3(n721), .A4(n722), .ZN(n1998) );
  AOI221_X1 U1483 ( .B1(\REGISTERS[15][18] ), .B2(n2124), .C1(DATA_OUT_2[18]), 
        .C2(n2119), .A(n754), .ZN(n719) );
  AOI221_X1 U1484 ( .B1(\REGISTERS[7][18] ), .B2(n2136), .C1(
        \REGISTERS[10][18] ), .C2(n2133), .A(n751), .ZN(n720) );
  NOR4_X1 U1485 ( .A1(n739), .A2(n740), .A3(n741), .A4(n742), .ZN(n721) );
  NAND4_X1 U1486 ( .A1(n757), .A2(n758), .A3(n759), .A4(n760), .ZN(n1999) );
  AOI221_X1 U1487 ( .B1(\REGISTERS[15][19] ), .B2(n2123), .C1(DATA_OUT_2[19]), 
        .C2(n2118), .A(n792), .ZN(n757) );
  AOI221_X1 U1488 ( .B1(\REGISTERS[7][19] ), .B2(n2135), .C1(
        \REGISTERS[10][19] ), .C2(n2132), .A(n789), .ZN(n758) );
  NOR4_X1 U1489 ( .A1(n777), .A2(n778), .A3(n779), .A4(n780), .ZN(n759) );
  NAND4_X1 U1490 ( .A1(n795), .A2(n796), .A3(n797), .A4(n798), .ZN(n2000) );
  AOI221_X1 U1491 ( .B1(\REGISTERS[15][20] ), .B2(n2123), .C1(DATA_OUT_2[20]), 
        .C2(n2118), .A(n830), .ZN(n795) );
  AOI221_X1 U1492 ( .B1(\REGISTERS[7][20] ), .B2(n2135), .C1(
        \REGISTERS[10][20] ), .C2(n2132), .A(n827), .ZN(n796) );
  NOR4_X1 U1493 ( .A1(n815), .A2(n816), .A3(n817), .A4(n818), .ZN(n797) );
  NAND4_X1 U1494 ( .A1(n833), .A2(n834), .A3(n835), .A4(n836), .ZN(n2001) );
  AOI221_X1 U1495 ( .B1(\REGISTERS[15][21] ), .B2(n2123), .C1(DATA_OUT_2[21]), 
        .C2(n2118), .A(n868), .ZN(n833) );
  AOI221_X1 U1496 ( .B1(\REGISTERS[7][21] ), .B2(n2135), .C1(
        \REGISTERS[10][21] ), .C2(n2132), .A(n865), .ZN(n834) );
  NOR4_X1 U1497 ( .A1(n853), .A2(n854), .A3(n855), .A4(n856), .ZN(n835) );
  NAND4_X1 U1498 ( .A1(n871), .A2(n872), .A3(n873), .A4(n874), .ZN(n2002) );
  AOI221_X1 U1499 ( .B1(\REGISTERS[15][22] ), .B2(n2123), .C1(DATA_OUT_2[22]), 
        .C2(n2118), .A(n906), .ZN(n871) );
  AOI221_X1 U1500 ( .B1(\REGISTERS[7][22] ), .B2(n2135), .C1(
        \REGISTERS[10][22] ), .C2(n2132), .A(n903), .ZN(n872) );
  NOR4_X1 U1501 ( .A1(n891), .A2(n892), .A3(n893), .A4(n894), .ZN(n873) );
  NAND4_X1 U1502 ( .A1(n909), .A2(n910), .A3(n911), .A4(n912), .ZN(n2003) );
  AOI221_X1 U1503 ( .B1(\REGISTERS[15][23] ), .B2(n2123), .C1(DATA_OUT_2[23]), 
        .C2(n2118), .A(n944), .ZN(n909) );
  AOI221_X1 U1504 ( .B1(\REGISTERS[7][23] ), .B2(n2135), .C1(
        \REGISTERS[10][23] ), .C2(n2132), .A(n941), .ZN(n910) );
  NOR4_X1 U1505 ( .A1(n929), .A2(n930), .A3(n931), .A4(n932), .ZN(n911) );
  NAND4_X1 U1506 ( .A1(n947), .A2(n948), .A3(n949), .A4(n950), .ZN(n2004) );
  AOI221_X1 U1507 ( .B1(\REGISTERS[15][24] ), .B2(n2123), .C1(DATA_OUT_2[24]), 
        .C2(n2118), .A(n982), .ZN(n947) );
  AOI221_X1 U1508 ( .B1(\REGISTERS[7][24] ), .B2(n2135), .C1(
        \REGISTERS[10][24] ), .C2(n2132), .A(n979), .ZN(n948) );
  NOR4_X1 U1509 ( .A1(n967), .A2(n968), .A3(n969), .A4(n970), .ZN(n949) );
  NAND4_X1 U1510 ( .A1(n985), .A2(n986), .A3(n987), .A4(n988), .ZN(n2005) );
  AOI221_X1 U1511 ( .B1(\REGISTERS[15][25] ), .B2(n2123), .C1(DATA_OUT_2[25]), 
        .C2(n2118), .A(n1020), .ZN(n985) );
  AOI221_X1 U1512 ( .B1(\REGISTERS[7][25] ), .B2(n2135), .C1(
        \REGISTERS[10][25] ), .C2(n2132), .A(n1017), .ZN(n986) );
  NOR4_X1 U1513 ( .A1(n1005), .A2(n1006), .A3(n1007), .A4(n1008), .ZN(n987) );
  NAND4_X1 U1514 ( .A1(n1023), .A2(n1024), .A3(n1025), .A4(n1026), .ZN(n2006)
         );
  AOI221_X1 U1515 ( .B1(\REGISTERS[15][26] ), .B2(n2123), .C1(DATA_OUT_2[26]), 
        .C2(n2118), .A(n1058), .ZN(n1023) );
  AOI221_X1 U1516 ( .B1(\REGISTERS[7][26] ), .B2(n2135), .C1(
        \REGISTERS[10][26] ), .C2(n2132), .A(n1055), .ZN(n1024) );
  NOR4_X1 U1517 ( .A1(n1043), .A2(n1044), .A3(n1045), .A4(n1046), .ZN(n1025)
         );
  NAND4_X1 U1518 ( .A1(n1061), .A2(n1062), .A3(n1063), .A4(n1064), .ZN(n2007)
         );
  AOI221_X1 U1519 ( .B1(\REGISTERS[15][27] ), .B2(n2123), .C1(DATA_OUT_2[27]), 
        .C2(n2118), .A(n1096), .ZN(n1061) );
  AOI221_X1 U1520 ( .B1(\REGISTERS[7][27] ), .B2(n2135), .C1(
        \REGISTERS[10][27] ), .C2(n2132), .A(n1093), .ZN(n1062) );
  NOR4_X1 U1521 ( .A1(n1081), .A2(n1082), .A3(n1083), .A4(n1084), .ZN(n1063)
         );
  NAND4_X1 U1522 ( .A1(n1099), .A2(n1100), .A3(n1101), .A4(n1102), .ZN(n2008)
         );
  AOI221_X1 U1523 ( .B1(\REGISTERS[15][28] ), .B2(n2123), .C1(DATA_OUT_2[28]), 
        .C2(n2118), .A(n1134), .ZN(n1099) );
  AOI221_X1 U1524 ( .B1(\REGISTERS[7][28] ), .B2(n2135), .C1(
        \REGISTERS[10][28] ), .C2(n2132), .A(n1131), .ZN(n1100) );
  NOR4_X1 U1525 ( .A1(n1119), .A2(n1120), .A3(n1121), .A4(n1122), .ZN(n1101)
         );
  NAND4_X1 U1526 ( .A1(n1137), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n2009)
         );
  AOI221_X1 U1527 ( .B1(\REGISTERS[15][29] ), .B2(n2123), .C1(DATA_OUT_2[29]), 
        .C2(n2118), .A(n1172), .ZN(n1137) );
  AOI221_X1 U1528 ( .B1(\REGISTERS[7][29] ), .B2(n2135), .C1(
        \REGISTERS[10][29] ), .C2(n2132), .A(n1169), .ZN(n1138) );
  NOR4_X1 U1529 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1139)
         );
  NAND4_X1 U1530 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n2010)
         );
  AOI221_X1 U1531 ( .B1(\REGISTERS[15][30] ), .B2(n2123), .C1(DATA_OUT_2[30]), 
        .C2(n2118), .A(n1210), .ZN(n1175) );
  AOI221_X1 U1532 ( .B1(\REGISTERS[7][30] ), .B2(n2135), .C1(
        \REGISTERS[10][30] ), .C2(n2132), .A(n1207), .ZN(n1176) );
  NOR4_X1 U1533 ( .A1(n1195), .A2(n1196), .A3(n1197), .A4(n1198), .ZN(n1177)
         );
  NAND4_X1 U1534 ( .A1(n1213), .A2(n1214), .A3(n1215), .A4(n1216), .ZN(n2011)
         );
  AOI221_X1 U1535 ( .B1(\REGISTERS[15][31] ), .B2(n2123), .C1(DATA_OUT_2[31]), 
        .C2(n2119), .A(n1266), .ZN(n1213) );
  AOI221_X1 U1536 ( .B1(\REGISTERS[7][31] ), .B2(n2135), .C1(
        \REGISTERS[10][31] ), .C2(n2132), .A(n1263), .ZN(n1214) );
  NOR4_X1 U1537 ( .A1(n1248), .A2(n1249), .A3(n1250), .A4(n1251), .ZN(n1215)
         );
  NAND4_X1 U1538 ( .A1(n1271), .A2(n1272), .A3(n1273), .A4(n1274), .ZN(n2012)
         );
  AOI221_X1 U1539 ( .B1(n1962), .B2(\REGISTERS[15][0] ), .C1(DATA_OUT_1[0]), 
        .C2(n1955), .A(n1319), .ZN(n1271) );
  AOI221_X1 U1540 ( .B1(n1974), .B2(\REGISTERS[7][0] ), .C1(n1971), .C2(
        \REGISTERS[10][0] ), .A(n1314), .ZN(n1272) );
  NOR4_X1 U1541 ( .A1(n1300), .A2(n1301), .A3(n1302), .A4(n1303), .ZN(n1273)
         );
  NAND4_X1 U1542 ( .A1(n1322), .A2(n1323), .A3(n1324), .A4(n1325), .ZN(n2013)
         );
  AOI221_X1 U1543 ( .B1(n1962), .B2(\REGISTERS[15][1] ), .C1(DATA_OUT_1[1]), 
        .C2(n1956), .A(n1339), .ZN(n1322) );
  AOI221_X1 U1544 ( .B1(n1974), .B2(\REGISTERS[7][1] ), .C1(n1971), .C2(
        \REGISTERS[10][1] ), .A(n1338), .ZN(n1323) );
  NOR4_X1 U1545 ( .A1(n1334), .A2(n1335), .A3(n1336), .A4(n1337), .ZN(n1324)
         );
  NAND4_X1 U1546 ( .A1(n1340), .A2(n1341), .A3(n1342), .A4(n1343), .ZN(n2014)
         );
  AOI221_X1 U1547 ( .B1(n1962), .B2(\REGISTERS[15][2] ), .C1(DATA_OUT_1[2]), 
        .C2(n1956), .A(n1357), .ZN(n1340) );
  AOI221_X1 U1548 ( .B1(n1974), .B2(\REGISTERS[7][2] ), .C1(n1971), .C2(
        \REGISTERS[10][2] ), .A(n1356), .ZN(n1341) );
  NOR4_X1 U1549 ( .A1(n1352), .A2(n1353), .A3(n1354), .A4(n1355), .ZN(n1342)
         );
  NAND4_X1 U1550 ( .A1(n1358), .A2(n1359), .A3(n1360), .A4(n1361), .ZN(n2015)
         );
  AOI221_X1 U1551 ( .B1(n1962), .B2(\REGISTERS[15][3] ), .C1(DATA_OUT_1[3]), 
        .C2(n1956), .A(n1375), .ZN(n1358) );
  AOI221_X1 U1552 ( .B1(n1974), .B2(\REGISTERS[7][3] ), .C1(n1971), .C2(
        \REGISTERS[10][3] ), .A(n1374), .ZN(n1359) );
  NOR4_X1 U1553 ( .A1(n1370), .A2(n1371), .A3(n1372), .A4(n1373), .ZN(n1360)
         );
  NAND4_X1 U1554 ( .A1(n1376), .A2(n1377), .A3(n1378), .A4(n1379), .ZN(n2016)
         );
  AOI221_X1 U1555 ( .B1(n1962), .B2(\REGISTERS[15][4] ), .C1(DATA_OUT_1[4]), 
        .C2(n1956), .A(n1393), .ZN(n1376) );
  AOI221_X1 U1556 ( .B1(n1974), .B2(\REGISTERS[7][4] ), .C1(n1971), .C2(
        \REGISTERS[10][4] ), .A(n1392), .ZN(n1377) );
  NOR4_X1 U1557 ( .A1(n1388), .A2(n1389), .A3(n1390), .A4(n1391), .ZN(n1378)
         );
  NAND4_X1 U1558 ( .A1(n1394), .A2(n1395), .A3(n1396), .A4(n1397), .ZN(n2017)
         );
  AOI221_X1 U1559 ( .B1(n1962), .B2(\REGISTERS[15][5] ), .C1(DATA_OUT_1[5]), 
        .C2(n1955), .A(n1411), .ZN(n1394) );
  AOI221_X1 U1560 ( .B1(n1974), .B2(\REGISTERS[7][5] ), .C1(n1971), .C2(
        \REGISTERS[10][5] ), .A(n1410), .ZN(n1395) );
  NOR4_X1 U1561 ( .A1(n1406), .A2(n1407), .A3(n1408), .A4(n1409), .ZN(n1396)
         );
  NAND4_X1 U1562 ( .A1(n1412), .A2(n1413), .A3(n1414), .A4(n1415), .ZN(n2018)
         );
  AOI221_X1 U1563 ( .B1(n1961), .B2(\REGISTERS[15][6] ), .C1(DATA_OUT_1[6]), 
        .C2(n1955), .A(n1429), .ZN(n1412) );
  AOI221_X1 U1564 ( .B1(n1973), .B2(\REGISTERS[7][6] ), .C1(n1970), .C2(
        \REGISTERS[10][6] ), .A(n1428), .ZN(n1413) );
  NOR4_X1 U1565 ( .A1(n1424), .A2(n1425), .A3(n1426), .A4(n1427), .ZN(n1414)
         );
  NAND4_X1 U1566 ( .A1(n1430), .A2(n1431), .A3(n1432), .A4(n1433), .ZN(n2019)
         );
  AOI221_X1 U1567 ( .B1(n1961), .B2(\REGISTERS[15][7] ), .C1(DATA_OUT_1[7]), 
        .C2(n1956), .A(n1447), .ZN(n1430) );
  AOI221_X1 U1568 ( .B1(n1973), .B2(\REGISTERS[7][7] ), .C1(n1970), .C2(
        \REGISTERS[10][7] ), .A(n1446), .ZN(n1431) );
  NOR4_X1 U1569 ( .A1(n1442), .A2(n1443), .A3(n1444), .A4(n1445), .ZN(n1432)
         );
  NAND4_X1 U1570 ( .A1(n1448), .A2(n1449), .A3(n1450), .A4(n1451), .ZN(n2020)
         );
  AOI221_X1 U1571 ( .B1(n1961), .B2(\REGISTERS[15][8] ), .C1(DATA_OUT_1[8]), 
        .C2(n1956), .A(n1465), .ZN(n1448) );
  AOI221_X1 U1572 ( .B1(n1973), .B2(\REGISTERS[7][8] ), .C1(n1970), .C2(
        \REGISTERS[10][8] ), .A(n1464), .ZN(n1449) );
  NOR4_X1 U1573 ( .A1(n1460), .A2(n1461), .A3(n1462), .A4(n1463), .ZN(n1450)
         );
  NAND4_X1 U1574 ( .A1(n1466), .A2(n1467), .A3(n1468), .A4(n1469), .ZN(n2021)
         );
  AOI221_X1 U1575 ( .B1(n1961), .B2(\REGISTERS[15][9] ), .C1(DATA_OUT_1[9]), 
        .C2(n1956), .A(n1483), .ZN(n1466) );
  AOI221_X1 U1576 ( .B1(n1973), .B2(\REGISTERS[7][9] ), .C1(n1970), .C2(
        \REGISTERS[10][9] ), .A(n1482), .ZN(n1467) );
  NOR4_X1 U1577 ( .A1(n1478), .A2(n1479), .A3(n1480), .A4(n1481), .ZN(n1468)
         );
  NAND4_X1 U1578 ( .A1(n1484), .A2(n1485), .A3(n1486), .A4(n1487), .ZN(n2022)
         );
  AOI221_X1 U1579 ( .B1(n1961), .B2(\REGISTERS[15][10] ), .C1(DATA_OUT_1[10]), 
        .C2(n1956), .A(n1501), .ZN(n1484) );
  AOI221_X1 U1580 ( .B1(n1973), .B2(\REGISTERS[7][10] ), .C1(n1970), .C2(
        \REGISTERS[10][10] ), .A(n1500), .ZN(n1485) );
  NOR4_X1 U1581 ( .A1(n1496), .A2(n1497), .A3(n1498), .A4(n1499), .ZN(n1486)
         );
  NAND4_X1 U1582 ( .A1(n1502), .A2(n1503), .A3(n1504), .A4(n1505), .ZN(n2023)
         );
  AOI221_X1 U1583 ( .B1(n1961), .B2(\REGISTERS[15][11] ), .C1(DATA_OUT_1[11]), 
        .C2(n1956), .A(n1519), .ZN(n1502) );
  AOI221_X1 U1584 ( .B1(n1973), .B2(\REGISTERS[7][11] ), .C1(n1970), .C2(
        \REGISTERS[10][11] ), .A(n1518), .ZN(n1503) );
  NOR4_X1 U1585 ( .A1(n1514), .A2(n1515), .A3(n1516), .A4(n1517), .ZN(n1504)
         );
  NAND4_X1 U1586 ( .A1(n1520), .A2(n1521), .A3(n1522), .A4(n1523), .ZN(n2024)
         );
  AOI221_X1 U1587 ( .B1(n1961), .B2(\REGISTERS[15][12] ), .C1(DATA_OUT_1[12]), 
        .C2(n1956), .A(n1537), .ZN(n1520) );
  AOI221_X1 U1588 ( .B1(n1973), .B2(\REGISTERS[7][12] ), .C1(n1970), .C2(
        \REGISTERS[10][12] ), .A(n1536), .ZN(n1521) );
  NOR4_X1 U1589 ( .A1(n1532), .A2(n1533), .A3(n1534), .A4(n1535), .ZN(n1522)
         );
  NAND4_X1 U1590 ( .A1(n1538), .A2(n1539), .A3(n1540), .A4(n1541), .ZN(n2025)
         );
  AOI221_X1 U1591 ( .B1(n1961), .B2(\REGISTERS[15][13] ), .C1(DATA_OUT_1[13]), 
        .C2(n1956), .A(n1555), .ZN(n1538) );
  AOI221_X1 U1592 ( .B1(n1973), .B2(\REGISTERS[7][13] ), .C1(n1970), .C2(
        \REGISTERS[10][13] ), .A(n1554), .ZN(n1539) );
  NOR4_X1 U1593 ( .A1(n1550), .A2(n1551), .A3(n1552), .A4(n1553), .ZN(n1540)
         );
  NAND4_X1 U1594 ( .A1(n1556), .A2(n1557), .A3(n1558), .A4(n1559), .ZN(n2026)
         );
  AOI221_X1 U1595 ( .B1(n1961), .B2(\REGISTERS[15][14] ), .C1(DATA_OUT_1[14]), 
        .C2(n1956), .A(n1573), .ZN(n1556) );
  AOI221_X1 U1596 ( .B1(n1973), .B2(\REGISTERS[7][14] ), .C1(n1970), .C2(
        \REGISTERS[10][14] ), .A(n1572), .ZN(n1557) );
  NOR4_X1 U1597 ( .A1(n1568), .A2(n1569), .A3(n1570), .A4(n1571), .ZN(n1558)
         );
  NAND4_X1 U1598 ( .A1(n1574), .A2(n1575), .A3(n1576), .A4(n1577), .ZN(n2027)
         );
  AOI221_X1 U1599 ( .B1(n1961), .B2(\REGISTERS[15][15] ), .C1(DATA_OUT_1[15]), 
        .C2(n1956), .A(n1591), .ZN(n1574) );
  AOI221_X1 U1600 ( .B1(n1973), .B2(\REGISTERS[7][15] ), .C1(n1970), .C2(
        \REGISTERS[10][15] ), .A(n1590), .ZN(n1575) );
  NOR4_X1 U1601 ( .A1(n1586), .A2(n1587), .A3(n1588), .A4(n1589), .ZN(n1576)
         );
  NAND4_X1 U1602 ( .A1(n1592), .A2(n1593), .A3(n1594), .A4(n1595), .ZN(n2028)
         );
  AOI221_X1 U1603 ( .B1(n1961), .B2(\REGISTERS[15][16] ), .C1(DATA_OUT_1[16]), 
        .C2(n1956), .A(n1609), .ZN(n1592) );
  AOI221_X1 U1604 ( .B1(n1973), .B2(\REGISTERS[7][16] ), .C1(n1970), .C2(
        \REGISTERS[10][16] ), .A(n1608), .ZN(n1593) );
  NOR4_X1 U1605 ( .A1(n1604), .A2(n1605), .A3(n1606), .A4(n1607), .ZN(n1594)
         );
  NAND4_X1 U1606 ( .A1(n1610), .A2(n1611), .A3(n1612), .A4(n1613), .ZN(n2029)
         );
  AOI221_X1 U1607 ( .B1(n1961), .B2(\REGISTERS[15][17] ), .C1(DATA_OUT_1[17]), 
        .C2(n1956), .A(n1627), .ZN(n1610) );
  AOI221_X1 U1608 ( .B1(n1973), .B2(\REGISTERS[7][17] ), .C1(n1970), .C2(
        \REGISTERS[10][17] ), .A(n1626), .ZN(n1611) );
  NOR4_X1 U1609 ( .A1(n1622), .A2(n1623), .A3(n1624), .A4(n1625), .ZN(n1612)
         );
  NAND4_X1 U1610 ( .A1(n1628), .A2(n1629), .A3(n1630), .A4(n1631), .ZN(n2030)
         );
  AOI221_X1 U1611 ( .B1(n1961), .B2(\REGISTERS[15][18] ), .C1(DATA_OUT_1[18]), 
        .C2(n1956), .A(n1645), .ZN(n1628) );
  AOI221_X1 U1612 ( .B1(n1973), .B2(\REGISTERS[7][18] ), .C1(n1970), .C2(
        \REGISTERS[10][18] ), .A(n1644), .ZN(n1629) );
  NOR4_X1 U1613 ( .A1(n1640), .A2(n1641), .A3(n1642), .A4(n1643), .ZN(n1630)
         );
  NAND4_X1 U1614 ( .A1(n1646), .A2(n1647), .A3(n1648), .A4(n1649), .ZN(n2031)
         );
  AOI221_X1 U1615 ( .B1(n1960), .B2(\REGISTERS[15][19] ), .C1(DATA_OUT_1[19]), 
        .C2(n1955), .A(n1663), .ZN(n1646) );
  AOI221_X1 U1616 ( .B1(n1972), .B2(\REGISTERS[7][19] ), .C1(n1969), .C2(
        \REGISTERS[10][19] ), .A(n1662), .ZN(n1647) );
  NOR4_X1 U1617 ( .A1(n1658), .A2(n1659), .A3(n1660), .A4(n1661), .ZN(n1648)
         );
  NAND4_X1 U1618 ( .A1(n1664), .A2(n1665), .A3(n1666), .A4(n1667), .ZN(n2032)
         );
  AOI221_X1 U1619 ( .B1(n1960), .B2(\REGISTERS[15][20] ), .C1(DATA_OUT_1[20]), 
        .C2(n1955), .A(n1681), .ZN(n1664) );
  AOI221_X1 U1620 ( .B1(n1972), .B2(\REGISTERS[7][20] ), .C1(n1969), .C2(
        \REGISTERS[10][20] ), .A(n1680), .ZN(n1665) );
  NOR4_X1 U1621 ( .A1(n1676), .A2(n1677), .A3(n1678), .A4(n1679), .ZN(n1666)
         );
  NAND4_X1 U1622 ( .A1(n1682), .A2(n1683), .A3(n1684), .A4(n1685), .ZN(n2033)
         );
  AOI221_X1 U1623 ( .B1(n1960), .B2(\REGISTERS[15][21] ), .C1(DATA_OUT_1[21]), 
        .C2(n1955), .A(n1699), .ZN(n1682) );
  AOI221_X1 U1624 ( .B1(n1972), .B2(\REGISTERS[7][21] ), .C1(n1969), .C2(
        \REGISTERS[10][21] ), .A(n1698), .ZN(n1683) );
  NOR4_X1 U1625 ( .A1(n1694), .A2(n1695), .A3(n1696), .A4(n1697), .ZN(n1684)
         );
  NAND4_X1 U1626 ( .A1(n1700), .A2(n1701), .A3(n1702), .A4(n1703), .ZN(n2034)
         );
  AOI221_X1 U1627 ( .B1(n1960), .B2(\REGISTERS[15][22] ), .C1(DATA_OUT_1[22]), 
        .C2(n1955), .A(n1717), .ZN(n1700) );
  AOI221_X1 U1628 ( .B1(n1972), .B2(\REGISTERS[7][22] ), .C1(n1969), .C2(
        \REGISTERS[10][22] ), .A(n1716), .ZN(n1701) );
  NOR4_X1 U1629 ( .A1(n1712), .A2(n1713), .A3(n1714), .A4(n1715), .ZN(n1702)
         );
  NAND4_X1 U1630 ( .A1(n1718), .A2(n1719), .A3(n1720), .A4(n1721), .ZN(n2035)
         );
  AOI221_X1 U1631 ( .B1(n1960), .B2(\REGISTERS[15][23] ), .C1(DATA_OUT_1[23]), 
        .C2(n1955), .A(n1735), .ZN(n1718) );
  AOI221_X1 U1632 ( .B1(n1972), .B2(\REGISTERS[7][23] ), .C1(n1969), .C2(
        \REGISTERS[10][23] ), .A(n1734), .ZN(n1719) );
  NOR4_X1 U1633 ( .A1(n1730), .A2(n1731), .A3(n1732), .A4(n1733), .ZN(n1720)
         );
  NAND4_X1 U1634 ( .A1(n1736), .A2(n1737), .A3(n1738), .A4(n1739), .ZN(n2036)
         );
  AOI221_X1 U1635 ( .B1(n1960), .B2(\REGISTERS[15][24] ), .C1(DATA_OUT_1[24]), 
        .C2(n1955), .A(n1753), .ZN(n1736) );
  AOI221_X1 U1636 ( .B1(n1972), .B2(\REGISTERS[7][24] ), .C1(n1969), .C2(
        \REGISTERS[10][24] ), .A(n1752), .ZN(n1737) );
  NOR4_X1 U1637 ( .A1(n1748), .A2(n1749), .A3(n1750), .A4(n1751), .ZN(n1738)
         );
  NAND4_X1 U1638 ( .A1(n1754), .A2(n1755), .A3(n1756), .A4(n1757), .ZN(n2037)
         );
  AOI221_X1 U1639 ( .B1(n1960), .B2(\REGISTERS[15][25] ), .C1(DATA_OUT_1[25]), 
        .C2(n1955), .A(n1771), .ZN(n1754) );
  AOI221_X1 U1640 ( .B1(n1972), .B2(\REGISTERS[7][25] ), .C1(n1969), .C2(
        \REGISTERS[10][25] ), .A(n1770), .ZN(n1755) );
  NOR4_X1 U1641 ( .A1(n1766), .A2(n1767), .A3(n1768), .A4(n1769), .ZN(n1756)
         );
  NAND4_X1 U1642 ( .A1(n1772), .A2(n1773), .A3(n1774), .A4(n1775), .ZN(n2038)
         );
  AOI221_X1 U1643 ( .B1(n1960), .B2(\REGISTERS[15][26] ), .C1(DATA_OUT_1[26]), 
        .C2(n1955), .A(n1789), .ZN(n1772) );
  AOI221_X1 U1644 ( .B1(n1972), .B2(\REGISTERS[7][26] ), .C1(n1969), .C2(
        \REGISTERS[10][26] ), .A(n1788), .ZN(n1773) );
  NOR4_X1 U1645 ( .A1(n1784), .A2(n1785), .A3(n1786), .A4(n1787), .ZN(n1774)
         );
  NAND4_X1 U1646 ( .A1(n1790), .A2(n1791), .A3(n1792), .A4(n1793), .ZN(n2039)
         );
  AOI221_X1 U1647 ( .B1(n1960), .B2(\REGISTERS[15][27] ), .C1(DATA_OUT_1[27]), 
        .C2(n1955), .A(n1807), .ZN(n1790) );
  AOI221_X1 U1648 ( .B1(n1972), .B2(\REGISTERS[7][27] ), .C1(n1969), .C2(
        \REGISTERS[10][27] ), .A(n1806), .ZN(n1791) );
  NOR4_X1 U1649 ( .A1(n1802), .A2(n1803), .A3(n1804), .A4(n1805), .ZN(n1792)
         );
  NAND4_X1 U1650 ( .A1(n1808), .A2(n1809), .A3(n1810), .A4(n1811), .ZN(n2040)
         );
  AOI221_X1 U1651 ( .B1(n1960), .B2(\REGISTERS[15][28] ), .C1(DATA_OUT_1[28]), 
        .C2(n1955), .A(n1825), .ZN(n1808) );
  AOI221_X1 U1652 ( .B1(n1972), .B2(\REGISTERS[7][28] ), .C1(n1969), .C2(
        \REGISTERS[10][28] ), .A(n1824), .ZN(n1809) );
  NOR4_X1 U1653 ( .A1(n1820), .A2(n1821), .A3(n1822), .A4(n1823), .ZN(n1810)
         );
  NAND4_X1 U1654 ( .A1(n1826), .A2(n1827), .A3(n1828), .A4(n1829), .ZN(n2041)
         );
  AOI221_X1 U1655 ( .B1(n1960), .B2(\REGISTERS[15][29] ), .C1(DATA_OUT_1[29]), 
        .C2(n1955), .A(n1843), .ZN(n1826) );
  AOI221_X1 U1656 ( .B1(n1972), .B2(\REGISTERS[7][29] ), .C1(n1969), .C2(
        \REGISTERS[10][29] ), .A(n1842), .ZN(n1827) );
  NOR4_X1 U1657 ( .A1(n1838), .A2(n1839), .A3(n1840), .A4(n1841), .ZN(n1828)
         );
  NAND4_X1 U1658 ( .A1(n1844), .A2(n1845), .A3(n1846), .A4(n1847), .ZN(n2042)
         );
  AOI221_X1 U1659 ( .B1(n1960), .B2(\REGISTERS[15][30] ), .C1(DATA_OUT_1[30]), 
        .C2(n1955), .A(n1861), .ZN(n1844) );
  AOI221_X1 U1660 ( .B1(n1972), .B2(\REGISTERS[7][30] ), .C1(n1969), .C2(
        \REGISTERS[10][30] ), .A(n1860), .ZN(n1845) );
  NOR4_X1 U1661 ( .A1(n1856), .A2(n1857), .A3(n1858), .A4(n1859), .ZN(n1846)
         );
  NAND4_X1 U1662 ( .A1(n1862), .A2(n1863), .A3(n1864), .A4(n1865), .ZN(n2043)
         );
  AOI221_X1 U1663 ( .B1(n1960), .B2(\REGISTERS[15][31] ), .C1(DATA_OUT_1[31]), 
        .C2(n1956), .A(n1897), .ZN(n1862) );
  AOI221_X1 U1664 ( .B1(n1972), .B2(\REGISTERS[7][31] ), .C1(n1969), .C2(
        \REGISTERS[10][31] ), .A(n1896), .ZN(n1863) );
  NOR4_X1 U1665 ( .A1(n1889), .A2(n1890), .A3(n1891), .A4(n1892), .ZN(n1864)
         );
  AOI221_X1 U1666 ( .B1(\REGISTERS[15][0] ), .B2(n2125), .C1(DATA_OUT_2[0]), 
        .C2(n2118), .A(n68), .ZN(n2) );
  AOI221_X1 U1667 ( .B1(\REGISTERS[7][0] ), .B2(n2137), .C1(\REGISTERS[10][0] ), .C2(n2134), .A(n61), .ZN(n3) );
  NOR4_X1 U1668 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(n4) );
  INV_X1 U1669 ( .A(ADDR_RD2[3]), .ZN(n1262) );
  INV_X1 U1670 ( .A(ADDR_RD2[0]), .ZN(n1259) );
  INV_X1 U1671 ( .A(ADDR_RD1[3]), .ZN(n1895) );
  INV_X1 U1672 ( .A(ADDR_RD1[0]), .ZN(n1894) );
  INV_X1 U1673 ( .A(ADDR_RD2[1]), .ZN(n1269) );
  INV_X1 U1674 ( .A(ADDR_RD2[2]), .ZN(n1256) );
  AND3_X1 U1675 ( .A1(ADDR_RD2[4]), .A2(n1259), .A3(ADDR_RD2[3]), .ZN(n1241)
         );
  AND3_X1 U1676 ( .A1(ADDR_RD2[4]), .A2(n1262), .A3(ADDR_RD2[0]), .ZN(n1245)
         );
  AND3_X1 U1677 ( .A1(ADDR_RD1[4]), .A2(n1894), .A3(ADDR_RD1[3]), .ZN(n1884)
         );
  AND3_X1 U1678 ( .A1(ADDR_RD1[4]), .A2(n1895), .A3(ADDR_RD1[0]), .ZN(n1886)
         );
  AND3_X1 U1679 ( .A1(ADDR_RD2[0]), .A2(ADDR_RD2[4]), .A3(ADDR_RD2[3]), .ZN(
        n1239) );
  AND3_X1 U1680 ( .A1(ADDR_RD1[0]), .A2(ADDR_RD1[4]), .A3(ADDR_RD1[3]), .ZN(
        n1882) );
  AND3_X1 U1681 ( .A1(n1259), .A2(n1262), .A3(ADDR_RD2[4]), .ZN(n1228) );
  AND3_X1 U1682 ( .A1(n1894), .A2(n1895), .A3(ADDR_RD1[4]), .ZN(n1875) );
  INV_X1 U1683 ( .A(ADDR_RD1[1]), .ZN(n1898) );
  INV_X1 U1684 ( .A(ADDR_RD1[2]), .ZN(n1893) );
  INV_X1 U1685 ( .A(ADDR_WR[2]), .ZN(n1915) );
  INV_X1 U1686 ( .A(ADDR_WR[0]), .ZN(n1913) );
  INV_X1 U1687 ( .A(ADDR_WR[1]), .ZN(n1914) );
  INV_X1 U1688 ( .A(\REGISTERS[9][0] ), .ZN(n11) );
  INV_X1 U1689 ( .A(\REGISTERS[1][0] ), .ZN(n18) );
  INV_X1 U1690 ( .A(\REGISTERS[25][0] ), .ZN(n25) );
  INV_X1 U1691 ( .A(\REGISTERS[9][1] ), .ZN(n81) );
  INV_X1 U1692 ( .A(\REGISTERS[1][1] ), .ZN(n84) );
  INV_X1 U1693 ( .A(\REGISTERS[25][1] ), .ZN(n87) );
  INV_X1 U1694 ( .A(\REGISTERS[17][2] ), .ZN(n128) );
  INV_X1 U1695 ( .A(\REGISTERS[9][2] ), .ZN(n119) );
  INV_X1 U1696 ( .A(\REGISTERS[1][2] ), .ZN(n122) );
  INV_X1 U1697 ( .A(\REGISTERS[25][2] ), .ZN(n125) );
  INV_X1 U1698 ( .A(\REGISTERS[17][3] ), .ZN(n166) );
  INV_X1 U1699 ( .A(\REGISTERS[9][3] ), .ZN(n157) );
  INV_X1 U1700 ( .A(\REGISTERS[1][3] ), .ZN(n160) );
  INV_X1 U1701 ( .A(\REGISTERS[25][3] ), .ZN(n163) );
  INV_X1 U1702 ( .A(\REGISTERS[17][4] ), .ZN(n204) );
  INV_X1 U1703 ( .A(\REGISTERS[9][4] ), .ZN(n195) );
  INV_X1 U1704 ( .A(\REGISTERS[1][4] ), .ZN(n198) );
  INV_X1 U1705 ( .A(\REGISTERS[25][4] ), .ZN(n201) );
  INV_X1 U1706 ( .A(\REGISTERS[17][5] ), .ZN(n242) );
  INV_X1 U1707 ( .A(\REGISTERS[9][5] ), .ZN(n233) );
  INV_X1 U1708 ( .A(\REGISTERS[1][5] ), .ZN(n236) );
  INV_X1 U1709 ( .A(\REGISTERS[25][5] ), .ZN(n239) );
  INV_X1 U1710 ( .A(\REGISTERS[17][6] ), .ZN(n280) );
  INV_X1 U1711 ( .A(\REGISTERS[9][6] ), .ZN(n271) );
  INV_X1 U1712 ( .A(\REGISTERS[1][6] ), .ZN(n274) );
  INV_X1 U1713 ( .A(\REGISTERS[25][6] ), .ZN(n277) );
  INV_X1 U1714 ( .A(\REGISTERS[17][7] ), .ZN(n318) );
  INV_X1 U1715 ( .A(\REGISTERS[9][7] ), .ZN(n309) );
  INV_X1 U1716 ( .A(\REGISTERS[1][7] ), .ZN(n312) );
  INV_X1 U1717 ( .A(\REGISTERS[25][7] ), .ZN(n315) );
  INV_X1 U1718 ( .A(\REGISTERS[17][8] ), .ZN(n356) );
  INV_X1 U1719 ( .A(\REGISTERS[9][8] ), .ZN(n347) );
  INV_X1 U1720 ( .A(\REGISTERS[1][8] ), .ZN(n350) );
  INV_X1 U1721 ( .A(\REGISTERS[25][8] ), .ZN(n353) );
  INV_X1 U1722 ( .A(\REGISTERS[17][9] ), .ZN(n394) );
  INV_X1 U1723 ( .A(\REGISTERS[9][9] ), .ZN(n385) );
  INV_X1 U1724 ( .A(\REGISTERS[1][9] ), .ZN(n388) );
  INV_X1 U1725 ( .A(\REGISTERS[25][9] ), .ZN(n391) );
  INV_X1 U1726 ( .A(\REGISTERS[17][10] ), .ZN(n432) );
  INV_X1 U1727 ( .A(\REGISTERS[9][10] ), .ZN(n423) );
  INV_X1 U1728 ( .A(\REGISTERS[1][10] ), .ZN(n426) );
  INV_X1 U1729 ( .A(\REGISTERS[25][10] ), .ZN(n429) );
  INV_X1 U1730 ( .A(\REGISTERS[17][11] ), .ZN(n470) );
  INV_X1 U1731 ( .A(\REGISTERS[9][11] ), .ZN(n461) );
  INV_X1 U1732 ( .A(\REGISTERS[1][11] ), .ZN(n464) );
  INV_X1 U1733 ( .A(\REGISTERS[25][11] ), .ZN(n467) );
  INV_X1 U1734 ( .A(\REGISTERS[17][12] ), .ZN(n508) );
  INV_X1 U1735 ( .A(\REGISTERS[9][12] ), .ZN(n499) );
  INV_X1 U1736 ( .A(\REGISTERS[1][12] ), .ZN(n502) );
  INV_X1 U1737 ( .A(\REGISTERS[25][12] ), .ZN(n505) );
  INV_X1 U1738 ( .A(\REGISTERS[17][13] ), .ZN(n546) );
  INV_X1 U1739 ( .A(\REGISTERS[9][13] ), .ZN(n537) );
  INV_X1 U1740 ( .A(\REGISTERS[1][13] ), .ZN(n540) );
  INV_X1 U1741 ( .A(\REGISTERS[25][13] ), .ZN(n543) );
  INV_X1 U1742 ( .A(\REGISTERS[17][14] ), .ZN(n584) );
  INV_X1 U1743 ( .A(\REGISTERS[9][14] ), .ZN(n575) );
  INV_X1 U1744 ( .A(\REGISTERS[1][14] ), .ZN(n578) );
  INV_X1 U1745 ( .A(\REGISTERS[25][14] ), .ZN(n581) );
  INV_X1 U1746 ( .A(\REGISTERS[17][15] ), .ZN(n622) );
  INV_X1 U1747 ( .A(\REGISTERS[9][15] ), .ZN(n613) );
  INV_X1 U1748 ( .A(\REGISTERS[1][15] ), .ZN(n616) );
  INV_X1 U1749 ( .A(\REGISTERS[25][15] ), .ZN(n619) );
  INV_X1 U1750 ( .A(\REGISTERS[17][16] ), .ZN(n660) );
  INV_X1 U1751 ( .A(\REGISTERS[9][16] ), .ZN(n651) );
  INV_X1 U1752 ( .A(\REGISTERS[1][16] ), .ZN(n654) );
  INV_X1 U1753 ( .A(\REGISTERS[25][16] ), .ZN(n657) );
  INV_X1 U1754 ( .A(\REGISTERS[17][17] ), .ZN(n698) );
  INV_X1 U1755 ( .A(\REGISTERS[9][17] ), .ZN(n689) );
  INV_X1 U1756 ( .A(\REGISTERS[1][17] ), .ZN(n692) );
  INV_X1 U1757 ( .A(\REGISTERS[25][17] ), .ZN(n695) );
  INV_X1 U1758 ( .A(\REGISTERS[17][18] ), .ZN(n736) );
  INV_X1 U1759 ( .A(\REGISTERS[9][18] ), .ZN(n727) );
  INV_X1 U1760 ( .A(\REGISTERS[1][18] ), .ZN(n730) );
  INV_X1 U1761 ( .A(\REGISTERS[25][18] ), .ZN(n733) );
  INV_X1 U1762 ( .A(\REGISTERS[17][19] ), .ZN(n774) );
  INV_X1 U1763 ( .A(\REGISTERS[9][19] ), .ZN(n765) );
  INV_X1 U1764 ( .A(\REGISTERS[1][19] ), .ZN(n768) );
  INV_X1 U1765 ( .A(\REGISTERS[25][19] ), .ZN(n771) );
  INV_X1 U1766 ( .A(\REGISTERS[17][20] ), .ZN(n812) );
  INV_X1 U1767 ( .A(\REGISTERS[9][20] ), .ZN(n803) );
  INV_X1 U1768 ( .A(\REGISTERS[1][20] ), .ZN(n806) );
  INV_X1 U1769 ( .A(\REGISTERS[25][20] ), .ZN(n809) );
  INV_X1 U1770 ( .A(\REGISTERS[17][21] ), .ZN(n850) );
  INV_X1 U1771 ( .A(\REGISTERS[9][21] ), .ZN(n841) );
  INV_X1 U1772 ( .A(\REGISTERS[1][21] ), .ZN(n844) );
  INV_X1 U1773 ( .A(\REGISTERS[25][21] ), .ZN(n847) );
  INV_X1 U1774 ( .A(\REGISTERS[17][22] ), .ZN(n888) );
  INV_X1 U1775 ( .A(\REGISTERS[9][22] ), .ZN(n879) );
  INV_X1 U1776 ( .A(\REGISTERS[1][22] ), .ZN(n882) );
  INV_X1 U1777 ( .A(\REGISTERS[25][22] ), .ZN(n885) );
  INV_X1 U1778 ( .A(\REGISTERS[17][23] ), .ZN(n926) );
  INV_X1 U1779 ( .A(\REGISTERS[9][23] ), .ZN(n917) );
  INV_X1 U1780 ( .A(\REGISTERS[1][23] ), .ZN(n920) );
  INV_X1 U1781 ( .A(\REGISTERS[25][23] ), .ZN(n923) );
  INV_X1 U1782 ( .A(\REGISTERS[17][24] ), .ZN(n964) );
  INV_X1 U1783 ( .A(\REGISTERS[9][24] ), .ZN(n955) );
  INV_X1 U1784 ( .A(\REGISTERS[1][24] ), .ZN(n958) );
  INV_X1 U1785 ( .A(\REGISTERS[25][24] ), .ZN(n961) );
  INV_X1 U1786 ( .A(\REGISTERS[17][25] ), .ZN(n1002) );
  INV_X1 U1787 ( .A(\REGISTERS[9][25] ), .ZN(n993) );
  INV_X1 U1788 ( .A(\REGISTERS[1][25] ), .ZN(n996) );
  INV_X1 U1789 ( .A(\REGISTERS[25][25] ), .ZN(n999) );
  INV_X1 U1790 ( .A(\REGISTERS[17][26] ), .ZN(n1040) );
  INV_X1 U1791 ( .A(\REGISTERS[9][26] ), .ZN(n1031) );
  INV_X1 U1792 ( .A(\REGISTERS[1][26] ), .ZN(n1034) );
  INV_X1 U1793 ( .A(\REGISTERS[25][26] ), .ZN(n1037) );
  INV_X1 U1794 ( .A(\REGISTERS[17][27] ), .ZN(n1078) );
  INV_X1 U1795 ( .A(\REGISTERS[9][27] ), .ZN(n1069) );
  INV_X1 U1796 ( .A(\REGISTERS[1][27] ), .ZN(n1072) );
  INV_X1 U1797 ( .A(\REGISTERS[25][27] ), .ZN(n1075) );
  INV_X1 U1798 ( .A(\REGISTERS[17][28] ), .ZN(n1116) );
  INV_X1 U1799 ( .A(\REGISTERS[9][28] ), .ZN(n1107) );
  INV_X1 U1800 ( .A(\REGISTERS[1][28] ), .ZN(n1110) );
  INV_X1 U1801 ( .A(\REGISTERS[25][28] ), .ZN(n1113) );
  INV_X1 U1802 ( .A(\REGISTERS[17][29] ), .ZN(n1154) );
  INV_X1 U1803 ( .A(\REGISTERS[9][29] ), .ZN(n1145) );
  INV_X1 U1804 ( .A(\REGISTERS[1][29] ), .ZN(n1148) );
  INV_X1 U1805 ( .A(\REGISTERS[25][29] ), .ZN(n1151) );
  INV_X1 U1806 ( .A(\REGISTERS[17][30] ), .ZN(n1192) );
  INV_X1 U1807 ( .A(\REGISTERS[9][30] ), .ZN(n1183) );
  INV_X1 U1808 ( .A(\REGISTERS[1][30] ), .ZN(n1186) );
  INV_X1 U1809 ( .A(\REGISTERS[25][30] ), .ZN(n1189) );
  INV_X1 U1810 ( .A(\REGISTERS[17][31] ), .ZN(n1242) );
  INV_X1 U1811 ( .A(\REGISTERS[9][31] ), .ZN(n1221) );
  INV_X1 U1812 ( .A(\REGISTERS[1][31] ), .ZN(n1231) );
  INV_X1 U1813 ( .A(\REGISTERS[25][31] ), .ZN(n1236) );
  INV_X1 U1814 ( .A(\REGISTERS[2][0] ), .ZN(n44) );
  INV_X1 U1815 ( .A(\REGISTERS[28][0] ), .ZN(n48) );
  INV_X1 U1816 ( .A(\REGISTERS[26][0] ), .ZN(n52) );
  INV_X1 U1817 ( .A(\REGISTERS[22][0] ), .ZN(n56) );
  INV_X1 U1818 ( .A(\REGISTERS[6][0] ), .ZN(n63) );
  INV_X1 U1819 ( .A(\REGISTERS[14][0] ), .ZN(n70) );
  INV_X1 U1820 ( .A(\REGISTERS[2][1] ), .ZN(n97) );
  INV_X1 U1821 ( .A(\REGISTERS[28][1] ), .ZN(n99) );
  INV_X1 U1822 ( .A(\REGISTERS[26][1] ), .ZN(n101) );
  INV_X1 U1823 ( .A(\REGISTERS[22][1] ), .ZN(n103) );
  INV_X1 U1824 ( .A(\REGISTERS[6][1] ), .ZN(n106) );
  INV_X1 U1825 ( .A(\REGISTERS[14][1] ), .ZN(n109) );
  INV_X1 U1826 ( .A(\REGISTERS[2][2] ), .ZN(n135) );
  INV_X1 U1827 ( .A(\REGISTERS[28][2] ), .ZN(n137) );
  INV_X1 U1828 ( .A(\REGISTERS[26][2] ), .ZN(n139) );
  INV_X1 U1829 ( .A(\REGISTERS[22][2] ), .ZN(n141) );
  INV_X1 U1830 ( .A(\REGISTERS[6][2] ), .ZN(n144) );
  INV_X1 U1831 ( .A(\REGISTERS[14][2] ), .ZN(n147) );
  INV_X1 U1832 ( .A(\REGISTERS[2][3] ), .ZN(n173) );
  INV_X1 U1833 ( .A(\REGISTERS[28][3] ), .ZN(n175) );
  INV_X1 U1834 ( .A(\REGISTERS[26][3] ), .ZN(n177) );
  INV_X1 U1835 ( .A(\REGISTERS[22][3] ), .ZN(n179) );
  INV_X1 U1836 ( .A(\REGISTERS[6][3] ), .ZN(n182) );
  INV_X1 U1837 ( .A(\REGISTERS[14][3] ), .ZN(n185) );
  INV_X1 U1838 ( .A(\REGISTERS[2][4] ), .ZN(n211) );
  INV_X1 U1839 ( .A(\REGISTERS[28][4] ), .ZN(n213) );
  INV_X1 U1840 ( .A(\REGISTERS[26][4] ), .ZN(n215) );
  INV_X1 U1841 ( .A(\REGISTERS[22][4] ), .ZN(n217) );
  INV_X1 U1842 ( .A(\REGISTERS[6][4] ), .ZN(n220) );
  INV_X1 U1843 ( .A(\REGISTERS[14][4] ), .ZN(n223) );
  INV_X1 U1844 ( .A(\REGISTERS[2][5] ), .ZN(n249) );
  INV_X1 U1845 ( .A(\REGISTERS[28][5] ), .ZN(n251) );
  INV_X1 U1846 ( .A(\REGISTERS[26][5] ), .ZN(n253) );
  INV_X1 U1847 ( .A(\REGISTERS[22][5] ), .ZN(n255) );
  INV_X1 U1848 ( .A(\REGISTERS[6][5] ), .ZN(n258) );
  INV_X1 U1849 ( .A(\REGISTERS[14][5] ), .ZN(n261) );
  INV_X1 U1850 ( .A(\REGISTERS[2][6] ), .ZN(n287) );
  INV_X1 U1851 ( .A(\REGISTERS[28][6] ), .ZN(n289) );
  INV_X1 U1852 ( .A(\REGISTERS[26][6] ), .ZN(n291) );
  INV_X1 U1853 ( .A(\REGISTERS[22][6] ), .ZN(n293) );
  INV_X1 U1854 ( .A(\REGISTERS[6][6] ), .ZN(n296) );
  INV_X1 U1855 ( .A(\REGISTERS[14][6] ), .ZN(n299) );
  INV_X1 U1856 ( .A(\REGISTERS[2][7] ), .ZN(n325) );
  INV_X1 U1857 ( .A(\REGISTERS[28][7] ), .ZN(n327) );
  INV_X1 U1858 ( .A(\REGISTERS[26][7] ), .ZN(n329) );
  INV_X1 U1859 ( .A(\REGISTERS[22][7] ), .ZN(n331) );
  INV_X1 U1860 ( .A(\REGISTERS[6][7] ), .ZN(n334) );
  INV_X1 U1861 ( .A(\REGISTERS[14][7] ), .ZN(n337) );
  INV_X1 U1862 ( .A(\REGISTERS[2][8] ), .ZN(n363) );
  INV_X1 U1863 ( .A(\REGISTERS[28][8] ), .ZN(n365) );
  INV_X1 U1864 ( .A(\REGISTERS[26][8] ), .ZN(n367) );
  INV_X1 U1865 ( .A(\REGISTERS[22][8] ), .ZN(n369) );
  INV_X1 U1866 ( .A(\REGISTERS[6][8] ), .ZN(n372) );
  INV_X1 U1867 ( .A(\REGISTERS[14][8] ), .ZN(n375) );
  INV_X1 U1868 ( .A(\REGISTERS[2][9] ), .ZN(n401) );
  INV_X1 U1869 ( .A(\REGISTERS[28][9] ), .ZN(n403) );
  INV_X1 U1870 ( .A(\REGISTERS[26][9] ), .ZN(n405) );
  INV_X1 U1871 ( .A(\REGISTERS[22][9] ), .ZN(n407) );
  INV_X1 U1872 ( .A(\REGISTERS[6][9] ), .ZN(n410) );
  INV_X1 U1873 ( .A(\REGISTERS[14][9] ), .ZN(n413) );
  INV_X1 U1874 ( .A(\REGISTERS[2][10] ), .ZN(n439) );
  INV_X1 U1875 ( .A(\REGISTERS[28][10] ), .ZN(n441) );
  INV_X1 U1876 ( .A(\REGISTERS[26][10] ), .ZN(n443) );
  INV_X1 U1877 ( .A(\REGISTERS[22][10] ), .ZN(n445) );
  INV_X1 U1879 ( .A(\REGISTERS[6][10] ), .ZN(n448) );
  INV_X1 U1881 ( .A(\REGISTERS[14][10] ), .ZN(n451) );
  INV_X1 U1882 ( .A(\REGISTERS[2][11] ), .ZN(n477) );
  INV_X1 U1883 ( .A(\REGISTERS[28][11] ), .ZN(n479) );
  INV_X1 U1884 ( .A(\REGISTERS[26][11] ), .ZN(n481) );
  INV_X1 U1885 ( .A(\REGISTERS[22][11] ), .ZN(n483) );
  INV_X1 U1887 ( .A(\REGISTERS[6][11] ), .ZN(n486) );
  INV_X1 U1889 ( .A(\REGISTERS[14][11] ), .ZN(n489) );
  INV_X1 U1890 ( .A(\REGISTERS[2][12] ), .ZN(n515) );
  INV_X1 U1891 ( .A(\REGISTERS[28][12] ), .ZN(n517) );
  INV_X1 U1892 ( .A(\REGISTERS[26][12] ), .ZN(n519) );
  INV_X1 U1893 ( .A(\REGISTERS[22][12] ), .ZN(n521) );
  INV_X1 U1895 ( .A(\REGISTERS[6][12] ), .ZN(n524) );
  INV_X1 U1897 ( .A(\REGISTERS[14][12] ), .ZN(n527) );
  INV_X1 U1898 ( .A(\REGISTERS[2][13] ), .ZN(n553) );
  INV_X1 U1899 ( .A(\REGISTERS[28][13] ), .ZN(n555) );
  INV_X1 U1900 ( .A(\REGISTERS[26][13] ), .ZN(n557) );
  INV_X1 U1901 ( .A(\REGISTERS[22][13] ), .ZN(n559) );
  INV_X1 U1902 ( .A(\REGISTERS[6][13] ), .ZN(n562) );
  INV_X1 U1903 ( .A(\REGISTERS[14][13] ), .ZN(n565) );
  INV_X1 U1905 ( .A(\REGISTERS[2][14] ), .ZN(n591) );
  INV_X1 U1906 ( .A(\REGISTERS[28][14] ), .ZN(n593) );
  INV_X1 U1908 ( .A(\REGISTERS[26][14] ), .ZN(n595) );
  INV_X1 U1909 ( .A(\REGISTERS[22][14] ), .ZN(n597) );
  INV_X1 U1910 ( .A(\REGISTERS[6][14] ), .ZN(n600) );
  INV_X1 U1911 ( .A(\REGISTERS[14][14] ), .ZN(n603) );
  INV_X1 U1913 ( .A(\REGISTERS[2][15] ), .ZN(n629) );
  INV_X1 U1915 ( .A(\REGISTERS[28][15] ), .ZN(n631) );
  INV_X1 U1916 ( .A(\REGISTERS[26][15] ), .ZN(n633) );
  INV_X1 U1918 ( .A(\REGISTERS[22][15] ), .ZN(n635) );
  INV_X1 U1919 ( .A(\REGISTERS[6][15] ), .ZN(n638) );
  INV_X1 U1921 ( .A(\REGISTERS[14][15] ), .ZN(n641) );
  INV_X1 U1922 ( .A(\REGISTERS[2][16] ), .ZN(n667) );
  INV_X1 U1923 ( .A(\REGISTERS[28][16] ), .ZN(n669) );
  INV_X1 U1925 ( .A(\REGISTERS[26][16] ), .ZN(n671) );
  INV_X1 U1927 ( .A(\REGISTERS[22][16] ), .ZN(n673) );
  INV_X1 U1928 ( .A(\REGISTERS[6][16] ), .ZN(n676) );
  INV_X1 U1929 ( .A(\REGISTERS[14][16] ), .ZN(n679) );
  INV_X1 U1931 ( .A(\REGISTERS[2][17] ), .ZN(n705) );
  INV_X1 U1932 ( .A(\REGISTERS[28][17] ), .ZN(n707) );
  INV_X1 U1934 ( .A(\REGISTERS[26][17] ), .ZN(n709) );
  INV_X1 U1935 ( .A(\REGISTERS[22][17] ), .ZN(n711) );
  INV_X1 U1936 ( .A(\REGISTERS[6][17] ), .ZN(n714) );
  INV_X1 U1937 ( .A(\REGISTERS[14][17] ), .ZN(n717) );
  INV_X1 U1939 ( .A(\REGISTERS[2][18] ), .ZN(n743) );
  INV_X1 U1941 ( .A(\REGISTERS[28][18] ), .ZN(n745) );
  INV_X1 U1942 ( .A(\REGISTERS[26][18] ), .ZN(n747) );
  INV_X1 U1943 ( .A(\REGISTERS[22][18] ), .ZN(n749) );
  INV_X1 U1944 ( .A(\REGISTERS[6][18] ), .ZN(n752) );
  INV_X1 U1945 ( .A(\REGISTERS[14][18] ), .ZN(n755) );
  INV_X1 U1946 ( .A(\REGISTERS[2][19] ), .ZN(n781) );
  INV_X1 U1947 ( .A(\REGISTERS[28][19] ), .ZN(n783) );
  INV_X1 U1949 ( .A(\REGISTERS[26][19] ), .ZN(n785) );
  INV_X1 U1950 ( .A(\REGISTERS[22][19] ), .ZN(n787) );
  INV_X1 U1952 ( .A(\REGISTERS[6][19] ), .ZN(n790) );
  INV_X1 U1953 ( .A(\REGISTERS[14][19] ), .ZN(n793) );
  INV_X1 U1954 ( .A(\REGISTERS[2][20] ), .ZN(n819) );
  INV_X1 U1955 ( .A(\REGISTERS[28][20] ), .ZN(n821) );
  INV_X1 U1956 ( .A(\REGISTERS[26][20] ), .ZN(n823) );
  INV_X1 U1957 ( .A(\REGISTERS[22][20] ), .ZN(n825) );
  INV_X1 U1958 ( .A(\REGISTERS[6][20] ), .ZN(n828) );
  INV_X1 U1960 ( .A(\REGISTERS[14][20] ), .ZN(n831) );
  INV_X1 U1961 ( .A(\REGISTERS[2][21] ), .ZN(n857) );
  INV_X1 U1962 ( .A(\REGISTERS[28][21] ), .ZN(n859) );
  INV_X1 U1963 ( .A(\REGISTERS[26][21] ), .ZN(n861) );
  INV_X1 U1964 ( .A(\REGISTERS[22][21] ), .ZN(n863) );
  INV_X1 U1965 ( .A(\REGISTERS[6][21] ), .ZN(n866) );
  INV_X1 U1966 ( .A(\REGISTERS[14][21] ), .ZN(n869) );
  INV_X1 U1967 ( .A(\REGISTERS[2][22] ), .ZN(n895) );
  INV_X1 U1968 ( .A(\REGISTERS[28][22] ), .ZN(n897) );
  INV_X1 U1969 ( .A(\REGISTERS[26][22] ), .ZN(n899) );
  INV_X1 U1970 ( .A(\REGISTERS[22][22] ), .ZN(n901) );
  INV_X1 U1971 ( .A(\REGISTERS[6][22] ), .ZN(n904) );
  INV_X1 U1972 ( .A(\REGISTERS[14][22] ), .ZN(n907) );
  INV_X1 U1973 ( .A(\REGISTERS[2][23] ), .ZN(n933) );
  INV_X1 U1974 ( .A(\REGISTERS[28][23] ), .ZN(n935) );
  INV_X1 U1975 ( .A(\REGISTERS[26][23] ), .ZN(n937) );
  INV_X1 U1976 ( .A(\REGISTERS[22][23] ), .ZN(n939) );
  INV_X1 U1977 ( .A(\REGISTERS[6][23] ), .ZN(n942) );
  INV_X1 U1978 ( .A(\REGISTERS[14][23] ), .ZN(n945) );
  INV_X1 U1979 ( .A(\REGISTERS[2][24] ), .ZN(n971) );
  INV_X1 U1980 ( .A(\REGISTERS[28][24] ), .ZN(n973) );
  INV_X1 U1981 ( .A(\REGISTERS[26][24] ), .ZN(n975) );
  INV_X1 U1982 ( .A(\REGISTERS[22][24] ), .ZN(n977) );
  INV_X1 U1983 ( .A(\REGISTERS[6][24] ), .ZN(n980) );
  INV_X1 U1984 ( .A(\REGISTERS[14][24] ), .ZN(n983) );
  INV_X1 U1985 ( .A(\REGISTERS[2][25] ), .ZN(n1009) );
  INV_X1 U1986 ( .A(\REGISTERS[28][25] ), .ZN(n1011) );
  INV_X1 U1987 ( .A(\REGISTERS[26][25] ), .ZN(n1013) );
  INV_X1 U1988 ( .A(\REGISTERS[22][25] ), .ZN(n1015) );
  INV_X1 U1989 ( .A(\REGISTERS[6][25] ), .ZN(n1018) );
  INV_X1 U1990 ( .A(\REGISTERS[14][25] ), .ZN(n1021) );
  INV_X1 U1991 ( .A(\REGISTERS[2][26] ), .ZN(n1047) );
  INV_X1 U1992 ( .A(\REGISTERS[28][26] ), .ZN(n1049) );
  INV_X1 U1993 ( .A(\REGISTERS[26][26] ), .ZN(n1051) );
  INV_X1 U1994 ( .A(\REGISTERS[22][26] ), .ZN(n1053) );
  INV_X1 U1995 ( .A(\REGISTERS[6][26] ), .ZN(n1056) );
  INV_X1 U1996 ( .A(\REGISTERS[14][26] ), .ZN(n1059) );
  INV_X1 U1997 ( .A(\REGISTERS[2][27] ), .ZN(n1085) );
  INV_X1 U1998 ( .A(\REGISTERS[28][27] ), .ZN(n1087) );
  INV_X1 U1999 ( .A(\REGISTERS[26][27] ), .ZN(n1089) );
  INV_X1 U2000 ( .A(\REGISTERS[22][27] ), .ZN(n1091) );
  INV_X1 U2001 ( .A(\REGISTERS[6][27] ), .ZN(n1094) );
  INV_X1 U2002 ( .A(\REGISTERS[14][27] ), .ZN(n1097) );
  INV_X1 U2004 ( .A(\REGISTERS[2][28] ), .ZN(n1123) );
  INV_X1 U2005 ( .A(\REGISTERS[28][28] ), .ZN(n1125) );
  INV_X1 U2006 ( .A(\REGISTERS[26][28] ), .ZN(n1127) );
  INV_X1 U2007 ( .A(\REGISTERS[22][28] ), .ZN(n1129) );
  INV_X1 U2008 ( .A(\REGISTERS[6][28] ), .ZN(n1132) );
  INV_X1 U2009 ( .A(\REGISTERS[14][28] ), .ZN(n1135) );
  INV_X1 U2010 ( .A(\REGISTERS[2][29] ), .ZN(n1161) );
  INV_X1 U2011 ( .A(\REGISTERS[28][29] ), .ZN(n1163) );
  INV_X1 U2013 ( .A(\REGISTERS[26][29] ), .ZN(n1165) );
  INV_X1 U2014 ( .A(\REGISTERS[22][29] ), .ZN(n1167) );
  INV_X1 U2015 ( .A(\REGISTERS[6][29] ), .ZN(n1170) );
  INV_X1 U2016 ( .A(\REGISTERS[14][29] ), .ZN(n1173) );
  INV_X1 U2017 ( .A(\REGISTERS[2][30] ), .ZN(n1199) );
  INV_X1 U2018 ( .A(\REGISTERS[28][30] ), .ZN(n1201) );
  INV_X1 U2019 ( .A(\REGISTERS[26][30] ), .ZN(n1203) );
  INV_X1 U2020 ( .A(\REGISTERS[22][30] ), .ZN(n1205) );
  INV_X1 U2022 ( .A(\REGISTERS[6][30] ), .ZN(n1208) );
  INV_X1 U2024 ( .A(\REGISTERS[14][30] ), .ZN(n1211) );
  INV_X1 U2026 ( .A(\REGISTERS[2][31] ), .ZN(n1252) );
  INV_X1 U2028 ( .A(\REGISTERS[28][31] ), .ZN(n1254) );
  INV_X1 U2030 ( .A(\REGISTERS[26][31] ), .ZN(n1257) );
  INV_X1 U2032 ( .A(\REGISTERS[22][31] ), .ZN(n1260) );
  INV_X1 U2034 ( .A(\REGISTERS[6][31] ), .ZN(n1264) );
  INV_X1 U2036 ( .A(\REGISTERS[14][31] ), .ZN(n1267) );
  INV_X1 U2037 ( .A(\REGISTERS[29][0] ), .ZN(n46) );
  INV_X1 U2039 ( .A(\REGISTERS[27][0] ), .ZN(n50) );
  INV_X1 U2040 ( .A(\REGISTERS[23][0] ), .ZN(n54) );
  INV_X1 U2042 ( .A(\REGISTERS[19][0] ), .ZN(n58) );
  INV_X1 U2043 ( .A(\REGISTERS[3][0] ), .ZN(n65) );
  INV_X1 U2044 ( .A(\REGISTERS[11][0] ), .ZN(n72) );
  INV_X1 U2046 ( .A(\REGISTERS[29][1] ), .ZN(n98) );
  INV_X1 U2047 ( .A(\REGISTERS[27][1] ), .ZN(n100) );
  INV_X1 U2048 ( .A(\REGISTERS[23][1] ), .ZN(n102) );
  INV_X1 U2049 ( .A(\REGISTERS[19][1] ), .ZN(n104) );
  INV_X1 U2050 ( .A(\REGISTERS[3][1] ), .ZN(n107) );
  INV_X1 U2051 ( .A(\REGISTERS[11][1] ), .ZN(n110) );
  INV_X1 U2052 ( .A(\REGISTERS[29][2] ), .ZN(n136) );
  INV_X1 U2053 ( .A(\REGISTERS[27][2] ), .ZN(n138) );
  INV_X1 U2054 ( .A(\REGISTERS[23][2] ), .ZN(n140) );
  INV_X1 U2055 ( .A(\REGISTERS[19][2] ), .ZN(n142) );
  INV_X1 U2056 ( .A(\REGISTERS[3][2] ), .ZN(n145) );
  INV_X1 U2057 ( .A(\REGISTERS[11][2] ), .ZN(n148) );
  INV_X1 U2058 ( .A(\REGISTERS[29][3] ), .ZN(n174) );
  INV_X1 U2059 ( .A(\REGISTERS[27][3] ), .ZN(n176) );
  INV_X1 U2060 ( .A(\REGISTERS[23][3] ), .ZN(n178) );
  INV_X1 U2061 ( .A(\REGISTERS[19][3] ), .ZN(n180) );
  INV_X1 U2062 ( .A(\REGISTERS[3][3] ), .ZN(n183) );
  INV_X1 U2063 ( .A(\REGISTERS[11][3] ), .ZN(n186) );
  INV_X1 U2064 ( .A(\REGISTERS[29][4] ), .ZN(n212) );
  INV_X1 U2065 ( .A(\REGISTERS[27][4] ), .ZN(n214) );
  INV_X1 U2066 ( .A(\REGISTERS[23][4] ), .ZN(n216) );
  INV_X1 U2067 ( .A(\REGISTERS[19][4] ), .ZN(n218) );
  INV_X1 U2068 ( .A(\REGISTERS[3][4] ), .ZN(n221) );
  INV_X1 U2069 ( .A(\REGISTERS[11][4] ), .ZN(n224) );
  INV_X1 U2070 ( .A(\REGISTERS[29][5] ), .ZN(n250) );
  INV_X1 U2071 ( .A(\REGISTERS[27][5] ), .ZN(n252) );
  INV_X1 U2072 ( .A(\REGISTERS[23][5] ), .ZN(n254) );
  INV_X1 U2073 ( .A(\REGISTERS[19][5] ), .ZN(n256) );
  INV_X1 U2074 ( .A(\REGISTERS[3][5] ), .ZN(n259) );
  INV_X1 U2075 ( .A(\REGISTERS[11][5] ), .ZN(n262) );
  INV_X1 U2076 ( .A(\REGISTERS[29][6] ), .ZN(n288) );
  INV_X1 U2077 ( .A(\REGISTERS[27][6] ), .ZN(n290) );
  INV_X1 U2078 ( .A(\REGISTERS[23][6] ), .ZN(n292) );
  INV_X1 U2079 ( .A(\REGISTERS[19][6] ), .ZN(n294) );
  INV_X1 U2080 ( .A(\REGISTERS[3][6] ), .ZN(n297) );
  INV_X1 U2081 ( .A(\REGISTERS[11][6] ), .ZN(n300) );
  INV_X1 U2082 ( .A(\REGISTERS[29][7] ), .ZN(n326) );
  INV_X1 U2083 ( .A(\REGISTERS[27][7] ), .ZN(n328) );
  INV_X1 U2084 ( .A(\REGISTERS[23][7] ), .ZN(n330) );
  INV_X1 U2085 ( .A(\REGISTERS[19][7] ), .ZN(n332) );
  INV_X1 U2086 ( .A(\REGISTERS[3][7] ), .ZN(n335) );
  INV_X1 U2087 ( .A(\REGISTERS[11][7] ), .ZN(n338) );
  INV_X1 U2088 ( .A(\REGISTERS[29][8] ), .ZN(n364) );
  INV_X1 U2089 ( .A(\REGISTERS[27][8] ), .ZN(n366) );
  INV_X1 U2090 ( .A(\REGISTERS[23][8] ), .ZN(n368) );
  INV_X1 U2091 ( .A(\REGISTERS[19][8] ), .ZN(n370) );
  INV_X1 U2092 ( .A(\REGISTERS[3][8] ), .ZN(n373) );
  INV_X1 U2093 ( .A(\REGISTERS[11][8] ), .ZN(n376) );
  INV_X1 U2094 ( .A(\REGISTERS[29][9] ), .ZN(n402) );
  INV_X1 U2095 ( .A(\REGISTERS[27][9] ), .ZN(n404) );
  INV_X1 U2096 ( .A(\REGISTERS[23][9] ), .ZN(n406) );
  INV_X1 U2097 ( .A(\REGISTERS[19][9] ), .ZN(n408) );
  INV_X1 U2098 ( .A(\REGISTERS[3][9] ), .ZN(n411) );
  INV_X1 U2099 ( .A(\REGISTERS[11][9] ), .ZN(n414) );
  INV_X1 U2100 ( .A(\REGISTERS[29][10] ), .ZN(n440) );
  INV_X1 U2101 ( .A(\REGISTERS[27][10] ), .ZN(n442) );
  INV_X1 U2102 ( .A(\REGISTERS[23][10] ), .ZN(n444) );
  INV_X1 U2103 ( .A(\REGISTERS[19][10] ), .ZN(n446) );
  INV_X1 U2104 ( .A(\REGISTERS[3][10] ), .ZN(n449) );
  INV_X1 U2105 ( .A(\REGISTERS[11][10] ), .ZN(n452) );
  INV_X1 U2106 ( .A(\REGISTERS[29][11] ), .ZN(n478) );
  INV_X1 U2107 ( .A(\REGISTERS[27][11] ), .ZN(n480) );
  INV_X1 U2108 ( .A(\REGISTERS[23][11] ), .ZN(n482) );
  INV_X1 U2109 ( .A(\REGISTERS[19][11] ), .ZN(n484) );
  INV_X1 U2110 ( .A(\REGISTERS[3][11] ), .ZN(n487) );
  INV_X1 U2111 ( .A(\REGISTERS[11][11] ), .ZN(n490) );
  INV_X1 U2112 ( .A(\REGISTERS[29][12] ), .ZN(n516) );
  INV_X1 U2113 ( .A(\REGISTERS[27][12] ), .ZN(n518) );
  INV_X1 U2114 ( .A(\REGISTERS[23][12] ), .ZN(n520) );
  INV_X1 U2115 ( .A(\REGISTERS[19][12] ), .ZN(n522) );
  INV_X1 U2116 ( .A(\REGISTERS[3][12] ), .ZN(n525) );
  INV_X1 U2117 ( .A(\REGISTERS[11][12] ), .ZN(n528) );
  INV_X1 U2118 ( .A(\REGISTERS[29][13] ), .ZN(n554) );
  INV_X1 U2119 ( .A(\REGISTERS[27][13] ), .ZN(n556) );
  INV_X1 U2120 ( .A(\REGISTERS[23][13] ), .ZN(n558) );
  INV_X1 U2121 ( .A(\REGISTERS[19][13] ), .ZN(n560) );
  INV_X1 U2122 ( .A(\REGISTERS[3][13] ), .ZN(n563) );
  INV_X1 U2123 ( .A(\REGISTERS[11][13] ), .ZN(n566) );
  INV_X1 U2124 ( .A(\REGISTERS[29][14] ), .ZN(n592) );
  INV_X1 U2125 ( .A(\REGISTERS[27][14] ), .ZN(n594) );
  INV_X1 U2126 ( .A(\REGISTERS[23][14] ), .ZN(n596) );
  INV_X1 U2127 ( .A(\REGISTERS[19][14] ), .ZN(n598) );
  INV_X1 U2128 ( .A(\REGISTERS[3][14] ), .ZN(n601) );
  INV_X1 U2129 ( .A(\REGISTERS[11][14] ), .ZN(n604) );
  INV_X1 U2130 ( .A(\REGISTERS[29][15] ), .ZN(n630) );
  INV_X1 U2131 ( .A(\REGISTERS[27][15] ), .ZN(n632) );
  INV_X1 U2132 ( .A(\REGISTERS[23][15] ), .ZN(n634) );
  INV_X1 U2133 ( .A(\REGISTERS[19][15] ), .ZN(n636) );
  INV_X1 U2134 ( .A(\REGISTERS[3][15] ), .ZN(n639) );
  INV_X1 U2135 ( .A(\REGISTERS[11][15] ), .ZN(n642) );
  INV_X1 U2136 ( .A(\REGISTERS[29][16] ), .ZN(n668) );
  INV_X1 U2137 ( .A(\REGISTERS[27][16] ), .ZN(n670) );
  INV_X1 U2138 ( .A(\REGISTERS[23][16] ), .ZN(n672) );
  INV_X1 U2139 ( .A(\REGISTERS[19][16] ), .ZN(n674) );
  INV_X1 U2140 ( .A(\REGISTERS[3][16] ), .ZN(n677) );
  INV_X1 U2141 ( .A(\REGISTERS[11][16] ), .ZN(n680) );
  INV_X1 U2142 ( .A(\REGISTERS[29][17] ), .ZN(n706) );
  INV_X1 U2143 ( .A(\REGISTERS[27][17] ), .ZN(n708) );
  INV_X1 U2144 ( .A(\REGISTERS[23][17] ), .ZN(n710) );
  INV_X1 U2145 ( .A(\REGISTERS[19][17] ), .ZN(n712) );
  INV_X1 U2146 ( .A(\REGISTERS[3][17] ), .ZN(n715) );
  INV_X1 U2147 ( .A(\REGISTERS[11][17] ), .ZN(n718) );
  INV_X1 U2148 ( .A(\REGISTERS[29][18] ), .ZN(n744) );
  INV_X1 U2149 ( .A(\REGISTERS[27][18] ), .ZN(n746) );
  INV_X1 U2150 ( .A(\REGISTERS[23][18] ), .ZN(n748) );
  INV_X1 U2151 ( .A(\REGISTERS[19][18] ), .ZN(n750) );
  INV_X1 U2152 ( .A(\REGISTERS[3][18] ), .ZN(n753) );
  INV_X1 U2153 ( .A(\REGISTERS[11][18] ), .ZN(n756) );
  INV_X1 U2154 ( .A(\REGISTERS[29][19] ), .ZN(n782) );
  INV_X1 U2155 ( .A(\REGISTERS[27][19] ), .ZN(n784) );
  INV_X1 U2156 ( .A(\REGISTERS[23][19] ), .ZN(n786) );
  INV_X1 U2157 ( .A(\REGISTERS[19][19] ), .ZN(n788) );
  INV_X1 U2158 ( .A(\REGISTERS[3][19] ), .ZN(n791) );
  INV_X1 U2159 ( .A(\REGISTERS[11][19] ), .ZN(n794) );
  INV_X1 U2160 ( .A(\REGISTERS[29][20] ), .ZN(n820) );
  INV_X1 U2161 ( .A(\REGISTERS[27][20] ), .ZN(n822) );
  INV_X1 U2162 ( .A(\REGISTERS[23][20] ), .ZN(n824) );
  INV_X1 U2163 ( .A(\REGISTERS[19][20] ), .ZN(n826) );
  INV_X1 U2164 ( .A(\REGISTERS[3][20] ), .ZN(n829) );
  INV_X1 U2165 ( .A(\REGISTERS[11][20] ), .ZN(n832) );
  INV_X1 U2166 ( .A(\REGISTERS[29][21] ), .ZN(n858) );
  INV_X1 U2167 ( .A(\REGISTERS[27][21] ), .ZN(n860) );
  INV_X1 U2168 ( .A(\REGISTERS[23][21] ), .ZN(n862) );
  INV_X1 U2169 ( .A(\REGISTERS[19][21] ), .ZN(n864) );
  INV_X1 U2170 ( .A(\REGISTERS[3][21] ), .ZN(n867) );
  INV_X1 U2171 ( .A(\REGISTERS[11][21] ), .ZN(n870) );
  INV_X1 U2172 ( .A(\REGISTERS[29][22] ), .ZN(n896) );
  INV_X1 U2173 ( .A(\REGISTERS[27][22] ), .ZN(n898) );
  INV_X1 U2174 ( .A(\REGISTERS[23][22] ), .ZN(n900) );
  INV_X1 U2175 ( .A(\REGISTERS[19][22] ), .ZN(n902) );
  INV_X1 U2176 ( .A(\REGISTERS[3][22] ), .ZN(n905) );
  INV_X1 U2177 ( .A(\REGISTERS[11][22] ), .ZN(n908) );
  INV_X1 U2178 ( .A(\REGISTERS[29][23] ), .ZN(n934) );
  INV_X1 U2179 ( .A(\REGISTERS[27][23] ), .ZN(n936) );
  INV_X1 U2180 ( .A(\REGISTERS[23][23] ), .ZN(n938) );
  INV_X1 U2181 ( .A(\REGISTERS[19][23] ), .ZN(n940) );
  INV_X1 U2182 ( .A(\REGISTERS[3][23] ), .ZN(n943) );
  INV_X1 U2183 ( .A(\REGISTERS[11][23] ), .ZN(n946) );
  INV_X1 U2184 ( .A(\REGISTERS[29][24] ), .ZN(n972) );
  INV_X1 U2185 ( .A(\REGISTERS[27][24] ), .ZN(n974) );
  INV_X1 U2186 ( .A(\REGISTERS[23][24] ), .ZN(n976) );
  INV_X1 U2187 ( .A(\REGISTERS[19][24] ), .ZN(n978) );
  INV_X1 U2188 ( .A(\REGISTERS[3][24] ), .ZN(n981) );
  INV_X1 U2189 ( .A(\REGISTERS[11][24] ), .ZN(n984) );
  INV_X1 U2190 ( .A(\REGISTERS[29][25] ), .ZN(n1010) );
  INV_X1 U2191 ( .A(\REGISTERS[27][25] ), .ZN(n1012) );
  INV_X1 U2192 ( .A(\REGISTERS[23][25] ), .ZN(n1014) );
  INV_X1 U2193 ( .A(\REGISTERS[19][25] ), .ZN(n1016) );
  INV_X1 U2194 ( .A(\REGISTERS[3][25] ), .ZN(n1019) );
  INV_X1 U2195 ( .A(\REGISTERS[11][25] ), .ZN(n1022) );
  INV_X1 U2196 ( .A(\REGISTERS[29][26] ), .ZN(n1048) );
  INV_X1 U2197 ( .A(\REGISTERS[27][26] ), .ZN(n1050) );
  INV_X1 U2198 ( .A(\REGISTERS[23][26] ), .ZN(n1052) );
  INV_X1 U2199 ( .A(\REGISTERS[19][26] ), .ZN(n1054) );
  INV_X1 U2200 ( .A(\REGISTERS[3][26] ), .ZN(n1057) );
  INV_X1 U2201 ( .A(\REGISTERS[11][26] ), .ZN(n1060) );
  INV_X1 U2202 ( .A(\REGISTERS[29][27] ), .ZN(n1086) );
  INV_X1 U2203 ( .A(\REGISTERS[27][27] ), .ZN(n1088) );
  INV_X1 U2204 ( .A(\REGISTERS[23][27] ), .ZN(n1090) );
  INV_X1 U2205 ( .A(\REGISTERS[19][27] ), .ZN(n1092) );
  INV_X1 U2206 ( .A(\REGISTERS[3][27] ), .ZN(n1095) );
  INV_X1 U2207 ( .A(\REGISTERS[11][27] ), .ZN(n1098) );
  INV_X1 U2208 ( .A(\REGISTERS[29][28] ), .ZN(n1124) );
  INV_X1 U2209 ( .A(\REGISTERS[27][28] ), .ZN(n1126) );
  INV_X1 U2210 ( .A(\REGISTERS[23][28] ), .ZN(n1128) );
  INV_X1 U2211 ( .A(\REGISTERS[19][28] ), .ZN(n1130) );
  INV_X1 U2212 ( .A(\REGISTERS[3][28] ), .ZN(n1133) );
  INV_X1 U2213 ( .A(\REGISTERS[11][28] ), .ZN(n1136) );
  INV_X1 U2214 ( .A(\REGISTERS[29][29] ), .ZN(n1162) );
  INV_X1 U2215 ( .A(\REGISTERS[27][29] ), .ZN(n1164) );
  INV_X1 U2216 ( .A(\REGISTERS[23][29] ), .ZN(n1166) );
  INV_X1 U2217 ( .A(\REGISTERS[19][29] ), .ZN(n1168) );
  INV_X1 U2218 ( .A(\REGISTERS[3][29] ), .ZN(n1171) );
  INV_X1 U2219 ( .A(\REGISTERS[11][29] ), .ZN(n1174) );
  INV_X1 U2220 ( .A(\REGISTERS[29][30] ), .ZN(n1200) );
  INV_X1 U2221 ( .A(\REGISTERS[27][30] ), .ZN(n1202) );
  INV_X1 U2222 ( .A(\REGISTERS[23][30] ), .ZN(n1204) );
  INV_X1 U2223 ( .A(\REGISTERS[19][30] ), .ZN(n1206) );
  INV_X1 U2224 ( .A(\REGISTERS[3][30] ), .ZN(n1209) );
  INV_X1 U2225 ( .A(\REGISTERS[11][30] ), .ZN(n1212) );
  INV_X1 U2226 ( .A(\REGISTERS[29][31] ), .ZN(n1253) );
  INV_X1 U2227 ( .A(\REGISTERS[27][31] ), .ZN(n1255) );
  INV_X1 U2228 ( .A(\REGISTERS[23][31] ), .ZN(n1258) );
  INV_X1 U2229 ( .A(\REGISTERS[19][31] ), .ZN(n1261) );
  INV_X1 U2230 ( .A(\REGISTERS[3][31] ), .ZN(n1265) );
  INV_X1 U2231 ( .A(\REGISTERS[11][31] ), .ZN(n1268) );
  INV_X1 U2232 ( .A(\REGISTERS[18][0] ), .ZN(n13) );
  INV_X1 U2233 ( .A(\REGISTERS[12][0] ), .ZN(n20) );
  INV_X1 U2234 ( .A(\REGISTERS[4][0] ), .ZN(n27) );
  INV_X1 U2235 ( .A(\REGISTERS[18][1] ), .ZN(n82) );
  INV_X1 U2236 ( .A(\REGISTERS[12][1] ), .ZN(n85) );
  INV_X1 U2237 ( .A(\REGISTERS[4][1] ), .ZN(n88) );
  INV_X1 U2238 ( .A(\REGISTERS[30][2] ), .ZN(n129) );
  INV_X1 U2239 ( .A(\REGISTERS[18][2] ), .ZN(n120) );
  INV_X1 U2240 ( .A(\REGISTERS[12][2] ), .ZN(n123) );
  INV_X1 U2241 ( .A(\REGISTERS[4][2] ), .ZN(n126) );
  INV_X1 U2242 ( .A(\REGISTERS[30][3] ), .ZN(n167) );
  INV_X1 U2243 ( .A(\REGISTERS[18][3] ), .ZN(n158) );
  INV_X1 U2244 ( .A(\REGISTERS[12][3] ), .ZN(n161) );
  INV_X1 U2245 ( .A(\REGISTERS[4][3] ), .ZN(n164) );
  INV_X1 U2246 ( .A(\REGISTERS[30][4] ), .ZN(n205) );
  INV_X1 U2247 ( .A(\REGISTERS[18][4] ), .ZN(n196) );
  INV_X1 U2248 ( .A(\REGISTERS[12][4] ), .ZN(n199) );
  INV_X1 U2249 ( .A(\REGISTERS[4][4] ), .ZN(n202) );
  INV_X1 U2250 ( .A(\REGISTERS[30][5] ), .ZN(n243) );
  INV_X1 U2251 ( .A(\REGISTERS[18][5] ), .ZN(n234) );
  INV_X1 U2252 ( .A(\REGISTERS[12][5] ), .ZN(n237) );
  INV_X1 U2253 ( .A(\REGISTERS[4][5] ), .ZN(n240) );
  INV_X1 U2254 ( .A(\REGISTERS[30][6] ), .ZN(n281) );
  INV_X1 U2255 ( .A(\REGISTERS[18][6] ), .ZN(n272) );
  INV_X1 U2256 ( .A(\REGISTERS[12][6] ), .ZN(n275) );
  INV_X1 U2257 ( .A(\REGISTERS[4][6] ), .ZN(n278) );
  INV_X1 U2258 ( .A(\REGISTERS[30][7] ), .ZN(n319) );
  INV_X1 U2259 ( .A(\REGISTERS[18][7] ), .ZN(n310) );
  INV_X1 U2260 ( .A(\REGISTERS[12][7] ), .ZN(n313) );
  INV_X1 U2261 ( .A(\REGISTERS[4][7] ), .ZN(n316) );
  INV_X1 U2262 ( .A(\REGISTERS[30][8] ), .ZN(n357) );
  INV_X1 U2263 ( .A(\REGISTERS[18][8] ), .ZN(n348) );
  INV_X1 U2264 ( .A(\REGISTERS[12][8] ), .ZN(n351) );
  INV_X1 U2265 ( .A(\REGISTERS[4][8] ), .ZN(n354) );
  INV_X1 U2266 ( .A(\REGISTERS[30][9] ), .ZN(n395) );
  INV_X1 U2267 ( .A(\REGISTERS[18][9] ), .ZN(n386) );
  INV_X1 U2268 ( .A(\REGISTERS[12][9] ), .ZN(n389) );
  INV_X1 U2269 ( .A(\REGISTERS[4][9] ), .ZN(n392) );
  INV_X1 U2270 ( .A(\REGISTERS[30][10] ), .ZN(n433) );
  INV_X1 U2271 ( .A(\REGISTERS[18][10] ), .ZN(n424) );
  INV_X1 U2272 ( .A(\REGISTERS[12][10] ), .ZN(n427) );
  INV_X1 U2273 ( .A(\REGISTERS[4][10] ), .ZN(n430) );
  INV_X1 U2274 ( .A(\REGISTERS[30][11] ), .ZN(n471) );
  INV_X1 U2275 ( .A(\REGISTERS[18][11] ), .ZN(n462) );
  INV_X1 U2276 ( .A(\REGISTERS[12][11] ), .ZN(n465) );
  INV_X1 U2277 ( .A(\REGISTERS[4][11] ), .ZN(n468) );
  INV_X1 U2278 ( .A(\REGISTERS[30][12] ), .ZN(n509) );
  INV_X1 U2279 ( .A(\REGISTERS[18][12] ), .ZN(n500) );
  INV_X1 U2280 ( .A(\REGISTERS[12][12] ), .ZN(n503) );
  INV_X1 U2281 ( .A(\REGISTERS[4][12] ), .ZN(n506) );
  INV_X1 U2282 ( .A(\REGISTERS[30][13] ), .ZN(n547) );
  INV_X1 U2283 ( .A(\REGISTERS[18][13] ), .ZN(n538) );
  INV_X1 U2284 ( .A(\REGISTERS[12][13] ), .ZN(n541) );
  INV_X1 U2285 ( .A(\REGISTERS[4][13] ), .ZN(n544) );
  INV_X1 U2286 ( .A(\REGISTERS[30][14] ), .ZN(n585) );
  INV_X1 U2287 ( .A(\REGISTERS[18][14] ), .ZN(n576) );
  INV_X1 U2288 ( .A(\REGISTERS[12][14] ), .ZN(n579) );
  INV_X1 U2289 ( .A(\REGISTERS[4][14] ), .ZN(n582) );
  INV_X1 U2290 ( .A(\REGISTERS[30][15] ), .ZN(n623) );
  INV_X1 U2291 ( .A(\REGISTERS[18][15] ), .ZN(n614) );
  INV_X1 U2292 ( .A(\REGISTERS[12][15] ), .ZN(n617) );
  INV_X1 U2293 ( .A(\REGISTERS[4][15] ), .ZN(n620) );
  INV_X1 U2294 ( .A(\REGISTERS[30][16] ), .ZN(n661) );
  INV_X1 U2295 ( .A(\REGISTERS[18][16] ), .ZN(n652) );
  INV_X1 U2296 ( .A(\REGISTERS[12][16] ), .ZN(n655) );
  INV_X1 U2297 ( .A(\REGISTERS[4][16] ), .ZN(n658) );
  INV_X1 U2298 ( .A(\REGISTERS[30][17] ), .ZN(n699) );
  INV_X1 U2299 ( .A(\REGISTERS[18][17] ), .ZN(n690) );
  INV_X1 U2300 ( .A(\REGISTERS[12][17] ), .ZN(n693) );
  INV_X1 U2301 ( .A(\REGISTERS[4][17] ), .ZN(n696) );
  INV_X1 U2302 ( .A(\REGISTERS[30][18] ), .ZN(n737) );
  INV_X1 U2303 ( .A(\REGISTERS[18][18] ), .ZN(n728) );
  INV_X1 U2304 ( .A(\REGISTERS[12][18] ), .ZN(n731) );
  INV_X1 U2305 ( .A(\REGISTERS[4][18] ), .ZN(n734) );
  INV_X1 U2306 ( .A(\REGISTERS[30][19] ), .ZN(n775) );
  INV_X1 U2307 ( .A(\REGISTERS[18][19] ), .ZN(n766) );
  INV_X1 U2308 ( .A(\REGISTERS[12][19] ), .ZN(n769) );
  INV_X1 U2309 ( .A(\REGISTERS[4][19] ), .ZN(n772) );
  INV_X1 U2310 ( .A(\REGISTERS[30][20] ), .ZN(n813) );
  INV_X1 U2311 ( .A(\REGISTERS[18][20] ), .ZN(n804) );
  INV_X1 U2312 ( .A(\REGISTERS[12][20] ), .ZN(n807) );
  INV_X1 U2313 ( .A(\REGISTERS[4][20] ), .ZN(n810) );
  INV_X1 U2314 ( .A(\REGISTERS[30][21] ), .ZN(n851) );
  INV_X1 U2315 ( .A(\REGISTERS[18][21] ), .ZN(n842) );
  INV_X1 U2316 ( .A(\REGISTERS[12][21] ), .ZN(n845) );
  INV_X1 U2317 ( .A(\REGISTERS[4][21] ), .ZN(n848) );
  INV_X1 U2318 ( .A(\REGISTERS[30][22] ), .ZN(n889) );
  INV_X1 U2319 ( .A(\REGISTERS[18][22] ), .ZN(n880) );
  INV_X1 U2320 ( .A(\REGISTERS[12][22] ), .ZN(n883) );
  INV_X1 U2321 ( .A(\REGISTERS[4][22] ), .ZN(n886) );
  INV_X1 U2322 ( .A(\REGISTERS[30][23] ), .ZN(n927) );
  INV_X1 U2323 ( .A(\REGISTERS[18][23] ), .ZN(n918) );
  INV_X1 U2324 ( .A(\REGISTERS[12][23] ), .ZN(n921) );
  INV_X1 U2325 ( .A(\REGISTERS[4][23] ), .ZN(n924) );
  INV_X1 U2326 ( .A(\REGISTERS[30][24] ), .ZN(n965) );
  INV_X1 U2327 ( .A(\REGISTERS[18][24] ), .ZN(n956) );
  INV_X1 U2328 ( .A(\REGISTERS[12][24] ), .ZN(n959) );
  INV_X1 U2329 ( .A(\REGISTERS[4][24] ), .ZN(n962) );
  INV_X1 U2330 ( .A(\REGISTERS[30][25] ), .ZN(n1003) );
  INV_X1 U2331 ( .A(\REGISTERS[18][25] ), .ZN(n994) );
  INV_X1 U2332 ( .A(\REGISTERS[12][25] ), .ZN(n997) );
  INV_X1 U2333 ( .A(\REGISTERS[4][25] ), .ZN(n1000) );
  INV_X1 U2334 ( .A(\REGISTERS[30][26] ), .ZN(n1041) );
  INV_X1 U2335 ( .A(\REGISTERS[18][26] ), .ZN(n1032) );
  INV_X1 U2336 ( .A(\REGISTERS[12][26] ), .ZN(n1035) );
  INV_X1 U2337 ( .A(\REGISTERS[4][26] ), .ZN(n1038) );
  INV_X1 U2338 ( .A(\REGISTERS[30][27] ), .ZN(n1079) );
  INV_X1 U2339 ( .A(\REGISTERS[18][27] ), .ZN(n1070) );
  INV_X1 U2340 ( .A(\REGISTERS[12][27] ), .ZN(n1073) );
  INV_X1 U2341 ( .A(\REGISTERS[4][27] ), .ZN(n1076) );
  INV_X1 U2342 ( .A(\REGISTERS[30][28] ), .ZN(n1117) );
  INV_X1 U2343 ( .A(\REGISTERS[18][28] ), .ZN(n1108) );
  INV_X1 U2344 ( .A(\REGISTERS[12][28] ), .ZN(n1111) );
  INV_X1 U2345 ( .A(\REGISTERS[4][28] ), .ZN(n1114) );
  INV_X1 U2346 ( .A(\REGISTERS[30][29] ), .ZN(n1155) );
  INV_X1 U2347 ( .A(\REGISTERS[18][29] ), .ZN(n1146) );
  INV_X1 U2348 ( .A(\REGISTERS[12][29] ), .ZN(n1149) );
  INV_X1 U2349 ( .A(\REGISTERS[4][29] ), .ZN(n1152) );
  INV_X1 U2350 ( .A(\REGISTERS[30][30] ), .ZN(n1193) );
  INV_X1 U2351 ( .A(\REGISTERS[18][30] ), .ZN(n1184) );
  INV_X1 U2352 ( .A(\REGISTERS[12][30] ), .ZN(n1187) );
  INV_X1 U2353 ( .A(\REGISTERS[4][30] ), .ZN(n1190) );
  INV_X1 U2354 ( .A(\REGISTERS[30][31] ), .ZN(n1243) );
  INV_X1 U2355 ( .A(\REGISTERS[18][31] ), .ZN(n1222) );
  INV_X1 U2356 ( .A(\REGISTERS[12][31] ), .ZN(n1232) );
  INV_X1 U2357 ( .A(\REGISTERS[4][31] ), .ZN(n1237) );
  INV_X1 U2358 ( .A(\REGISTERS[17][0] ), .ZN(n32) );
  INV_X1 U2359 ( .A(\REGISTERS[30][1] ), .ZN(n91) );
  INV_X1 U2360 ( .A(\REGISTERS[17][1] ), .ZN(n90) );
  INV_X1 U2361 ( .A(\REGISTERS[30][0] ), .ZN(n34) );
  INV_X1 U2362 ( .A(ADDR_WR[4]), .ZN(n1911) );
  INV_X1 U2363 ( .A(ADDR_WR[3]), .ZN(n1909) );
  OAI221_X1 U2364 ( .B1(n90), .B2(n2073), .C1(n91), .C2(n2070), .A(n1333), 
        .ZN(n1326) );
  NAND4_X1 U2365 ( .A1(n2), .A2(n3), .A3(n4), .A4(n5), .ZN(n1980) );
  OAI221_X1 U2366 ( .B1(n2172), .B2(n32), .C1(n2169), .C2(n34), .A(n35), .ZN(
        n6) );
  AOI222_X1 U2367 ( .A1(\REGISTERS[21][0] ), .A2(n2168), .B1(
        \REGISTERS[20][0] ), .B2(n2165), .C1(\REGISTERS[16][0] ), .C2(n2164), 
        .ZN(n35) );
  INV_X1 U2368 ( .A(n1318), .ZN(n1957) );
  INV_X1 U2369 ( .A(n1318), .ZN(n1958) );
  INV_X1 U2370 ( .A(n1318), .ZN(n1959) );
  INV_X1 U2371 ( .A(n67), .ZN(n2120) );
  INV_X1 U2372 ( .A(n67), .ZN(n2121) );
  INV_X1 U2373 ( .A(n67), .ZN(n2122) );
endmodule


module N_OR_N3 ( A, Y );
  input [2:0] A;
  output Y;


  OR3_X1 U1 ( .A1(A[2]), .A2(A[1]), .A3(A[0]), .ZN(Y) );
endmodule


module AND_GATE_1_0 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module FD_1_0 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n2, n3, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n2), .ZN(n5) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n3), .ZN(n2) );
  INV_X1 U5 ( .A(EN), .ZN(n3) );
endmodule


module CU_BPU ( HIT_MISS, BRANCH_FETCH, CLK, RST, BRANCH_TAKEN, NEW_BRANCH, 
        EN_FSM );
  input HIT_MISS, BRANCH_FETCH, CLK, RST, BRANCH_TAKEN;
  output NEW_BRANCH, EN_FSM;
  wire   \CURRENT_STATE[1] , N16, N17, n4, n5, n6, n7, n8, n1, n2;

  DFFR_X1 \CURRENT_STATE_reg[0]  ( .D(N16), .CK(CLK), .RN(n2), .QN(n8) );
  DFFR_X1 \CURRENT_STATE_reg[1]  ( .D(N17), .CK(CLK), .RN(n2), .Q(
        \CURRENT_STATE[1] ), .QN(n1) );
  NAND2_X1 U11 ( .A1(\CURRENT_STATE[1] ), .A2(n8), .ZN(n4) );
  NOR3_X1 U3 ( .A1(n5), .A2(HIT_MISS), .A3(n6), .ZN(N17) );
  NOR3_X1 U4 ( .A1(n7), .A2(n6), .A3(n5), .ZN(N16) );
  INV_X1 U5 ( .A(HIT_MISS), .ZN(n7) );
  INV_X1 U6 ( .A(n4), .ZN(NEW_BRANCH) );
  INV_X1 U7 ( .A(BRANCH_FETCH), .ZN(n5) );
  OAI21_X1 U8 ( .B1(\CURRENT_STATE[1] ), .B2(n8), .A(n4), .ZN(EN_FSM) );
  NOR2_X1 U9 ( .A1(n8), .A2(n1), .ZN(n6) );
  INV_X1 U10 ( .A(RST), .ZN(n2) );
endmodule


module FSM_BPU ( RST, CLK, BRANCH_TAKEN, EN_FSM, FSM_SEL, MUX_SEL );
  input [1:0] FSM_SEL;
  input RST, CLK, BRANCH_TAKEN, EN_FSM;
  output MUX_SEL;
  wire   MUX_SEL_A, MUX_SEL_B, MUX_SEL_C, MUX_SEL_D, n2, n3, n4, n5, n6, n8,
         n9, n10, n11, n13, n14, n15, n16, n18, n19, n20, n21, n23, n24, n25,
         n27, n28, n29, n31, n32, n33, n35, n36, n37, n39, n40, n41, n42, n43,
         n44, n45, n47, n48, n49, n50, n51, n1, n7, n12, n17, n22, n26, n30,
         n34, n38;

  DFFR_X1 \CURRENT_STATE_D_reg[0]  ( .D(n47), .CK(CLK), .RN(n38), .Q(n12), 
        .QN(n48) );
  DFFS_X1 \CURRENT_STATE_D_reg[1]  ( .D(n45), .CK(CLK), .SN(n38), .Q(n30), 
        .QN(MUX_SEL_D) );
  DFFR_X1 \CURRENT_STATE_A_reg[0]  ( .D(n44), .CK(CLK), .RN(n38), .Q(n17), 
        .QN(n51) );
  DFFS_X1 \CURRENT_STATE_A_reg[1]  ( .D(n43), .CK(CLK), .SN(n38), .Q(n34), 
        .QN(MUX_SEL_A) );
  DFFR_X1 \CURRENT_STATE_B_reg[0]  ( .D(n42), .CK(CLK), .RN(n38), .Q(n7), .QN(
        n50) );
  DFFS_X1 \CURRENT_STATE_B_reg[1]  ( .D(n41), .CK(CLK), .SN(n38), .Q(n22), 
        .QN(MUX_SEL_B) );
  DFFR_X1 \CURRENT_STATE_C_reg[0]  ( .D(n40), .CK(CLK), .RN(n38), .Q(n1), .QN(
        n49) );
  DFFS_X1 \CURRENT_STATE_C_reg[1]  ( .D(n39), .CK(CLK), .SN(n38), .Q(n26), 
        .QN(MUX_SEL_C) );
  NAND2_X1 U24 ( .A1(BRANCH_TAKEN), .A2(n6), .ZN(n9) );
  NAND3_X1 U27 ( .A1(n51), .A2(n16), .A3(n29), .ZN(n28) );
  NAND2_X1 U31 ( .A1(EN_FSM), .A2(n31), .ZN(n18) );
  NAND2_X1 U38 ( .A1(FSM_SEL[0]), .A2(BRANCH_TAKEN), .ZN(n19) );
  NAND3_X1 U42 ( .A1(n48), .A2(FSM_SEL[0]), .A3(n37), .ZN(n36) );
  NAND2_X1 U45 ( .A1(FSM_SEL[1]), .A2(EN_FSM), .ZN(n8) );
  MUX41_0 MUX_OUT ( .A(MUX_SEL_D), .B(MUX_SEL_C), .C(MUX_SEL_B), .D(MUX_SEL_A), 
        .SEL(FSM_SEL), .Y(MUX_SEL) );
  INV_X1 U3 ( .A(BRANCH_TAKEN), .ZN(n5) );
  INV_X1 U4 ( .A(n18), .ZN(n16) );
  INV_X1 U5 ( .A(n8), .ZN(n4) );
  INV_X1 U6 ( .A(FSM_SEL[1]), .ZN(n31) );
  INV_X1 U7 ( .A(FSM_SEL[0]), .ZN(n6) );
  NOR2_X1 U8 ( .A1(n8), .A2(n1), .ZN(n13) );
  NOR2_X1 U9 ( .A1(n6), .A2(n7), .ZN(n23) );
  OAI21_X1 U10 ( .B1(MUX_SEL_C), .B2(n2), .A(n3), .ZN(n39) );
  NAND4_X1 U11 ( .A1(n4), .A2(n5), .A3(n6), .A4(n1), .ZN(n3) );
  NOR3_X1 U12 ( .A1(n1), .A2(n8), .A3(n9), .ZN(n2) );
  OAI21_X1 U13 ( .B1(MUX_SEL_D), .B2(n32), .A(n33), .ZN(n45) );
  NAND4_X1 U14 ( .A1(FSM_SEL[0]), .A2(n4), .A3(n5), .A4(n12), .ZN(n33) );
  NOR3_X1 U15 ( .A1(n12), .A2(n8), .A3(n19), .ZN(n32) );
  AOI21_X1 U16 ( .B1(MUX_SEL_A), .B2(BRANCH_TAKEN), .A(FSM_SEL[0]), .ZN(n29)
         );
  AOI21_X1 U17 ( .B1(MUX_SEL_D), .B2(BRANCH_TAKEN), .A(n8), .ZN(n37) );
  OAI21_X1 U18 ( .B1(MUX_SEL_A), .B2(n24), .A(n25), .ZN(n43) );
  NAND4_X1 U19 ( .A1(n16), .A2(n5), .A3(n6), .A4(n17), .ZN(n25) );
  NOR3_X1 U20 ( .A1(n17), .A2(n9), .A3(n18), .ZN(n24) );
  OAI21_X1 U21 ( .B1(MUX_SEL_B), .B2(n14), .A(n15), .ZN(n41) );
  NAND4_X1 U22 ( .A1(FSM_SEL[0]), .A2(n16), .A3(n5), .A4(n7), .ZN(n15) );
  NOR3_X1 U23 ( .A1(n7), .A2(n18), .A3(n19), .ZN(n14) );
  OAI21_X1 U25 ( .B1(n49), .B2(n10), .A(n11), .ZN(n40) );
  OAI211_X1 U26 ( .C1(n5), .C2(n26), .A(n6), .B(n13), .ZN(n11) );
  AOI211_X1 U28 ( .C1(n5), .C2(n26), .A(n8), .B(FSM_SEL[0]), .ZN(n10) );
  OAI21_X1 U29 ( .B1(n51), .B2(n27), .A(n28), .ZN(n44) );
  AOI211_X1 U30 ( .C1(n5), .C2(n34), .A(n18), .B(FSM_SEL[0]), .ZN(n27) );
  OAI21_X1 U32 ( .B1(n48), .B2(n35), .A(n36), .ZN(n47) );
  AOI211_X1 U33 ( .C1(n5), .C2(n30), .A(n6), .B(n8), .ZN(n35) );
  OAI21_X1 U34 ( .B1(n50), .B2(n20), .A(n21), .ZN(n42) );
  OAI211_X1 U35 ( .C1(n5), .C2(n22), .A(n16), .B(n23), .ZN(n21) );
  AOI211_X1 U36 ( .C1(n5), .C2(n22), .A(n6), .B(n18), .ZN(n20) );
  INV_X1 U37 ( .A(RST), .ZN(n38) );
endmodule


module CACHE_BPU_N32_SET_BIT2 ( ADDR, DATA_IN, DATA_OUT, ENC, RST, LOAD, CLK, 
        HIT_MISS );
  input [31:0] ADDR;
  input [31:0] DATA_IN;
  output [31:0] DATA_OUT;
  output [1:0] ENC;
  input RST, LOAD, CLK;
  output HIT_MISS;
  wire   VALID_BIT_1, VALID_BIT_2, VALID_BIT_3, VALID_BIT_4, COMP_OUT_1,
         COMP_OUT_2, COMP_OUT_3, COMP_OUT_4;
  wire   [31:0] IN_A_MUX;
  wire   [31:0] OUT_MUX;
  wire   [1:0] COUNT_OUT;
  wire   [31:0] CAM_OUT_1;
  wire   [31:0] CAM_OUT_2;
  wire   [31:0] CAM_OUT_3;
  wire   [31:0] CAM_OUT_4;
  wire   [3:0] IN_OR;
  wire   [1:0] IN_B_MUX_2;

  REG_N32_1 PC_REG ( .D(ADDR), .Q(IN_A_MUX), .EN(1'b1), .RST(RST), .CLK(CLK)
         );
  MUX21_GEN_N32_3 MUX_1 ( .A(IN_A_MUX), .B(ADDR), .SEL(LOAD), .Y(OUT_MUX) );
  CAM_BPU_N32_SET_BIT2 CAM_INST ( .ADDR(COUNT_OUT), .RST(RST), .WE(LOAD), 
        .DATA_IN(OUT_MUX), .ADDR_OUT_1(CAM_OUT_1), .ADDR_OUT_2(CAM_OUT_2), 
        .ADDR_OUT_3(CAM_OUT_3), .ADDR_OUT_4(CAM_OUT_4), .VALID_1(VALID_BIT_1), 
        .VALID_2(VALID_BIT_2), .VALID_3(VALID_BIT_3), .VALID_4(VALID_BIT_4) );
  EQU_COMPARATOR_N32_0 COMP_INST_1 ( .A(CAM_OUT_1), .B(OUT_MUX), .Y(COMP_OUT_1) );
  EQU_COMPARATOR_N32_4 COMP_INST_2 ( .A(CAM_OUT_2), .B(OUT_MUX), .Y(COMP_OUT_2) );
  EQU_COMPARATOR_N32_3 COMP_INST_3 ( .A(CAM_OUT_3), .B(OUT_MUX), .Y(COMP_OUT_3) );
  EQU_COMPARATOR_N32_2 COMP_INST_4 ( .A(CAM_OUT_4), .B(OUT_MUX), .Y(COMP_OUT_4) );
  AND_GATE_1_711 HIT_MISS_OUT_1 ( .A(COMP_OUT_1), .B(VALID_BIT_1), .Y(IN_OR[0]) );
  AND_GATE_1_710 HIT_MISS_OUT_2 ( .A(COMP_OUT_2), .B(VALID_BIT_2), .Y(IN_OR[1]) );
  AND_GATE_1_709 HIT_MISS_OUT_3 ( .A(COMP_OUT_3), .B(VALID_BIT_3), .Y(IN_OR[2]) );
  AND_GATE_1_708 HIT_MISS_OUT_4 ( .A(COMP_OUT_4), .B(VALID_BIT_4), .Y(IN_OR[3]) );
  N_OR_N4 HIT_MISS_OUT ( .A(IN_OR), .Y(HIT_MISS) );
  BPU_ENCODER ENCODER ( .A(IN_OR), .Y(IN_B_MUX_2) );
  SYNC_COUNTER_2BIT CNT_INST ( .EN(LOAD), .RST(RST), .CLK(CLK), .COUNT(
        COUNT_OUT) );
  MUX21_GEN_N2 MUX_2 ( .A(COUNT_OUT), .B(IN_B_MUX_2), .SEL(LOAD), .Y(ENC) );
  CACHE_DATA_BPU_N32_SET_BIT2 DATA_INST ( .DATA_IN(DATA_IN), .DATA_OUT(
        DATA_OUT), .ADDR(ENC), .CLK(CLK), .WE(LOAD) );
endmodule


module MUX21_GEN_N32_0 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   SB, n1, n2, n3, n4, n5, n6;
  wire   [31:0] Y1;
  wire   [31:0] Y2;

  INV_1_0 UIV ( .A(n1), .Y(SB) );
  NAND_GATE_0 UND1_0 ( .A(A[0]), .B(n1), .Y(Y1[0]) );
  NAND_GATE_1613 UND2_0 ( .A(B[0]), .B(n6), .Y(Y2[0]) );
  NAND_GATE_1612 UND3_0 ( .A(Y1[0]), .B(Y2[0]), .Y(Y[0]) );
  NAND_GATE_1611 UND1_1 ( .A(A[1]), .B(n3), .Y(Y1[1]) );
  NAND_GATE_1610 UND2_1 ( .A(B[1]), .B(n6), .Y(Y2[1]) );
  NAND_GATE_1609 UND3_1 ( .A(Y1[1]), .B(Y2[1]), .Y(Y[1]) );
  NAND_GATE_1608 UND1_2 ( .A(A[2]), .B(n3), .Y(Y1[2]) );
  NAND_GATE_1607 UND2_2 ( .A(B[2]), .B(n6), .Y(Y2[2]) );
  NAND_GATE_1606 UND3_2 ( .A(Y1[2]), .B(Y2[2]), .Y(Y[2]) );
  NAND_GATE_1605 UND1_3 ( .A(A[3]), .B(n3), .Y(Y1[3]) );
  NAND_GATE_1604 UND2_3 ( .A(B[3]), .B(n6), .Y(Y2[3]) );
  NAND_GATE_1603 UND3_3 ( .A(Y1[3]), .B(Y2[3]), .Y(Y[3]) );
  NAND_GATE_1602 UND1_4 ( .A(A[4]), .B(n3), .Y(Y1[4]) );
  NAND_GATE_1601 UND2_4 ( .A(B[4]), .B(n6), .Y(Y2[4]) );
  NAND_GATE_1600 UND3_4 ( .A(Y1[4]), .B(Y2[4]), .Y(Y[4]) );
  NAND_GATE_1599 UND1_5 ( .A(A[5]), .B(n3), .Y(Y1[5]) );
  NAND_GATE_1598 UND2_5 ( .A(B[5]), .B(n6), .Y(Y2[5]) );
  NAND_GATE_1597 UND3_5 ( .A(Y1[5]), .B(Y2[5]), .Y(Y[5]) );
  NAND_GATE_1596 UND1_6 ( .A(A[6]), .B(n3), .Y(Y1[6]) );
  NAND_GATE_1595 UND2_6 ( .A(B[6]), .B(n5), .Y(Y2[6]) );
  NAND_GATE_1594 UND3_6 ( .A(Y1[6]), .B(Y2[6]), .Y(Y[6]) );
  NAND_GATE_1593 UND1_7 ( .A(A[7]), .B(n3), .Y(Y1[7]) );
  NAND_GATE_1592 UND2_7 ( .A(B[7]), .B(n5), .Y(Y2[7]) );
  NAND_GATE_1591 UND3_7 ( .A(Y1[7]), .B(Y2[7]), .Y(Y[7]) );
  NAND_GATE_1590 UND1_8 ( .A(A[8]), .B(n2), .Y(Y1[8]) );
  NAND_GATE_1589 UND2_8 ( .A(B[8]), .B(n5), .Y(Y2[8]) );
  NAND_GATE_1588 UND3_8 ( .A(Y1[8]), .B(Y2[8]), .Y(Y[8]) );
  NAND_GATE_1587 UND1_9 ( .A(A[9]), .B(n2), .Y(Y1[9]) );
  NAND_GATE_1586 UND2_9 ( .A(B[9]), .B(n5), .Y(Y2[9]) );
  NAND_GATE_1585 UND3_9 ( .A(Y1[9]), .B(Y2[9]), .Y(Y[9]) );
  NAND_GATE_1584 UND1_10 ( .A(A[10]), .B(n2), .Y(Y1[10]) );
  NAND_GATE_1583 UND2_10 ( .A(B[10]), .B(n5), .Y(Y2[10]) );
  NAND_GATE_1582 UND3_10 ( .A(Y1[10]), .B(Y2[10]), .Y(Y[10]) );
  NAND_GATE_1581 UND1_11 ( .A(A[11]), .B(n2), .Y(Y1[11]) );
  NAND_GATE_1580 UND2_11 ( .A(B[11]), .B(n5), .Y(Y2[11]) );
  NAND_GATE_1579 UND3_11 ( .A(Y1[11]), .B(Y2[11]), .Y(Y[11]) );
  NAND_GATE_1578 UND1_12 ( .A(A[12]), .B(n2), .Y(Y1[12]) );
  NAND_GATE_1577 UND2_12 ( .A(B[12]), .B(n5), .Y(Y2[12]) );
  NAND_GATE_1576 UND3_12 ( .A(Y1[12]), .B(Y2[12]), .Y(Y[12]) );
  NAND_GATE_1575 UND1_13 ( .A(A[13]), .B(n2), .Y(Y1[13]) );
  NAND_GATE_1574 UND2_13 ( .A(B[13]), .B(n5), .Y(Y2[13]) );
  NAND_GATE_1573 UND3_13 ( .A(Y1[13]), .B(Y2[13]), .Y(Y[13]) );
  NAND_GATE_1572 UND1_14 ( .A(A[14]), .B(n2), .Y(Y1[14]) );
  NAND_GATE_1571 UND2_14 ( .A(B[14]), .B(n5), .Y(Y2[14]) );
  NAND_GATE_1570 UND3_14 ( .A(Y1[14]), .B(Y2[14]), .Y(Y[14]) );
  NAND_GATE_1569 UND1_15 ( .A(A[15]), .B(n2), .Y(Y1[15]) );
  NAND_GATE_1568 UND2_15 ( .A(B[15]), .B(n5), .Y(Y2[15]) );
  NAND_GATE_1567 UND3_15 ( .A(Y1[15]), .B(Y2[15]), .Y(Y[15]) );
  NAND_GATE_1566 UND1_16 ( .A(A[16]), .B(n2), .Y(Y1[16]) );
  NAND_GATE_1565 UND2_16 ( .A(B[16]), .B(n5), .Y(Y2[16]) );
  NAND_GATE_1564 UND3_16 ( .A(Y1[16]), .B(Y2[16]), .Y(Y[16]) );
  NAND_GATE_1563 UND1_17 ( .A(A[17]), .B(n2), .Y(Y1[17]) );
  NAND_GATE_1562 UND2_17 ( .A(B[17]), .B(n5), .Y(Y2[17]) );
  NAND_GATE_1561 UND3_17 ( .A(Y1[17]), .B(Y2[17]), .Y(Y[17]) );
  NAND_GATE_1560 UND1_18 ( .A(A[18]), .B(n2), .Y(Y1[18]) );
  NAND_GATE_1559 UND2_18 ( .A(B[18]), .B(n5), .Y(Y2[18]) );
  NAND_GATE_1558 UND3_18 ( .A(Y1[18]), .B(Y2[18]), .Y(Y[18]) );
  NAND_GATE_1557 UND1_19 ( .A(A[19]), .B(n2), .Y(Y1[19]) );
  NAND_GATE_1556 UND2_19 ( .A(B[19]), .B(n4), .Y(Y2[19]) );
  NAND_GATE_1555 UND3_19 ( .A(Y1[19]), .B(Y2[19]), .Y(Y[19]) );
  NAND_GATE_1554 UND1_20 ( .A(A[20]), .B(n2), .Y(Y1[20]) );
  NAND_GATE_1553 UND2_20 ( .A(B[20]), .B(n4), .Y(Y2[20]) );
  NAND_GATE_1552 UND3_20 ( .A(Y1[20]), .B(Y2[20]), .Y(Y[20]) );
  NAND_GATE_1551 UND1_21 ( .A(A[21]), .B(n1), .Y(Y1[21]) );
  NAND_GATE_1550 UND2_21 ( .A(B[21]), .B(n4), .Y(Y2[21]) );
  NAND_GATE_1549 UND3_21 ( .A(Y1[21]), .B(Y2[21]), .Y(Y[21]) );
  NAND_GATE_1548 UND1_22 ( .A(A[22]), .B(n1), .Y(Y1[22]) );
  NAND_GATE_1547 UND2_22 ( .A(B[22]), .B(n4), .Y(Y2[22]) );
  NAND_GATE_1546 UND3_22 ( .A(Y1[22]), .B(Y2[22]), .Y(Y[22]) );
  NAND_GATE_1545 UND1_23 ( .A(A[23]), .B(n1), .Y(Y1[23]) );
  NAND_GATE_1544 UND2_23 ( .A(B[23]), .B(n4), .Y(Y2[23]) );
  NAND_GATE_1543 UND3_23 ( .A(Y1[23]), .B(Y2[23]), .Y(Y[23]) );
  NAND_GATE_1542 UND1_24 ( .A(A[24]), .B(n1), .Y(Y1[24]) );
  NAND_GATE_1541 UND2_24 ( .A(B[24]), .B(n4), .Y(Y2[24]) );
  NAND_GATE_1540 UND3_24 ( .A(Y1[24]), .B(Y2[24]), .Y(Y[24]) );
  NAND_GATE_1539 UND1_25 ( .A(A[25]), .B(n1), .Y(Y1[25]) );
  NAND_GATE_1538 UND2_25 ( .A(B[25]), .B(n4), .Y(Y2[25]) );
  NAND_GATE_1537 UND3_25 ( .A(Y1[25]), .B(Y2[25]), .Y(Y[25]) );
  NAND_GATE_1536 UND1_26 ( .A(A[26]), .B(n1), .Y(Y1[26]) );
  NAND_GATE_1535 UND2_26 ( .A(B[26]), .B(n4), .Y(Y2[26]) );
  NAND_GATE_1534 UND3_26 ( .A(Y1[26]), .B(Y2[26]), .Y(Y[26]) );
  NAND_GATE_1533 UND1_27 ( .A(A[27]), .B(n1), .Y(Y1[27]) );
  NAND_GATE_1532 UND2_27 ( .A(B[27]), .B(n4), .Y(Y2[27]) );
  NAND_GATE_1531 UND3_27 ( .A(Y1[27]), .B(Y2[27]), .Y(Y[27]) );
  NAND_GATE_1530 UND1_28 ( .A(A[28]), .B(n1), .Y(Y1[28]) );
  NAND_GATE_1529 UND2_28 ( .A(B[28]), .B(n4), .Y(Y2[28]) );
  NAND_GATE_1528 UND3_28 ( .A(Y1[28]), .B(Y2[28]), .Y(Y[28]) );
  NAND_GATE_1527 UND1_29 ( .A(A[29]), .B(n1), .Y(Y1[29]) );
  NAND_GATE_1526 UND2_29 ( .A(B[29]), .B(n4), .Y(Y2[29]) );
  NAND_GATE_1525 UND3_29 ( .A(Y1[29]), .B(Y2[29]), .Y(Y[29]) );
  NAND_GATE_1524 UND1_30 ( .A(A[30]), .B(n1), .Y(Y1[30]) );
  NAND_GATE_1523 UND2_30 ( .A(B[30]), .B(n4), .Y(Y2[30]) );
  NAND_GATE_1522 UND3_30 ( .A(Y1[30]), .B(Y2[30]), .Y(Y[30]) );
  NAND_GATE_1521 UND1_31 ( .A(A[31]), .B(n1), .Y(Y1[31]) );
  NAND_GATE_1520 UND2_31 ( .A(B[31]), .B(n4), .Y(Y2[31]) );
  NAND_GATE_1519 UND3_31 ( .A(Y1[31]), .B(Y2[31]), .Y(Y[31]) );
  BUF_X1 U1 ( .A(SB), .Z(n4) );
  BUF_X1 U2 ( .A(SB), .Z(n5) );
  BUF_X1 U3 ( .A(SB), .Z(n6) );
  BUF_X1 U4 ( .A(SEL), .Z(n3) );
  BUF_X1 U5 ( .A(SEL), .Z(n1) );
  BUF_X1 U6 ( .A(SEL), .Z(n2) );
endmodule


module RCA_GEN_NO_C_N30 ( A, B, S, Co );
  input [29:0] A;
  input [29:0] B;
  output [29:0] S;
  output Co;

  wire   [28:0] CTMP;

  HA_0 HA_INST ( .A(A[0]), .B(B[0]), .S(S[0]), .Co(CTMP[0]) );
  FA_0 FAI_0 ( .A(A[1]), .B(B[1]), .Ci(CTMP[0]), .S(S[1]), .Co(CTMP[1]) );
  FA_297 FAI_1 ( .A(A[2]), .B(B[2]), .Ci(CTMP[1]), .S(S[2]), .Co(CTMP[2]) );
  FA_296 FAI_2 ( .A(A[3]), .B(B[3]), .Ci(CTMP[2]), .S(S[3]), .Co(CTMP[3]) );
  FA_295 FAI_3 ( .A(A[4]), .B(B[4]), .Ci(CTMP[3]), .S(S[4]), .Co(CTMP[4]) );
  FA_294 FAI_4 ( .A(A[5]), .B(B[5]), .Ci(CTMP[4]), .S(S[5]), .Co(CTMP[5]) );
  FA_293 FAI_5 ( .A(A[6]), .B(B[6]), .Ci(CTMP[5]), .S(S[6]), .Co(CTMP[6]) );
  FA_292 FAI_6 ( .A(A[7]), .B(B[7]), .Ci(CTMP[6]), .S(S[7]), .Co(CTMP[7]) );
  FA_291 FAI_7 ( .A(A[8]), .B(B[8]), .Ci(CTMP[7]), .S(S[8]), .Co(CTMP[8]) );
  FA_290 FAI_8 ( .A(A[9]), .B(B[9]), .Ci(CTMP[8]), .S(S[9]), .Co(CTMP[9]) );
  FA_289 FAI_9 ( .A(A[10]), .B(B[10]), .Ci(CTMP[9]), .S(S[10]), .Co(CTMP[10])
         );
  FA_288 FAI_10 ( .A(A[11]), .B(B[11]), .Ci(CTMP[10]), .S(S[11]), .Co(CTMP[11]) );
  FA_287 FAI_11 ( .A(A[12]), .B(B[12]), .Ci(CTMP[11]), .S(S[12]), .Co(CTMP[12]) );
  FA_286 FAI_12 ( .A(A[13]), .B(B[13]), .Ci(CTMP[12]), .S(S[13]), .Co(CTMP[13]) );
  FA_285 FAI_13 ( .A(A[14]), .B(B[14]), .Ci(CTMP[13]), .S(S[14]), .Co(CTMP[14]) );
  FA_284 FAI_14 ( .A(A[15]), .B(B[15]), .Ci(CTMP[14]), .S(S[15]), .Co(CTMP[15]) );
  FA_283 FAI_15 ( .A(A[16]), .B(B[16]), .Ci(CTMP[15]), .S(S[16]), .Co(CTMP[16]) );
  FA_282 FAI_16 ( .A(A[17]), .B(B[17]), .Ci(CTMP[16]), .S(S[17]), .Co(CTMP[17]) );
  FA_281 FAI_17 ( .A(A[18]), .B(B[18]), .Ci(CTMP[17]), .S(S[18]), .Co(CTMP[18]) );
  FA_280 FAI_18 ( .A(A[19]), .B(B[19]), .Ci(CTMP[18]), .S(S[19]), .Co(CTMP[19]) );
  FA_279 FAI_19 ( .A(A[20]), .B(B[20]), .Ci(CTMP[19]), .S(S[20]), .Co(CTMP[20]) );
  FA_278 FAI_20 ( .A(A[21]), .B(B[21]), .Ci(CTMP[20]), .S(S[21]), .Co(CTMP[21]) );
  FA_277 FAI_21 ( .A(A[22]), .B(B[22]), .Ci(CTMP[21]), .S(S[22]), .Co(CTMP[22]) );
  FA_276 FAI_22 ( .A(A[23]), .B(B[23]), .Ci(CTMP[22]), .S(S[23]), .Co(CTMP[23]) );
  FA_275 FAI_23 ( .A(A[24]), .B(B[24]), .Ci(CTMP[23]), .S(S[24]), .Co(CTMP[24]) );
  FA_274 FAI_24 ( .A(A[25]), .B(B[25]), .Ci(CTMP[24]), .S(S[25]), .Co(CTMP[25]) );
  FA_273 FAI_25 ( .A(A[26]), .B(B[26]), .Ci(CTMP[25]), .S(S[26]), .Co(CTMP[26]) );
  FA_272 FAI_26 ( .A(A[27]), .B(B[27]), .Ci(CTMP[26]), .S(S[27]), .Co(CTMP[27]) );
  FA_271 FAI_27 ( .A(A[28]), .B(B[28]), .Ci(CTMP[27]), .S(S[28]), .Co(CTMP[28]) );
  FA_270 FAI_28 ( .A(A[29]), .B(B[29]), .Ci(CTMP[28]), .S(S[29]), .Co(Co) );
endmodule


module CACHE_N32_TAG_BIT23_SET_BIT4_N_DATA5 ( ADDR, ADDR_OUT, DATA_IN, 
        DATA_OUT, RST, LOAD, CLK, HIT_MISS );
  input [31:0] ADDR;
  output [31:0] ADDR_OUT;
  input [7:0] DATA_IN;
  output [31:0] DATA_OUT;
  input RST, LOAD, CLK;
  output HIT_MISS;
  wire   \ADDR[31] , \ADDR[30] , \ADDR[29] , \ADDR[28] , \ADDR[27] ,
         \ADDR[26] , \ADDR[25] , \ADDR[24] , \ADDR[23] , \ADDR[22] ,
         \ADDR[21] , \ADDR[20] , \ADDR[19] , \ADDR[18] , \ADDR[17] ,
         \ADDR[16] , \ADDR[15] , \ADDR[14] , \ADDR[13] , \ADDR[12] ,
         \ADDR[11] , \ADDR[10] , \ADDR[9] , \ADDR[8] , \ADDR[7] , \ADDR[6] ,
         \ADDR[5] , VALID_BIT, COMP_OUT, CNT_RST, n1, n2;
  wire   [4:0] OFF_DATA;
  wire   [22:0] IN_COMP;
  assign ADDR_OUT[31] = \ADDR[31] ;
  assign \ADDR[31]  = ADDR[31];
  assign ADDR_OUT[30] = \ADDR[30] ;
  assign \ADDR[30]  = ADDR[30];
  assign ADDR_OUT[29] = \ADDR[29] ;
  assign \ADDR[29]  = ADDR[29];
  assign ADDR_OUT[28] = \ADDR[28] ;
  assign \ADDR[28]  = ADDR[28];
  assign ADDR_OUT[27] = \ADDR[27] ;
  assign \ADDR[27]  = ADDR[27];
  assign ADDR_OUT[26] = \ADDR[26] ;
  assign \ADDR[26]  = ADDR[26];
  assign ADDR_OUT[25] = \ADDR[25] ;
  assign \ADDR[25]  = ADDR[25];
  assign ADDR_OUT[24] = \ADDR[24] ;
  assign \ADDR[24]  = ADDR[24];
  assign ADDR_OUT[23] = \ADDR[23] ;
  assign \ADDR[23]  = ADDR[23];
  assign ADDR_OUT[22] = \ADDR[22] ;
  assign \ADDR[22]  = ADDR[22];
  assign ADDR_OUT[21] = \ADDR[21] ;
  assign \ADDR[21]  = ADDR[21];
  assign ADDR_OUT[20] = \ADDR[20] ;
  assign \ADDR[20]  = ADDR[20];
  assign ADDR_OUT[19] = \ADDR[19] ;
  assign \ADDR[19]  = ADDR[19];
  assign ADDR_OUT[18] = \ADDR[18] ;
  assign \ADDR[18]  = ADDR[18];
  assign ADDR_OUT[17] = \ADDR[17] ;
  assign \ADDR[17]  = ADDR[17];
  assign ADDR_OUT[16] = \ADDR[16] ;
  assign \ADDR[16]  = ADDR[16];
  assign ADDR_OUT[15] = \ADDR[15] ;
  assign \ADDR[15]  = ADDR[15];
  assign ADDR_OUT[14] = \ADDR[14] ;
  assign \ADDR[14]  = ADDR[14];
  assign ADDR_OUT[13] = \ADDR[13] ;
  assign \ADDR[13]  = ADDR[13];
  assign ADDR_OUT[12] = \ADDR[12] ;
  assign \ADDR[12]  = ADDR[12];
  assign ADDR_OUT[11] = \ADDR[11] ;
  assign \ADDR[11]  = ADDR[11];
  assign ADDR_OUT[10] = \ADDR[10] ;
  assign \ADDR[10]  = ADDR[10];
  assign ADDR_OUT[9] = \ADDR[9] ;
  assign \ADDR[9]  = ADDR[9];
  assign ADDR_OUT[8] = \ADDR[8] ;
  assign \ADDR[8]  = ADDR[8];
  assign ADDR_OUT[7] = \ADDR[7] ;
  assign \ADDR[7]  = ADDR[7];
  assign ADDR_OUT[6] = \ADDR[6] ;
  assign \ADDR[6]  = ADDR[6];
  assign ADDR_OUT[5] = \ADDR[5] ;
  assign \ADDR[5]  = ADDR[5];

  NAND2_X1 U2 ( .A1(n2), .A2(n1), .ZN(CNT_RST) );
  MUX21_GEN_N5 MUX_1 ( .A(ADDR_OUT[4:0]), .B(ADDR[4:0]), .SEL(n2), .Y(OFF_DATA) );
  CAM_TAG_BIT23_SET_BIT4 CAM_INST ( .TAG_IN({\ADDR[31] , \ADDR[30] , 
        \ADDR[29] , \ADDR[28] , \ADDR[27] , \ADDR[26] , \ADDR[25] , \ADDR[24] , 
        \ADDR[23] , \ADDR[22] , \ADDR[21] , \ADDR[20] , \ADDR[19] , \ADDR[18] , 
        \ADDR[17] , \ADDR[16] , \ADDR[15] , \ADDR[14] , \ADDR[13] , \ADDR[12] , 
        \ADDR[11] , \ADDR[10] , \ADDR[9] }), .TAG_OUT(IN_COMP), .SET_INDEX({
        \ADDR[8] , \ADDR[7] , \ADDR[6] , \ADDR[5] }), .COUNT(ADDR_OUT[4:0]), 
        .VALID(VALID_BIT), .CLK(CLK), .RST(RST), .WE(n2) );
  CACHE_DATA_N32_N_DATA5_SET_BIT4 DATA_INST ( .DATA_IN(DATA_IN), .DATA_OUT(
        DATA_OUT), .ADDR({\ADDR[8] , \ADDR[7] , \ADDR[6] , \ADDR[5] }), 
        .OFFSET(OFF_DATA), .CLK(CLK), .WE(n2) );
  EQU_COMPARATOR_N23 COMP_INST ( .A(IN_COMP), .B({\ADDR[31] , \ADDR[30] , 
        \ADDR[29] , \ADDR[28] , \ADDR[27] , \ADDR[26] , \ADDR[25] , \ADDR[24] , 
        \ADDR[23] , \ADDR[22] , \ADDR[21] , \ADDR[20] , \ADDR[19] , \ADDR[18] , 
        \ADDR[17] , \ADDR[16] , \ADDR[15] , \ADDR[14] , \ADDR[13] , \ADDR[12] , 
        \ADDR[11] , \ADDR[10] , \ADDR[9] }), .Y(COMP_OUT) );
  SYNC_COUNTER_5BIT CNT_INST ( .EN(n2), .RST(CNT_RST), .CLK(CLK), .COUNT(
        ADDR_OUT[4:0]) );
  AND_GATE_339 HIT_MISS_OUT ( .A(COMP_OUT), .B(VALID_BIT), .Y(HIT_MISS) );
  BUF_X1 U1 ( .A(LOAD), .Z(n2) );
  INV_X1 U3 ( .A(RST), .ZN(n1) );
endmodule


module FORWARD_UNIT_OPCODE_SIZE6_N_ADDR5 ( CLK, RST, OPCODE_IF, REG_A_IF, 
        OPCODE_ID, REG_DEST_ID, REG_DEST_EXE, REG_DEST_MEM, REG_A, REG_B, 
        MUX_A, MUX_B, MUX_C, MUX_D, RST_DIV, STALL_BRANCH, STALL );
  input [5:0] OPCODE_IF;
  input [4:0] REG_A_IF;
  input [5:0] OPCODE_ID;
  input [4:0] REG_DEST_ID;
  input [4:0] REG_DEST_EXE;
  input [4:0] REG_DEST_MEM;
  input [4:0] REG_A;
  input [4:0] REG_B;
  output [1:0] MUX_A;
  output [1:0] MUX_B;
  output [1:0] MUX_C;
  output [1:0] MUX_D;
  input CLK, RST;
  output RST_DIV, STALL_BRANCH, STALL;
  wire   EN_REG, CMP_A_EXE, CMP_A_MEM, CMP_B_EXE, CMP_B_MEM, CMP_BRANCH_ID,
         CMP_BRANCH_EXE, CMP_BRANCH_MEM, CMP_C_EXE, CMP_C_MEM, n1;
  wire   [5:0] OPCODE_EXE;
  wire   [5:0] OPCODE_MEM;
  wire   [5:0] OPCODE_WB;

  EQU_COMPARATOR_N5_0 CMP_EXE_A ( .A(REG_A), .B(REG_DEST_EXE), .Y(CMP_A_EXE)
         );
  EQU_COMPARATOR_N5_6 CMP_MEM_A ( .A(REG_A), .B(REG_DEST_MEM), .Y(CMP_A_MEM)
         );
  EQU_COMPARATOR_N5_5 CMP_EXE_B ( .A(REG_B), .B(REG_DEST_EXE), .Y(CMP_B_EXE)
         );
  EQU_COMPARATOR_N5_4 CMP_MEM_B ( .A(REG_B), .B(REG_DEST_MEM), .Y(CMP_B_MEM)
         );
  EQU_COMPARATOR_N5_3 CMP_ID_IF ( .A(REG_A_IF), .B(REG_DEST_ID), .Y(
        CMP_BRANCH_ID) );
  EQU_COMPARATOR_N5_2 CMP_ID_EXE ( .A(REG_A_IF), .B(REG_DEST_EXE), .Y(
        CMP_BRANCH_EXE) );
  EQU_COMPARATOR_N5_1 CMP_ID_MEM ( .A(REG_A_IF), .B(REG_DEST_MEM), .Y(
        CMP_BRANCH_MEM) );
  REG_N6_0 OP_PIPE_ID_EXE ( .D(OPCODE_ID), .Q(OPCODE_EXE), .EN(EN_REG), .RST(
        n1), .CLK(CLK) );
  REG_N6_2 OP_PIPE_EXE_MEM ( .D(OPCODE_EXE), .Q(OPCODE_MEM), .EN(EN_REG), 
        .RST(n1), .CLK(CLK) );
  REG_N6_1 OP_PIPE_MEM_WB ( .D(OPCODE_MEM), .Q(OPCODE_WB), .EN(1'b1), .RST(n1), 
        .CLK(CLK) );
  FD_1_149 CMP_PIPE_C_EXE ( .D(CMP_B_EXE), .CLK(CLK), .EN(EN_REG), .RST(n1), 
        .Q(CMP_C_EXE) );
  FD_1_148 CMP_PIPE_C_MEM ( .D(CMP_B_MEM), .CLK(CLK), .EN(EN_REG), .RST(n1), 
        .Q(CMP_C_MEM) );
  FORW_FSM_OPCODE_SIZE6_N_ADDR5 FSM_FORWARD ( .CLK(CLK), .RST(n1), .CMP_A_EXE(
        CMP_A_EXE), .CMP_A_MEM(CMP_A_MEM), .CMP_B_EXE(CMP_B_EXE), .CMP_B_MEM(
        CMP_B_MEM), .CMP_C_EXE(CMP_C_EXE), .CMP_C_MEM(CMP_C_MEM), 
        .CMP_BRANCH_ID(CMP_BRANCH_ID), .CMP_BRANCH_EXE(CMP_BRANCH_EXE), 
        .CMP_BRANCH_MEM(CMP_BRANCH_MEM), .OPCODE_IF(OPCODE_IF), .OPCODE_ID(
        OPCODE_ID), .OPCODE_EXE(OPCODE_EXE), .OPCODE_MEM(OPCODE_MEM), 
        .OPCODE_WB(OPCODE_WB), .MUX_A(MUX_A), .MUX_B(MUX_B), .MUX_C(MUX_C), 
        .MUX_D(MUX_D), .RST_DIV(RST_DIV), .STALL_BRANCH(STALL_BRANCH), .STALL(
        STALL) );
  BUF_X1 U2 ( .A(RST), .Z(n1) );
  INV_X1 U3 ( .A(STALL), .ZN(EN_REG) );
endmodule


module WB_N32_N_ADDR5 ( IN_MEM, IN_ALU, IN_NPC, SEL, DEST_REG_IN, DEST_REG_OUT, 
        OUT_WB );
  input [31:0] IN_MEM;
  input [31:0] IN_ALU;
  input [31:0] IN_NPC;
  input [1:0] SEL;
  input [4:0] DEST_REG_IN;
  output [4:0] DEST_REG_OUT;
  output [31:0] OUT_WB;

  assign DEST_REG_OUT[4] = DEST_REG_IN[4];
  assign DEST_REG_OUT[3] = DEST_REG_IN[3];
  assign DEST_REG_OUT[2] = DEST_REG_IN[2];
  assign DEST_REG_OUT[1] = DEST_REG_IN[1];
  assign DEST_REG_OUT[0] = DEST_REG_IN[0];

  MUX41_GEN_N32_1 MUX_INST ( .A(IN_MEM), .B(IN_ALU), .C(IN_NPC), .D({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL(SEL), .Y(OUT_WB) );
endmodule


module MEMORY_N32_N_ADDR5 ( IN_ALU, DEST_REG_IN, REG_B_IN, FORW_ALU_WB, 
        FORW_MEM_WB, FORW_REG, SEL_DATA, RESET, ENABLE, DATA_IN_MEM, LOAD_TYPE, 
        STORE_MASK, ADDR_MEM, DATA_OUT_MEM, DEST_REG_OUT, MEMORY_OUT, OUT_ALU
 );
  input [31:0] IN_ALU;
  input [4:0] DEST_REG_IN;
  input [31:0] REG_B_IN;
  input [31:0] FORW_ALU_WB;
  input [31:0] FORW_MEM_WB;
  input [31:0] FORW_REG;
  input [1:0] SEL_DATA;
  input [31:0] DATA_IN_MEM;
  input [2:0] LOAD_TYPE;
  input [1:0] STORE_MASK;
  output [31:0] ADDR_MEM;
  output [31:0] DATA_OUT_MEM;
  output [4:0] DEST_REG_OUT;
  output [31:0] MEMORY_OUT;
  output [31:0] OUT_ALU;
  input RESET, ENABLE;
  wire   n1, n2, n3;
  wire   [31:8] OUT_MUX;
  assign ADDR_MEM[31] = IN_ALU[31];
  assign OUT_ALU[31] = IN_ALU[31];
  assign ADDR_MEM[30] = IN_ALU[30];
  assign OUT_ALU[30] = IN_ALU[30];
  assign ADDR_MEM[29] = IN_ALU[29];
  assign OUT_ALU[29] = IN_ALU[29];
  assign ADDR_MEM[28] = IN_ALU[28];
  assign OUT_ALU[28] = IN_ALU[28];
  assign ADDR_MEM[27] = IN_ALU[27];
  assign OUT_ALU[27] = IN_ALU[27];
  assign ADDR_MEM[26] = IN_ALU[26];
  assign OUT_ALU[26] = IN_ALU[26];
  assign ADDR_MEM[25] = IN_ALU[25];
  assign OUT_ALU[25] = IN_ALU[25];
  assign ADDR_MEM[24] = IN_ALU[24];
  assign OUT_ALU[24] = IN_ALU[24];
  assign ADDR_MEM[23] = IN_ALU[23];
  assign OUT_ALU[23] = IN_ALU[23];
  assign ADDR_MEM[22] = IN_ALU[22];
  assign OUT_ALU[22] = IN_ALU[22];
  assign ADDR_MEM[21] = IN_ALU[21];
  assign OUT_ALU[21] = IN_ALU[21];
  assign ADDR_MEM[20] = IN_ALU[20];
  assign OUT_ALU[20] = IN_ALU[20];
  assign ADDR_MEM[19] = IN_ALU[19];
  assign OUT_ALU[19] = IN_ALU[19];
  assign ADDR_MEM[18] = IN_ALU[18];
  assign OUT_ALU[18] = IN_ALU[18];
  assign ADDR_MEM[17] = IN_ALU[17];
  assign OUT_ALU[17] = IN_ALU[17];
  assign ADDR_MEM[16] = IN_ALU[16];
  assign OUT_ALU[16] = IN_ALU[16];
  assign ADDR_MEM[15] = IN_ALU[15];
  assign OUT_ALU[15] = IN_ALU[15];
  assign ADDR_MEM[14] = IN_ALU[14];
  assign OUT_ALU[14] = IN_ALU[14];
  assign ADDR_MEM[13] = IN_ALU[13];
  assign OUT_ALU[13] = IN_ALU[13];
  assign ADDR_MEM[12] = IN_ALU[12];
  assign OUT_ALU[12] = IN_ALU[12];
  assign ADDR_MEM[11] = IN_ALU[11];
  assign OUT_ALU[11] = IN_ALU[11];
  assign ADDR_MEM[10] = IN_ALU[10];
  assign OUT_ALU[10] = IN_ALU[10];
  assign ADDR_MEM[9] = IN_ALU[9];
  assign OUT_ALU[9] = IN_ALU[9];
  assign ADDR_MEM[8] = IN_ALU[8];
  assign OUT_ALU[8] = IN_ALU[8];
  assign ADDR_MEM[7] = IN_ALU[7];
  assign OUT_ALU[7] = IN_ALU[7];
  assign ADDR_MEM[6] = IN_ALU[6];
  assign OUT_ALU[6] = IN_ALU[6];
  assign ADDR_MEM[5] = IN_ALU[5];
  assign OUT_ALU[5] = IN_ALU[5];
  assign ADDR_MEM[4] = IN_ALU[4];
  assign OUT_ALU[4] = IN_ALU[4];
  assign ADDR_MEM[3] = IN_ALU[3];
  assign OUT_ALU[3] = IN_ALU[3];
  assign ADDR_MEM[2] = IN_ALU[2];
  assign OUT_ALU[2] = IN_ALU[2];
  assign ADDR_MEM[1] = IN_ALU[1];
  assign OUT_ALU[1] = IN_ALU[1];
  assign ADDR_MEM[0] = IN_ALU[0];
  assign OUT_ALU[0] = IN_ALU[0];
  assign DEST_REG_OUT[4] = DEST_REG_IN[4];
  assign DEST_REG_OUT[3] = DEST_REG_IN[3];
  assign DEST_REG_OUT[2] = DEST_REG_IN[2];
  assign DEST_REG_OUT[1] = DEST_REG_IN[1];
  assign DEST_REG_OUT[0] = DEST_REG_IN[0];

  AND_GATE_1_735 SH_MASK_0 ( .A(OUT_MUX[31]), .B(STORE_MASK[0]), .Y(
        DATA_OUT_MEM[31]) );
  AND_GATE_1_734 SH_MASK_1 ( .A(OUT_MUX[30]), .B(STORE_MASK[0]), .Y(
        DATA_OUT_MEM[30]) );
  AND_GATE_1_733 SH_MASK_2 ( .A(OUT_MUX[29]), .B(STORE_MASK[0]), .Y(
        DATA_OUT_MEM[29]) );
  AND_GATE_1_732 SH_MASK_3 ( .A(OUT_MUX[28]), .B(STORE_MASK[0]), .Y(
        DATA_OUT_MEM[28]) );
  AND_GATE_1_731 SH_MASK_4 ( .A(OUT_MUX[27]), .B(STORE_MASK[0]), .Y(
        DATA_OUT_MEM[27]) );
  AND_GATE_1_730 SH_MASK_5 ( .A(OUT_MUX[26]), .B(STORE_MASK[0]), .Y(
        DATA_OUT_MEM[26]) );
  AND_GATE_1_729 SH_MASK_6 ( .A(OUT_MUX[25]), .B(STORE_MASK[0]), .Y(
        DATA_OUT_MEM[25]) );
  AND_GATE_1_728 SH_MASK_7 ( .A(OUT_MUX[24]), .B(STORE_MASK[0]), .Y(
        DATA_OUT_MEM[24]) );
  AND_GATE_1_727 SH_MASK_8 ( .A(OUT_MUX[23]), .B(STORE_MASK[0]), .Y(
        DATA_OUT_MEM[23]) );
  AND_GATE_1_726 SH_MASK_9 ( .A(OUT_MUX[22]), .B(STORE_MASK[0]), .Y(
        DATA_OUT_MEM[22]) );
  AND_GATE_1_725 SH_MASK_10 ( .A(OUT_MUX[21]), .B(STORE_MASK[0]), .Y(
        DATA_OUT_MEM[21]) );
  AND_GATE_1_724 SH_MASK_11 ( .A(OUT_MUX[20]), .B(STORE_MASK[0]), .Y(
        DATA_OUT_MEM[20]) );
  AND_GATE_1_723 SH_MASK_12 ( .A(OUT_MUX[19]), .B(STORE_MASK[0]), .Y(
        DATA_OUT_MEM[19]) );
  AND_GATE_1_722 SH_MASK_13 ( .A(OUT_MUX[18]), .B(STORE_MASK[0]), .Y(
        DATA_OUT_MEM[18]) );
  AND_GATE_1_721 SH_MASK_14 ( .A(OUT_MUX[17]), .B(STORE_MASK[0]), .Y(
        DATA_OUT_MEM[17]) );
  AND_GATE_1_720 SH_MASK_15 ( .A(OUT_MUX[16]), .B(STORE_MASK[0]), .Y(
        DATA_OUT_MEM[16]) );
  AND_GATE_1_719 SB_MASK_16 ( .A(OUT_MUX[15]), .B(STORE_MASK[1]), .Y(
        DATA_OUT_MEM[15]) );
  AND_GATE_1_718 SB_MASK_17 ( .A(OUT_MUX[14]), .B(STORE_MASK[1]), .Y(
        DATA_OUT_MEM[14]) );
  AND_GATE_1_717 SB_MASK_18 ( .A(OUT_MUX[13]), .B(STORE_MASK[1]), .Y(
        DATA_OUT_MEM[13]) );
  AND_GATE_1_716 SB_MASK_19 ( .A(OUT_MUX[12]), .B(STORE_MASK[1]), .Y(
        DATA_OUT_MEM[12]) );
  AND_GATE_1_715 SB_MASK_20 ( .A(OUT_MUX[11]), .B(STORE_MASK[1]), .Y(
        DATA_OUT_MEM[11]) );
  AND_GATE_1_714 SB_MASK_21 ( .A(OUT_MUX[10]), .B(STORE_MASK[1]), .Y(
        DATA_OUT_MEM[10]) );
  AND_GATE_1_713 SB_MASK_22 ( .A(OUT_MUX[9]), .B(STORE_MASK[1]), .Y(
        DATA_OUT_MEM[9]) );
  AND_GATE_1_712 SB_MASK_23 ( .A(OUT_MUX[8]), .B(STORE_MASK[1]), .Y(
        DATA_OUT_MEM[8]) );
  MUX41_GEN_N32_2 REGB_MUX ( .A(REG_B_IN), .B(FORW_ALU_WB), .C(FORW_MEM_WB), 
        .D(FORW_REG), .SEL(SEL_DATA), .Y({OUT_MUX, DATA_OUT_MEM[7:0]}) );
  MUX51_GEN_N32_1 LOAD_MUX ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n3, DATA_IN_MEM[6:0]}), .B({n1, n1, n1, 
        n1, n1, n2, n1, n1, n1, n1, n1, n1, n2, n2, n2, n2, n2, n2, n2, n2, n2, 
        n2, n2, n2, n3, DATA_IN_MEM[6:0]}), .C({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        DATA_IN_MEM[15:8], n1, DATA_IN_MEM[6:0]}), .D({DATA_IN_MEM[15], 
        DATA_IN_MEM[15], DATA_IN_MEM[15], DATA_IN_MEM[15], DATA_IN_MEM[15], 
        DATA_IN_MEM[15], DATA_IN_MEM[15], DATA_IN_MEM[15], DATA_IN_MEM[15], 
        DATA_IN_MEM[15], DATA_IN_MEM[15], DATA_IN_MEM[15], DATA_IN_MEM[15], 
        DATA_IN_MEM[15], DATA_IN_MEM[15], DATA_IN_MEM[15], DATA_IN_MEM[15:8], 
        n3, DATA_IN_MEM[6:0]}), .E({DATA_IN_MEM[31:8], n1, DATA_IN_MEM[6:0]}), 
        .SEL(LOAD_TYPE), .Y(MEMORY_OUT) );
  BUF_X1 U2 ( .A(DATA_IN_MEM[7]), .Z(n3) );
  BUF_X1 U3 ( .A(DATA_IN_MEM[7]), .Z(n1) );
  BUF_X1 U4 ( .A(DATA_IN_MEM[7]), .Z(n2) );
endmodule


module EXECUTE_N32_N_ADDR5_ALUSIZE5 ( REG_A, REG_B, IMMEDIATE, FORW_ALU_MEM, 
        FORW_ALU_WB, FORW_MEM_WB, DEST_REG_IN, ALU_CODE, OP_SEL_A, OP_SEL_B, 
        CLK, RST, DEST_REG_OUT, OUTPUT_ALU, RST_DIV, REG_B_OUT );
  input [31:0] REG_A;
  input [31:0] REG_B;
  input [31:0] IMMEDIATE;
  input [31:0] FORW_ALU_MEM;
  input [31:0] FORW_ALU_WB;
  input [31:0] FORW_MEM_WB;
  input [4:0] DEST_REG_IN;
  input [4:0] ALU_CODE;
  input [1:0] OP_SEL_A;
  input [2:0] OP_SEL_B;
  output [4:0] DEST_REG_OUT;
  output [31:0] OUTPUT_ALU;
  output [31:0] REG_B_OUT;
  input CLK, RST, RST_DIV;

  wire   [31:0] IN_A_ALU_SIG;
  wire   [31:0] IN_B_ALU_SIG;
  assign DEST_REG_OUT[4] = DEST_REG_IN[4];
  assign DEST_REG_OUT[3] = DEST_REG_IN[3];
  assign DEST_REG_OUT[2] = DEST_REG_IN[2];
  assign DEST_REG_OUT[1] = DEST_REG_IN[1];
  assign DEST_REG_OUT[0] = DEST_REG_IN[0];
  assign REG_B_OUT[31] = REG_B[31];
  assign REG_B_OUT[30] = REG_B[30];
  assign REG_B_OUT[29] = REG_B[29];
  assign REG_B_OUT[28] = REG_B[28];
  assign REG_B_OUT[27] = REG_B[27];
  assign REG_B_OUT[26] = REG_B[26];
  assign REG_B_OUT[25] = REG_B[25];
  assign REG_B_OUT[24] = REG_B[24];
  assign REG_B_OUT[23] = REG_B[23];
  assign REG_B_OUT[22] = REG_B[22];
  assign REG_B_OUT[21] = REG_B[21];
  assign REG_B_OUT[20] = REG_B[20];
  assign REG_B_OUT[19] = REG_B[19];
  assign REG_B_OUT[18] = REG_B[18];
  assign REG_B_OUT[17] = REG_B[17];
  assign REG_B_OUT[16] = REG_B[16];
  assign REG_B_OUT[15] = REG_B[15];
  assign REG_B_OUT[14] = REG_B[14];
  assign REG_B_OUT[13] = REG_B[13];
  assign REG_B_OUT[12] = REG_B[12];
  assign REG_B_OUT[11] = REG_B[11];
  assign REG_B_OUT[10] = REG_B[10];
  assign REG_B_OUT[9] = REG_B[9];
  assign REG_B_OUT[8] = REG_B[8];
  assign REG_B_OUT[7] = REG_B[7];
  assign REG_B_OUT[6] = REG_B[6];
  assign REG_B_OUT[5] = REG_B[5];
  assign REG_B_OUT[4] = REG_B[4];
  assign REG_B_OUT[3] = REG_B[3];
  assign REG_B_OUT[2] = REG_B[2];
  assign REG_B_OUT[1] = REG_B[1];
  assign REG_B_OUT[0] = REG_B[0];

  MUX41_GEN_N32_3 OP_A_SEL_MUX ( .A(REG_A), .B(FORW_ALU_MEM), .C(FORW_ALU_WB), 
        .D(FORW_MEM_WB), .SEL(OP_SEL_A), .Y(IN_A_ALU_SIG) );
  MUX51_GEN_N32_0 OP_B_SEL_MUX ( .A(REG_B), .B(FORW_ALU_MEM), .C(FORW_ALU_WB), 
        .D(FORW_MEM_WB), .E(IMMEDIATE), .SEL(OP_SEL_B), .Y(IN_B_ALU_SIG) );
  ALU_N32_ALU_SIZE5 ALUCOMP ( .IN_A(IN_A_ALU_SIG), .IN_B(IN_B_ALU_SIG), 
        .ALU_OP_CODE(ALU_CODE), .CLK(CLK), .RST(RST), .RST_DIV(RST_DIV), 
        .OUT_ALU(OUTPUT_ALU) );
endmodule


module REG_N5_0 ( D, Q, EN, RST, CLK );
  input [4:0] D;
  output [4:0] Q;
  input EN, RST, CLK;


  FD_1_420 FF_0 ( .D(D[0]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[0]) );
  FD_1_419 FF_1 ( .D(D[1]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[1]) );
  FD_1_418 FF_2 ( .D(D[2]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[2]) );
  FD_1_417 FF_3 ( .D(D[3]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[3]) );
  FD_1_416 FF_4 ( .D(D[4]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[4]) );
endmodule


module XOR_GATE_0 ( A, B, Y );
  input A, B;
  output Y;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(Y) );
endmodule


module AND_GATE_0 ( A, B, Y );
  input A, B;
  output Y;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module INV_0 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module DECODE_N32_N_ADDR5_IMM_SIZE16_OP_CODE_SIZE6 ( CLK, INSTRUCTION, NPC, 
        CONFIRM_JMP, CONFIRM_BRANCH, BRANCH_TYPE, EN, RST, RD1, RD2, WR, 
        SEL_DEST, LHI_SEL, JMP_SEL, SEL_MUX_BRANCH, FORW_ALU_MEM, FORW_ALU_WB, 
        FORW_MEM_WB, DATA_IN, ADDR_WR, PC_SEL_MUX, NPC_OUT, NPC_ADDED, REG_A, 
        REG_B, IMMEDIATE, DEST_REG );
  input [31:0] INSTRUCTION;
  input [31:0] NPC;
  input [1:0] SEL_DEST;
  input [1:0] SEL_MUX_BRANCH;
  input [31:0] FORW_ALU_MEM;
  input [31:0] FORW_ALU_WB;
  input [31:0] FORW_MEM_WB;
  input [31:0] DATA_IN;
  input [4:0] ADDR_WR;
  output [31:0] NPC_OUT;
  output [31:0] NPC_ADDED;
  output [31:0] REG_A;
  output [31:0] REG_B;
  output [31:0] IMMEDIATE;
  output [4:0] DEST_REG;
  input CLK, CONFIRM_JMP, CONFIRM_BRANCH, BRANCH_TYPE, EN, RST, RD1, RD2, WR,
         LHI_SEL, JMP_SEL;
  output PC_SEL_MUX;
  wire   n1, n2;
  wire   [31:0] OUT_ADDER;
  wire   [31:0] IN_A_BRANCH;
  assign NPC_OUT[31] = NPC[31];
  assign NPC_OUT[30] = NPC[30];
  assign NPC_OUT[29] = NPC[29];
  assign NPC_OUT[28] = NPC[28];
  assign NPC_OUT[27] = NPC[27];
  assign NPC_OUT[26] = NPC[26];
  assign NPC_OUT[25] = NPC[25];
  assign NPC_OUT[24] = NPC[24];
  assign NPC_OUT[23] = NPC[23];
  assign NPC_OUT[22] = NPC[22];
  assign NPC_OUT[21] = NPC[21];
  assign NPC_OUT[20] = NPC[20];
  assign NPC_OUT[19] = NPC[19];
  assign NPC_OUT[18] = NPC[18];
  assign NPC_OUT[17] = NPC[17];
  assign NPC_OUT[16] = NPC[16];
  assign NPC_OUT[15] = NPC[15];
  assign NPC_OUT[14] = NPC[14];
  assign NPC_OUT[13] = NPC[13];
  assign NPC_OUT[12] = NPC[12];
  assign NPC_OUT[11] = NPC[11];
  assign NPC_OUT[10] = NPC[10];
  assign NPC_OUT[9] = NPC[9];
  assign NPC_OUT[8] = NPC[8];
  assign NPC_OUT[7] = NPC[7];
  assign NPC_OUT[6] = NPC[6];
  assign NPC_OUT[5] = NPC[5];
  assign NPC_OUT[4] = NPC[4];
  assign NPC_OUT[3] = NPC[3];
  assign NPC_OUT[2] = NPC[2];
  assign NPC_OUT[1] = NPC[1];
  assign NPC_OUT[0] = NPC[0];

  REG_FILE_N32_N_ADDR5 REG_FILE_INST ( .CLK(CLK), .RST(RST), .EN(EN), .RD1(RD1), .RD2(RD2), .WR(WR), .ADDR_WR(ADDR_WR), .ADDR_RD1(INSTRUCTION[25:21]), 
        .ADDR_RD2(INSTRUCTION[20:16]), .DATA_IN(DATA_IN), .DATA_OUT_1(REG_A), 
        .DATA_OUT_2(REG_B) );
  MUX31_GEN_N5 DEST_MUX ( .A(INSTRUCTION[20:16]), .B({n2, INSTRUCTION[14:11]}), 
        .C({1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .SEL(SEL_DEST), .Y(DEST_REG) );
  MUX21_GEN_N32_5 IMMEDIATE_MUX ( .A({n2, INSTRUCTION[14:0], 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({n2, n2, n2, n2, n2, n2, n2, n2, n2, n2, n2, n2, n2, n2, n2, 
        n2, n2, INSTRUCTION[14:0]}), .SEL(LHI_SEL), .Y(IMMEDIATE) );
  MUX21_GEN_N32_4 NPC_MUX ( .A(REG_A), .B(OUT_ADDER), .SEL(JMP_SEL), .Y(
        NPC_ADDED) );
  CSA_N4_0 BRANCH_JMP_ADDER_0 ( .A(NPC[3:0]), .B(INSTRUCTION[3:0]), .Ci(1'b0), 
        .S(OUT_ADDER[3:0]) );
  CSA_N4_15 BRANCH_JMP_ADDER_1 ( .A(NPC[7:4]), .B(INSTRUCTION[7:4]), .Ci(1'b0), 
        .S(OUT_ADDER[7:4]) );
  CSA_N4_14 BRANCH_JMP_ADDER_2 ( .A(NPC[11:8]), .B(INSTRUCTION[11:8]), .Ci(
        1'b0), .S(OUT_ADDER[11:8]) );
  CSA_N4_13 BRANCH_JMP_ADDER_3 ( .A(NPC[15:12]), .B({n1, INSTRUCTION[14:12]}), 
        .Ci(1'b0), .S(OUT_ADDER[15:12]) );
  CSA_N4_12 BRANCH_JMP_ADDER_4 ( .A(NPC[19:16]), .B({n1, n1, n1, n1}), .Ci(
        1'b0), .S(OUT_ADDER[19:16]) );
  CSA_N4_11 BRANCH_JMP_ADDER_5 ( .A(NPC[23:20]), .B({n1, n1, n1, n1}), .Ci(
        1'b0), .S(OUT_ADDER[23:20]) );
  CSA_N4_10 BRANCH_JMP_ADDER_6 ( .A(NPC[27:24]), .B({n1, n1, n1, n1}), .Ci(
        1'b0), .S(OUT_ADDER[27:24]) );
  CSA_N4_9 BRANCH_JMP_ADDER_7 ( .A(NPC[31:28]), .B({n2, n2, n2, n2}), .Ci(1'b0), .S(OUT_ADDER[31:28]) );
  MUX41_GEN_N32_0 FORW_BRANCH_MUX ( .A(FORW_MEM_WB), .B(FORW_ALU_WB), .C(
        FORW_ALU_MEM), .D(REG_A), .SEL(SEL_MUX_BRANCH), .Y(IN_A_BRANCH) );
  BRANCH_N32 INST_BRANCH ( .REG_A(IN_A_BRANCH), .BNEZ_SEL(BRANCH_TYPE), 
        .CONFIRM_BRANCH(CONFIRM_BRANCH), .CONFIRM_JMP(CONFIRM_JMP), 
        .BRANCH_SEL(PC_SEL_MUX) );
  BUF_X2 U3 ( .A(INSTRUCTION[15]), .Z(n1) );
  BUF_X1 U4 ( .A(INSTRUCTION[15]), .Z(n2) );
endmodule


module REG_N32_0 ( D, Q, EN, RST, CLK );
  input [31:0] D;
  output [31:0] Q;
  input EN, RST, CLK;
  wire   n1, n2, n3, n4, n5, n6;

  FD_1_580 FF_0 ( .D(D[0]), .CLK(CLK), .EN(n4), .RST(n2), .Q(Q[0]) );
  FD_1_579 FF_1 ( .D(D[1]), .CLK(CLK), .EN(n4), .RST(n2), .Q(Q[1]) );
  FD_1_578 FF_2 ( .D(D[2]), .CLK(CLK), .EN(n4), .RST(n2), .Q(Q[2]) );
  FD_1_577 FF_3 ( .D(D[3]), .CLK(CLK), .EN(n4), .RST(n2), .Q(Q[3]) );
  FD_1_576 FF_4 ( .D(D[4]), .CLK(CLK), .EN(n4), .RST(n2), .Q(Q[4]) );
  FD_1_575 FF_5 ( .D(D[5]), .CLK(CLK), .EN(n4), .RST(n2), .Q(Q[5]) );
  FD_1_574 FF_6 ( .D(D[6]), .CLK(CLK), .EN(n4), .RST(n2), .Q(Q[6]) );
  FD_1_573 FF_7 ( .D(D[7]), .CLK(CLK), .EN(n4), .RST(n3), .Q(Q[7]) );
  FD_1_572 FF_8 ( .D(D[8]), .CLK(CLK), .EN(n4), .RST(n3), .Q(Q[8]) );
  FD_1_571 FF_9 ( .D(D[9]), .CLK(CLK), .EN(n4), .RST(n3), .Q(Q[9]) );
  FD_1_570 FF_10 ( .D(D[10]), .CLK(CLK), .EN(n4), .RST(n3), .Q(Q[10]) );
  FD_1_569 FF_11 ( .D(D[11]), .CLK(CLK), .EN(n4), .RST(n3), .Q(Q[11]) );
  FD_1_568 FF_12 ( .D(D[12]), .CLK(CLK), .EN(n4), .RST(n1), .Q(Q[12]) );
  FD_1_567 FF_13 ( .D(D[13]), .CLK(CLK), .EN(n5), .RST(n1), .Q(Q[13]) );
  FD_1_566 FF_14 ( .D(D[14]), .CLK(CLK), .EN(n5), .RST(n1), .Q(Q[14]) );
  FD_1_565 FF_15 ( .D(D[15]), .CLK(CLK), .EN(n5), .RST(n1), .Q(Q[15]) );
  FD_1_564 FF_16 ( .D(D[16]), .CLK(CLK), .EN(n5), .RST(n1), .Q(Q[16]) );
  FD_1_563 FF_17 ( .D(D[17]), .CLK(CLK), .EN(n5), .RST(n1), .Q(Q[17]) );
  FD_1_562 FF_18 ( .D(D[18]), .CLK(CLK), .EN(n5), .RST(n1), .Q(Q[18]) );
  FD_1_561 FF_19 ( .D(D[19]), .CLK(CLK), .EN(n5), .RST(n1), .Q(Q[19]) );
  FD_1_560 FF_20 ( .D(D[20]), .CLK(CLK), .EN(n5), .RST(n1), .Q(Q[20]) );
  FD_1_559 FF_21 ( .D(D[21]), .CLK(CLK), .EN(n5), .RST(n2), .Q(Q[21]) );
  FD_1_558 FF_22 ( .D(D[22]), .CLK(CLK), .EN(n5), .RST(n2), .Q(Q[22]) );
  FD_1_557 FF_23 ( .D(D[23]), .CLK(CLK), .EN(n5), .RST(n2), .Q(Q[23]) );
  FD_1_556 FF_24 ( .D(D[24]), .CLK(CLK), .EN(n5), .RST(n2), .Q(Q[24]) );
  FD_1_555 FF_25 ( .D(D[25]), .CLK(CLK), .EN(n5), .RST(n2), .Q(Q[25]) );
  FD_1_554 FF_26 ( .D(D[26]), .CLK(CLK), .EN(n6), .RST(n2), .Q(Q[26]) );
  FD_1_553 FF_27 ( .D(D[27]), .CLK(CLK), .EN(n6), .RST(n1), .Q(Q[27]) );
  FD_1_552 FF_28 ( .D(D[28]), .CLK(CLK), .EN(n6), .RST(n1), .Q(Q[28]) );
  FD_1_551 FF_29 ( .D(D[29]), .CLK(CLK), .EN(n6), .RST(n1), .Q(Q[29]) );
  FD_1_550 FF_30 ( .D(D[30]), .CLK(CLK), .EN(n6), .RST(n1), .Q(Q[30]) );
  FD_1_549 FF_31 ( .D(D[31]), .CLK(CLK), .EN(n6), .RST(n3), .Q(Q[31]) );
  BUF_X1 U1 ( .A(EN), .Z(n4) );
  BUF_X1 U2 ( .A(EN), .Z(n5) );
  BUF_X1 U3 ( .A(EN), .Z(n6) );
  BUF_X1 U4 ( .A(RST), .Z(n2) );
  BUF_X1 U5 ( .A(RST), .Z(n1) );
  BUF_X1 U6 ( .A(RST), .Z(n3) );
endmodule


module BPU_N32_OP_CODE_SIZE6_SET_BIT2 ( CLK, RST, STALL_BRANCH, BRANCH_DEC, 
        BRANCH_FETCH, DEST_DEC, PC_IN, PC_OUT, MUX_SEL );
  input [5:0] BRANCH_FETCH;
  input [31:0] DEST_DEC;
  input [31:0] PC_IN;
  output [31:0] PC_OUT;
  input CLK, RST, STALL_BRANCH, BRANCH_DEC;
  output MUX_SEL;
  wire   EN_BPU, MUX_SEL_SIG, HIT_MISS, DIS_FSM, LOAD, EN_FSM_SIG, n4, n5, n6;
  wire   [1:0] FSM_SEL;
  wire   [2:0] EN_FSM_VECT;
  wire   [2:0] OUT_AND;

  CACHE_BPU_N32_SET_BIT2 CACHE_INST ( .ADDR(PC_IN), .DATA_IN(DEST_DEC), 
        .DATA_OUT(PC_OUT), .ENC(FSM_SEL), .RST(RST), .LOAD(LOAD), .CLK(CLK), 
        .HIT_MISS(HIT_MISS) );
  FSM_BPU FSM_INST ( .RST(RST), .CLK(CLK), .BRANCH_TAKEN(BRANCH_DEC), .EN_FSM(
        EN_FSM_SIG), .FSM_SEL(FSM_SEL), .MUX_SEL(MUX_SEL_SIG) );
  CU_BPU CU_INST ( .HIT_MISS(HIT_MISS), .BRANCH_FETCH(EN_BPU), .CLK(CLK), 
        .RST(RST), .BRANCH_TAKEN(BRANCH_DEC), .NEW_BRANCH(LOAD), .EN_FSM(
        EN_FSM_VECT[0]) );
  FD_1_0 FDs_0 ( .D(EN_FSM_VECT[0]), .CLK(CLK), .EN(STALL_BRANCH), .RST(
        DIS_FSM), .Q(EN_FSM_VECT[1]) );
  FD_1_581 FDs_1 ( .D(EN_FSM_VECT[1]), .CLK(CLK), .EN(STALL_BRANCH), .RST(
        DIS_FSM), .Q(EN_FSM_VECT[2]) );
  AND_GATE_1_0 ANDs_0 ( .A(EN_FSM_VECT[0]), .B(DIS_FSM), .Y(OUT_AND[0]) );
  AND_GATE_1_737 ANDs_1 ( .A(EN_FSM_VECT[1]), .B(DIS_FSM), .Y(OUT_AND[1]) );
  AND_GATE_1_736 ANDs_2 ( .A(EN_FSM_VECT[2]), .B(DIS_FSM), .Y(OUT_AND[2]) );
  N_OR_N3 OR_INST ( .A(OUT_AND), .Y(EN_FSM_SIG) );
  INV_X1 U2 ( .A(STALL_BRANCH), .ZN(DIS_FSM) );
  NOR3_X1 U3 ( .A1(BRANCH_FETCH[3]), .A2(BRANCH_FETCH[5]), .A3(n4), .ZN(EN_BPU) );
  AOI22_X1 U4 ( .A1(n5), .A2(BRANCH_FETCH[2]), .B1(BRANCH_FETCH[1]), .B2(n6), 
        .ZN(n4) );
  INV_X1 U5 ( .A(BRANCH_FETCH[2]), .ZN(n6) );
  NOR2_X1 U6 ( .A1(BRANCH_FETCH[4]), .A2(BRANCH_FETCH[1]), .ZN(n5) );
  AND2_X1 U7 ( .A1(MUX_SEL_SIG), .A2(HIT_MISS), .ZN(MUX_SEL) );
endmodule


module FETCH_N32 ( JUMP_ADDR, BPU_ADDR, NPC_IN, BRANCH_SEL, BRANCH_SEL_BPU, 
        SEL_N_TAKEN, EN, RST, CLK, DATA_IN_INSTR, H_M_CACHE, ADDR_IRAM, PC_OUT, 
        NPC, INSTRUCTION );
  input [31:0] JUMP_ADDR;
  input [31:0] BPU_ADDR;
  input [31:0] NPC_IN;
  input [7:0] DATA_IN_INSTR;
  output [31:0] ADDR_IRAM;
  output [31:0] PC_OUT;
  output [31:0] NPC;
  output [31:0] INSTRUCTION;
  input BRANCH_SEL, BRANCH_SEL_BPU, SEL_N_TAKEN, EN, RST, CLK;
  output H_M_CACHE;
  wire   CACHE_LOAD;
  wire   [31:0] OUT_MUX_2;
  wire   [31:0] OUT_MUX;
  wire   [31:0] OUT_MUX_1;
  assign PC_OUT[1] = NPC[1];
  assign PC_OUT[0] = NPC[0];

  REG_N32_2 PC ( .D(OUT_MUX_2), .Q({PC_OUT[31:2], NPC[1:0]}), .EN(EN), .RST(
        RST), .CLK(CLK) );
  CACHE_N32_TAG_BIT23_SET_BIT4_N_DATA5 INSTRUCTION_CACHE ( .ADDR({PC_OUT[31:2], 
        NPC[1:0]}), .ADDR_OUT(ADDR_IRAM), .DATA_IN(DATA_IN_INSTR), .DATA_OUT(
        INSTRUCTION), .RST(RST), .LOAD(CACHE_LOAD), .CLK(CLK), .HIT_MISS(
        H_M_CACHE) );
  RCA_GEN_NO_C_N30 PC_ADDER ( .A(PC_OUT[31:2]), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b1}), .S(NPC[31:2]) );
  MUX21_GEN_N32_0 MUX_PC ( .A(JUMP_ADDR), .B(NPC), .SEL(BRANCH_SEL), .Y(
        OUT_MUX) );
  MUX21_GEN_N32_7 MUX_BPU ( .A(BPU_ADDR), .B(OUT_MUX), .SEL(BRANCH_SEL_BPU), 
        .Y(OUT_MUX_1) );
  MUX21_GEN_N32_6 MUX_N_TAKEN ( .A(NPC_IN), .B(OUT_MUX_1), .SEL(SEL_N_TAKEN), 
        .Y(OUT_MUX_2) );
  NOR2_X1 U3 ( .A1(RST), .A2(H_M_CACHE), .ZN(CACHE_LOAD) );
endmodule


module FD_0 ( D, CLK, EN, RST, Q );
  input D, CLK, EN, RST;
  output Q;
  wire   n2, n3, n5;

  DFF_X1 Q_reg ( .D(n5), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(RST), .A2(n2), .ZN(n5) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n3), .ZN(n2) );
  INV_X1 U5 ( .A(EN), .ZN(n3) );
endmodule


module REG_N3 ( D, Q, EN, RST, CLK );
  input [2:0] D;
  output [2:0] Q;
  input EN, RST, CLK;


  FD_147 FF_0 ( .D(D[0]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[0]) );
  FD_146 FF_1 ( .D(D[1]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[1]) );
  FD_145 FF_2 ( .D(D[2]), .CLK(CLK), .EN(EN), .RST(RST), .Q(Q[2]) );
endmodule


module REG_N11 ( D, Q, EN, RST, CLK );
  input [10:0] D;
  output [10:0] Q;
  input EN, RST, CLK;
  wire   n1;

  FD_158 FF_0 ( .D(D[0]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[0]) );
  FD_157 FF_1 ( .D(D[1]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[1]) );
  FD_156 FF_2 ( .D(D[2]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[2]) );
  FD_155 FF_3 ( .D(D[3]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[3]) );
  FD_154 FF_4 ( .D(D[4]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[4]) );
  FD_153 FF_5 ( .D(D[5]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[5]) );
  FD_152 FF_6 ( .D(D[6]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[6]) );
  FD_151 FF_7 ( .D(D[7]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[7]) );
  FD_150 FF_8 ( .D(D[8]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[8]) );
  FD_149 FF_9 ( .D(D[9]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[9]) );
  FD_148 FF_10 ( .D(D[10]), .CLK(CLK), .EN(EN), .RST(n1), .Q(Q[10]) );
  BUF_X1 U1 ( .A(RST), .Z(n1) );
endmodule


module REG_N18 ( D, Q, EN, RST, CLK );
  input [17:0] D;
  output [17:0] Q;
  input EN, RST, CLK;
  wire   n1, n2, n3, n4;

  FD_176 FF_0 ( .D(D[0]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[0]) );
  FD_175 FF_1 ( .D(D[1]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[1]) );
  FD_174 FF_2 ( .D(D[2]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[2]) );
  FD_173 FF_3 ( .D(D[3]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[3]) );
  FD_172 FF_4 ( .D(D[4]), .CLK(CLK), .EN(n1), .RST(n4), .Q(Q[4]) );
  FD_171 FF_5 ( .D(D[5]), .CLK(CLK), .EN(n1), .RST(n3), .Q(Q[5]) );
  FD_170 FF_6 ( .D(D[6]), .CLK(CLK), .EN(n1), .RST(n3), .Q(Q[6]) );
  FD_169 FF_7 ( .D(D[7]), .CLK(CLK), .EN(n1), .RST(n3), .Q(Q[7]) );
  FD_168 FF_8 ( .D(D[8]), .CLK(CLK), .EN(n1), .RST(n3), .Q(Q[8]) );
  FD_167 FF_9 ( .D(D[9]), .CLK(CLK), .EN(n1), .RST(n3), .Q(Q[9]) );
  FD_166 FF_10 ( .D(D[10]), .CLK(CLK), .EN(n1), .RST(n3), .Q(Q[10]) );
  FD_165 FF_11 ( .D(D[11]), .CLK(CLK), .EN(n1), .RST(n3), .Q(Q[11]) );
  FD_164 FF_12 ( .D(D[12]), .CLK(CLK), .EN(n1), .RST(n3), .Q(Q[12]) );
  FD_163 FF_13 ( .D(D[13]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[13]) );
  FD_162 FF_14 ( .D(D[14]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[14]) );
  FD_161 FF_15 ( .D(D[15]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[15]) );
  FD_160 FF_16 ( .D(D[16]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[16]) );
  FD_159 FF_17 ( .D(D[17]), .CLK(CLK), .EN(n2), .RST(n3), .Q(Q[17]) );
  BUF_X1 U1 ( .A(EN), .Z(n2) );
  BUF_X1 U2 ( .A(EN), .Z(n1) );
  BUF_X1 U3 ( .A(RST), .Z(n4) );
  BUF_X1 U4 ( .A(RST), .Z(n3) );
endmodule


module DATAPATH_N32_N_ADDR5_IMM_SIZE16_OP_CODE_SIZE6_M5_ALUSIZE5 ( CLK, RST, 
        EN_PC, EN_1, EN_2, CONFIRM_JMP, CONFIRM_BRANCH, BRANCH_TYPE, RD1, RD2, 
        WR, SEL_DEST, LHI_SEL, JMP_SEL, EN_3, ALU_CODE, OP_SEL, EN_4, 
        STORE_MASK, LOAD_TYPE, SEL, DATA_IN_IRAM, DATA_IN_MEM, DATA_OUT_MEM, 
        ADDR_MEM, INSTR_CACHE_H_M, ADDR_IRAM, INSTR, STALL, STALL_BRANCH, 
        WRONG_FETCH );
  input [1:0] SEL_DEST;
  input [4:0] ALU_CODE;
  input [1:0] STORE_MASK;
  input [2:0] LOAD_TYPE;
  input [1:0] SEL;
  input [7:0] DATA_IN_IRAM;
  input [31:0] DATA_IN_MEM;
  output [31:0] DATA_OUT_MEM;
  output [31:0] ADDR_MEM;
  output [31:0] ADDR_IRAM;
  output [31:0] INSTR;
  input CLK, RST, EN_PC, EN_1, EN_2, CONFIRM_JMP, CONFIRM_BRANCH, BRANCH_TYPE,
         RD1, RD2, WR, LHI_SEL, JMP_SEL, EN_3, OP_SEL, EN_4;
  output INSTR_CACHE_H_M, STALL, STALL_BRANCH, WRONG_FETCH;
  wire   BPU_SEL, WRONG_FETCH_SIG_1, BPU_SEL_SIG, BRANCH_SEL_DECODE_FETCH,
         SEL_N_TAKEN, BRANCH_SEL_ID, BPU_ID, N_BPU_ID, RST_DIV_SIG, n2, n1, n3,
         n4, n5, n6;
  wire   [1:0] OP_SEL_B_SIG;
  wire   [31:0] NPC_DECODE_OUT_FETCH_IN;
  wire   [31:0] PC_BPU_OUT;
  wire   [31:0] NPC_DECODE_OUT_FETCH_IN_OLD;
  wire   [31:0] PC_BPU_IN;
  wire   [31:0] NPC_FETCH_OUT;
  wire   [31:0] NPC_DECODE_IN;
  wire   [31:0] INSTRUCTION_DECODE_IN;
  wire   [1:0] FORW_SEL_D;
  wire   [31:0] ALU_MEM_IN;
  wire   [31:0] OUT_ALU_WB_IN;
  wire   [31:0] MEMORY_OUT_WB_IN;
  wire   [31:0] DATA_DECODE_IN;
  wire   [4:0] ADDR_WR_DECODE_IN;
  wire   [31:0] REG_A_DECODE_OUT;
  wire   [31:0] REG_B_DECODE_OUT;
  wire   [31:0] IMMEDIATE_DECODE_OUT;
  wire   [4:0] DEST_REG_DECODE_OUT;
  wire   [31:0] REG_A_EXECUTE_IN;
  wire   [31:0] REG_B_EXECUTE_IN;
  wire   [31:0] IMMEDIATE_EXECUTE_IN;
  wire   [4:0] DEST_REG_EXECUTE_IN;
  wire   [31:0] NPC_OUT_EX_IN_MEM;
  wire   [1:0] FORW_SEL_A;
  wire   [4:0] DEST_REG_EXECUTE_OUT;
  wire   [31:0] ALU_EXECUTE_OUT;
  wire   [31:0] REG_B_EXECUTE_OUT;
  wire   [4:0] DEST_REG_MEM_IN;
  wire   [31:0] REG_B_MEM_IN;
  wire   [31:0] NPC_OUT_MEM_IN_WB;
  wire   [31:0] WB_OUT_REG_B;
  wire   [1:0] FORW_SEL_C;
  wire   [4:0] DEST_REG_MEM_OUT;
  wire   [31:0] MEMORY_OUT_MEM_OUT;
  wire   [31:0] OUT_ALU_MEM_OUT;
  wire   [4:0] DEST_REG_WB_IN;
  wire   [31:0] NPC_OUT_WB_IN;

  FETCH_N32 INST_FETCH ( .JUMP_ADDR(NPC_DECODE_OUT_FETCH_IN), .BPU_ADDR(
        PC_BPU_OUT), .NPC_IN(NPC_DECODE_OUT_FETCH_IN_OLD), .BRANCH_SEL(
        BRANCH_SEL_DECODE_FETCH), .BRANCH_SEL_BPU(BPU_SEL_SIG), .SEL_N_TAKEN(
        SEL_N_TAKEN), .EN(EN_1), .RST(n5), .CLK(CLK), .DATA_IN_INSTR(
        DATA_IN_IRAM), .H_M_CACHE(INSTR_CACHE_H_M), .ADDR_IRAM(ADDR_IRAM), 
        .PC_OUT(PC_BPU_IN), .NPC(NPC_FETCH_OUT), .INSTRUCTION(INSTR) );
  BPU_N32_OP_CODE_SIZE6_SET_BIT2 INST_BPU ( .CLK(CLK), .RST(n4), 
        .STALL_BRANCH(STALL_BRANCH), .BRANCH_DEC(BRANCH_SEL_ID), 
        .BRANCH_FETCH(INSTR[31:26]), .DEST_DEC(NPC_DECODE_OUT_FETCH_IN), 
        .PC_IN(PC_BPU_IN), .PC_OUT(PC_BPU_OUT), .MUX_SEL(BPU_SEL) );
  REG_N32_0 PIPE_IF_ID_NPC ( .D(NPC_FETCH_OUT), .Q(NPC_DECODE_IN), .EN(EN_1), 
        .RST(n5), .CLK(CLK) );
  REG_N32_14 PIPE_IF_ID_INSTRUCTION ( .D(INSTR), .Q(INSTRUCTION_DECODE_IN), 
        .EN(EN_1), .RST(n5), .CLK(CLK) );
  FD_178 PIPE_IF_ID_BPU ( .D(BPU_SEL), .CLK(CLK), .EN(EN_1), .RST(n4), .Q(
        BPU_ID) );
  DECODE_N32_N_ADDR5_IMM_SIZE16_OP_CODE_SIZE6 INST_DECODE ( .CLK(CLK), 
        .INSTRUCTION(INSTRUCTION_DECODE_IN), .NPC(NPC_DECODE_IN), 
        .CONFIRM_JMP(CONFIRM_JMP), .CONFIRM_BRANCH(CONFIRM_BRANCH), 
        .BRANCH_TYPE(BRANCH_TYPE), .EN(n3), .RST(n5), .RD1(RD1), .RD2(RD2), 
        .WR(WR), .SEL_DEST(SEL_DEST), .LHI_SEL(LHI_SEL), .JMP_SEL(JMP_SEL), 
        .SEL_MUX_BRANCH(FORW_SEL_D), .FORW_ALU_MEM(ALU_MEM_IN), .FORW_ALU_WB(
        OUT_ALU_WB_IN), .FORW_MEM_WB(MEMORY_OUT_WB_IN), .DATA_IN(
        DATA_DECODE_IN), .ADDR_WR(ADDR_WR_DECODE_IN), .PC_SEL_MUX(
        BRANCH_SEL_ID), .NPC_OUT(NPC_DECODE_OUT_FETCH_IN_OLD), .NPC_ADDED(
        NPC_DECODE_OUT_FETCH_IN), .REG_A(REG_A_DECODE_OUT), .REG_B(
        REG_B_DECODE_OUT), .IMMEDIATE(IMMEDIATE_DECODE_OUT), .DEST_REG(
        DEST_REG_DECODE_OUT) );
  INV_0 INV_BPU ( .A(BPU_ID), .Y(N_BPU_ID) );
  AND_GATE_0 CORR_BRANCH ( .A(N_BPU_ID), .B(BRANCH_SEL_ID), .Y(
        BRANCH_SEL_DECODE_FETCH) );
  AND_GATE_340 SEL_MUX_N_TAKEN ( .A(WRONG_FETCH), .B(BPU_ID), .Y(SEL_N_TAKEN)
         );
  XOR_GATE_0 PREDICTION ( .A(BPU_ID), .B(BRANCH_SEL_ID), .Y(WRONG_FETCH) );
  FD_177 DELAY_MUX ( .D(WRONG_FETCH), .CLK(CLK), .EN(1'b1), .RST(n5), .Q(
        WRONG_FETCH_SIG_1) );
  REG_N32_13 PIPE_ID_EX_REG_A ( .D(REG_A_DECODE_OUT), .Q(REG_A_EXECUTE_IN), 
        .EN(n3), .RST(n6), .CLK(CLK) );
  REG_N32_12 PIPE_ID_EX_REG_B ( .D(REG_B_DECODE_OUT), .Q(REG_B_EXECUTE_IN), 
        .EN(n3), .RST(n6), .CLK(CLK) );
  REG_N32_11 PIPE_ID_EX_IMMEDIATE ( .D(IMMEDIATE_DECODE_OUT), .Q(
        IMMEDIATE_EXECUTE_IN), .EN(n3), .RST(n6), .CLK(CLK) );
  REG_N5_0 PIPE_ID_EX_DEST_REG ( .D(DEST_REG_DECODE_OUT), .Q(
        DEST_REG_EXECUTE_IN), .EN(n3), .RST(n5), .CLK(CLK) );
  REG_N32_10 PIPE_ID_EX_OUT_NPC ( .D(NPC_DECODE_IN), .Q(NPC_OUT_EX_IN_MEM), 
        .EN(n3), .RST(n6), .CLK(CLK) );
  EXECUTE_N32_N_ADDR5_ALUSIZE5 INST_EXECUTE ( .REG_A(REG_A_EXECUTE_IN), 
        .REG_B(REG_B_EXECUTE_IN), .IMMEDIATE(IMMEDIATE_EXECUTE_IN), 
        .FORW_ALU_MEM(ALU_MEM_IN), .FORW_ALU_WB(OUT_ALU_WB_IN), .FORW_MEM_WB(
        MEMORY_OUT_WB_IN), .DEST_REG_IN(DEST_REG_EXECUTE_IN), .ALU_CODE(
        ALU_CODE), .OP_SEL_A(FORW_SEL_A), .OP_SEL_B({OP_SEL, OP_SEL_B_SIG}), 
        .CLK(CLK), .RST(n5), .DEST_REG_OUT(DEST_REG_EXECUTE_OUT), .OUTPUT_ALU(
        ALU_EXECUTE_OUT), .RST_DIV(RST_DIV_SIG), .REG_B_OUT(REG_B_EXECUTE_OUT)
         );
  REG_N5_2 PIPE_EX_MEM_DEST_REG ( .D(DEST_REG_EXECUTE_OUT), .Q(DEST_REG_MEM_IN), .EN(EN_3), .RST(n4), .CLK(CLK) );
  REG_N32_9 PIPE_EX_MEM_OUTPUT_ALU ( .D(ALU_EXECUTE_OUT), .Q(ALU_MEM_IN), .EN(
        EN_3), .RST(n6), .CLK(CLK) );
  REG_N32_8 PIPE_EX_MEM_REG_B ( .D(REG_B_EXECUTE_OUT), .Q(REG_B_MEM_IN), .EN(
        EN_3), .RST(n6), .CLK(CLK) );
  REG_N32_7 PIPE_EX_MEM_OUT_NPC ( .D(NPC_OUT_EX_IN_MEM), .Q(NPC_OUT_MEM_IN_WB), 
        .EN(EN_3), .RST(n6), .CLK(CLK) );
  MEMORY_N32_N_ADDR5 INST_MEMORY ( .IN_ALU(ALU_MEM_IN), .DEST_REG_IN(
        DEST_REG_MEM_IN), .REG_B_IN(REG_B_MEM_IN), .FORW_ALU_WB(OUT_ALU_WB_IN), 
        .FORW_MEM_WB(MEMORY_OUT_WB_IN), .FORW_REG(WB_OUT_REG_B), .SEL_DATA(
        FORW_SEL_C), .RESET(n4), .ENABLE(n1), .DATA_IN_MEM(DATA_IN_MEM), 
        .LOAD_TYPE(LOAD_TYPE), .STORE_MASK(STORE_MASK), .ADDR_MEM(ADDR_MEM), 
        .DATA_OUT_MEM(DATA_OUT_MEM), .DEST_REG_OUT(DEST_REG_MEM_OUT), 
        .MEMORY_OUT(MEMORY_OUT_MEM_OUT), .OUT_ALU(OUT_ALU_MEM_OUT) );
  REG_N5_1 PIPE_MEM_WB_DEST_REG ( .D(DEST_REG_MEM_OUT), .Q(DEST_REG_WB_IN), 
        .EN(n1), .RST(n4), .CLK(CLK) );
  REG_N32_6 PIPE_MEM_WB_MEMORY_OUT ( .D(MEMORY_OUT_MEM_OUT), .Q(
        MEMORY_OUT_WB_IN), .EN(n1), .RST(n6), .CLK(CLK) );
  REG_N32_5 PIPE_MEM_WB_OUT_ALU ( .D(OUT_ALU_MEM_OUT), .Q(OUT_ALU_WB_IN), .EN(
        n1), .RST(n6), .CLK(CLK) );
  REG_N32_4 PIPE_MEM_WB_OUT_NPC ( .D(NPC_OUT_MEM_IN_WB), .Q(NPC_OUT_WB_IN), 
        .EN(n1), .RST(n6), .CLK(CLK) );
  WB_N32_N_ADDR5 INST_WB ( .IN_MEM(MEMORY_OUT_WB_IN), .IN_ALU(OUT_ALU_WB_IN), 
        .IN_NPC(NPC_OUT_WB_IN), .SEL(SEL), .DEST_REG_IN(DEST_REG_WB_IN), 
        .DEST_REG_OUT(ADDR_WR_DECODE_IN), .OUT_WB(DATA_DECODE_IN) );
  REG_N32_3 PIPE_WB_OUT ( .D(DATA_DECODE_IN), .Q(WB_OUT_REG_B), .EN(1'b1), 
        .RST(n5), .CLK(CLK) );
  FORWARD_UNIT_OPCODE_SIZE6_N_ADDR5 FORW_INST ( .CLK(CLK), .RST(n6), 
        .OPCODE_IF(INSTR[31:26]), .REG_A_IF(INSTR[25:21]), .OPCODE_ID(
        INSTRUCTION_DECODE_IN[31:26]), .REG_DEST_ID(DEST_REG_DECODE_OUT), 
        .REG_DEST_EXE(DEST_REG_EXECUTE_IN), .REG_DEST_MEM(DEST_REG_MEM_IN), 
        .REG_A(INSTRUCTION_DECODE_IN[25:21]), .REG_B(
        INSTRUCTION_DECODE_IN[20:16]), .MUX_A(FORW_SEL_A), .MUX_B(OP_SEL_B_SIG), .MUX_C(FORW_SEL_C), .MUX_D(FORW_SEL_D), .RST_DIV(RST_DIV_SIG), 
        .STALL_BRANCH(STALL_BRANCH), .STALL(STALL) );
  BUF_X2 U2 ( .A(EN_2), .Z(n3) );
  BUF_X1 U3 ( .A(RST), .Z(n6) );
  NOR2_X1 U4 ( .A1(WRONG_FETCH_SIG_1), .A2(n2), .ZN(BPU_SEL_SIG) );
  INV_X1 U5 ( .A(BPU_SEL), .ZN(n2) );
  CLKBUF_X1 U6 ( .A(EN_4), .Z(n1) );
  CLKBUF_X1 U7 ( .A(RST), .Z(n4) );
  CLKBUF_X1 U8 ( .A(RST), .Z(n5) );
endmodule



    module FSM_CU_CW_SIZE29_FETCH_SIGs1_DECODE_SIGs10_EXECUTE_SIGs7_MEM_SIGs8_WB_SIG3_ALU_CODE_SIZE5_IR_SIZE32_OPCODE_SIZE6_FUNC_SIZE11 ( 
        CLK, RST, STALL_BRANCH, STALL, INSTR_HIT_MISS, WRONG_FETCH, OPCODE, 
        FUNC, EN_IF, EN_ID, CONFIRM_JMP, CONFIRM_BRANCH, BRANCH_TYPE, RD1, RD2, 
        SEL_DEST, LHI_SEL, JMP_SEL, EN_EXE, ALU_CODE, OP_SEL, EN_MEM, 
        STORE_MASK, RM, WM, LOAD_TYPE, WB_SEL, WR );
  input [5:0] OPCODE;
  input [10:0] FUNC;
  output [1:0] SEL_DEST;
  output [4:0] ALU_CODE;
  output [1:0] STORE_MASK;
  output [2:0] LOAD_TYPE;
  output [1:0] WB_SEL;
  input CLK, RST, STALL_BRANCH, STALL, INSTR_HIT_MISS, WRONG_FETCH;
  output EN_IF, EN_ID, CONFIRM_JMP, CONFIRM_BRANCH, BRANCH_TYPE, RD1, RD2,
         LHI_SEL, JMP_SEL, EN_EXE, OP_SEL, EN_MEM, RM, WM, WR;
  wire   n265, n266, n267, REG_EN, DIS_DEC, CW1_0, DIS_EXE, \CW3[2] ,
         DISABLE_WR_2, DISABLE_WR_1, n291, n292, n293, n294, n295, n297, n298,
         n299, n300, n301, n1, n2, n3, n4, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264;
  wire   [17:7] CW1;
  wire   [10:8] CW2;
  wire   [6:1] EXE_CW;
  wire   [7:0] MEM_CW;
  wire   [2:0] WB_CW;

  DFFR_X1 \CURRENT_STATE_reg[0]  ( .D(n297), .CK(CLK), .RN(n8), .QN(n301) );
  DFFR_X1 \CURRENT_STATE_reg[2]  ( .D(n295), .CK(CLK), .RN(n8), .Q(n1), .QN(
        n299) );
  DFFR_X1 \CURRENT_STATE_reg[4]  ( .D(n294), .CK(CLK), .RN(n8), .QN(n300) );
  DFFR_X1 \CURRENT_STATE_reg[5]  ( .D(n293), .CK(CLK), .RN(n8), .Q(n2), .QN(
        n263) );
  DFFR_X1 \CURRENT_STATE_reg[3]  ( .D(n292), .CK(CLK), .RN(n8), .QN(n298) );
  DFFR_X1 \CURRENT_STATE_reg[1]  ( .D(n291), .CK(CLK), .RN(n8), .Q(n3), .QN(
        n264) );
  REG_N18 CW_01_REG ( .D({WB_CW, MEM_CW, EXE_CW, MEM_CW[0]}), .Q({CW1, OP_SEL, 
        ALU_CODE, CW1_0}), .EN(REG_EN), .RST(RST), .CLK(CLK) );
  REG_N11 CW_02_REG ( .D(CW1), .Q({CW2, LOAD_TYPE, WM, RM, STORE_MASK, EN_MEM}), .EN(1'b1), .RST(RST), .CLK(CLK) );
  REG_N3 CW_03_REG ( .D(CW2), .Q({\CW3[2] , WB_SEL}), .EN(1'b1), .RST(RST), 
        .CLK(CLK) );
  FD_0 PIPE_DISABLE_WR_1 ( .D(STALL), .CLK(CLK), .EN(1'b1), .RST(RST), .Q(
        DISABLE_WR_1) );
  FD_181 PIPE_DISABLE_WR_2 ( .D(DISABLE_WR_1), .CLK(CLK), .EN(1'b1), .RST(RST), 
        .Q(DISABLE_WR_2) );
  FD_180 FLUSH_DECODE ( .D(WRONG_FETCH), .CLK(CLK), .EN(1'b1), .RST(RST), .Q(
        DIS_DEC) );
  FD_179 FLUSH_EXECUTE ( .D(STALL_BRANCH), .CLK(CLK), .EN(1'b1), .RST(RST), 
        .Q(DIS_EXE) );
  AOI221_X2 U3 ( .B1(n196), .B2(n229), .C1(n243), .C2(n206), .A(n259), .ZN(
        n199) );
  NOR2_X1 U4 ( .A1(MEM_CW[4]), .A2(WB_CW[1]), .ZN(n189) );
  NOR2_X1 U5 ( .A1(n181), .A2(n256), .ZN(n219) );
  BUF_X1 U6 ( .A(n265), .Z(EN_ID) );
  OR2_X1 U7 ( .A1(n3), .A2(n301), .ZN(n220) );
  NAND2_X1 U8 ( .A1(n301), .A2(n3), .ZN(n237) );
  NOR3_X2 U9 ( .A1(n180), .A2(CONFIRM_JMP), .A3(n178), .ZN(n246) );
  NAND4_X1 U10 ( .A1(n257), .A2(n213), .A3(n211), .A4(n258), .ZN(EXE_CW[6]) );
  INV_X1 U11 ( .A(n189), .ZN(n178) );
  AND2_X1 U12 ( .A1(n214), .A2(n199), .ZN(n258) );
  BUF_X1 U13 ( .A(n267), .Z(JMP_SEL) );
  INV_X1 U14 ( .A(n237), .ZN(n181) );
  INV_X1 U15 ( .A(n234), .ZN(n216) );
  BUF_X1 U16 ( .A(n266), .Z(LHI_SEL) );
  INV_X1 U17 ( .A(OPCODE[4]), .ZN(n23) );
  INV_X1 U18 ( .A(RST), .ZN(n8) );
  INV_X1 U19 ( .A(REG_EN), .ZN(n4) );
  OAI21_X1 U20 ( .B1(n301), .B2(n9), .A(n10), .ZN(n297) );
  NAND3_X1 U21 ( .A1(INSTR_HIT_MISS), .A2(n11), .A3(n12), .ZN(n10) );
  NAND4_X1 U22 ( .A1(n13), .A2(n14), .A3(n15), .A4(n16), .ZN(n11) );
  AND3_X1 U23 ( .A1(n17), .A2(n18), .A3(n19), .ZN(n16) );
  MUX2_X1 U24 ( .A(n20), .B(n21), .S(OPCODE[0]), .Z(n15) );
  AOI221_X1 U25 ( .B1(n22), .B2(n23), .C1(n24), .C2(n25), .A(n26), .ZN(n21) );
  AOI221_X1 U26 ( .B1(n27), .B2(n23), .C1(n24), .C2(n28), .A(n29), .ZN(n20) );
  OAI21_X1 U27 ( .B1(n30), .B2(n31), .A(n25), .ZN(n28) );
  OAI221_X1 U28 ( .B1(FUNC[4]), .B2(n32), .C1(n33), .C2(n34), .A(n35), .ZN(n31) );
  AOI21_X1 U29 ( .B1(n36), .B2(n37), .A(n38), .ZN(n35) );
  OAI211_X1 U30 ( .C1(n34), .C2(n39), .A(n40), .B(n41), .ZN(n30) );
  AND3_X1 U31 ( .A1(n42), .A2(n43), .A3(n44), .ZN(n41) );
  NAND2_X1 U32 ( .A1(FUNC[0]), .A2(n45), .ZN(n39) );
  OAI21_X1 U33 ( .B1(n46), .B2(n47), .A(n48), .ZN(n14) );
  MUX2_X1 U34 ( .A(n49), .B(n50), .S(OPCODE[4]), .Z(n47) );
  NOR2_X1 U35 ( .A1(OPCODE[2]), .A2(n51), .ZN(n50) );
  INV_X1 U36 ( .A(n52), .ZN(n13) );
  NAND4_X1 U37 ( .A1(n53), .A2(n54), .A3(n55), .A4(n56), .ZN(n295) );
  NAND4_X1 U38 ( .A1(n57), .A2(n12), .A3(n58), .A4(n34), .ZN(n56) );
  NAND4_X1 U39 ( .A1(n59), .A2(n60), .A3(n61), .A4(n40), .ZN(n58) );
  INV_X1 U40 ( .A(n38), .ZN(n61) );
  OAI21_X1 U41 ( .B1(n62), .B2(n63), .A(n64), .ZN(n55) );
  NAND2_X1 U42 ( .A1(n65), .A2(n1), .ZN(n54) );
  NAND3_X1 U43 ( .A1(n66), .A2(n67), .A3(n68), .ZN(n294) );
  AOI21_X1 U44 ( .B1(n65), .B2(n69), .A(n70), .ZN(n68) );
  NAND4_X1 U45 ( .A1(n71), .A2(n59), .A3(n32), .A4(n72), .ZN(n67) );
  INV_X1 U46 ( .A(n73), .ZN(n59) );
  OAI21_X1 U47 ( .B1(n74), .B2(n75), .A(n64), .ZN(n66) );
  NOR3_X1 U48 ( .A1(n76), .A2(n77), .A3(n78), .ZN(n74) );
  NAND3_X1 U49 ( .A1(n79), .A2(n80), .A3(n81), .ZN(n76) );
  OAI211_X1 U50 ( .C1(n263), .C2(n9), .A(n53), .B(n82), .ZN(n293) );
  AOI22_X1 U51 ( .A1(n83), .A2(n84), .B1(n85), .B2(n64), .ZN(n82) );
  NOR2_X1 U52 ( .A1(n86), .A2(n75), .ZN(n85) );
  NOR3_X1 U53 ( .A1(n87), .A2(OPCODE[4]), .A3(OPCODE[1]), .ZN(n86) );
  AND4_X1 U54 ( .A1(n72), .A2(n40), .A3(n32), .A4(n34), .ZN(n84) );
  NAND2_X1 U55 ( .A1(n88), .A2(FUNC[3]), .ZN(n32) );
  NOR3_X1 U56 ( .A1(n89), .A2(n73), .A3(n90), .ZN(n83) );
  NAND4_X1 U57 ( .A1(n91), .A2(n92), .A3(n42), .A4(n44), .ZN(n73) );
  NAND4_X1 U58 ( .A1(FUNC[4]), .A2(FUNC[3]), .A3(n93), .A4(n94), .ZN(n42) );
  NOR2_X1 U59 ( .A1(FUNC[2]), .A2(n33), .ZN(n93) );
  NAND2_X1 U60 ( .A1(n37), .A2(n45), .ZN(n91) );
  INV_X1 U61 ( .A(n70), .ZN(n53) );
  NAND3_X1 U62 ( .A1(n95), .A2(n96), .A3(n97), .ZN(n292) );
  AOI21_X1 U63 ( .B1(n65), .B2(n98), .A(n70), .ZN(n97) );
  OAI22_X1 U64 ( .A1(INSTR_HIT_MISS), .A2(n99), .B1(n65), .B2(n100), .ZN(n70)
         );
  INV_X1 U65 ( .A(n9), .ZN(n65) );
  OAI221_X1 U66 ( .B1(n101), .B2(n75), .C1(OPCODE[4]), .C2(n102), .A(n64), 
        .ZN(n96) );
  NOR2_X1 U67 ( .A1(n99), .A2(n57), .ZN(n64) );
  NOR3_X1 U68 ( .A1(n103), .A2(n104), .A3(n78), .ZN(n101) );
  OAI21_X1 U69 ( .B1(n105), .B2(n106), .A(n107), .ZN(n103) );
  NAND4_X1 U70 ( .A1(n108), .A2(n71), .A3(n34), .A4(n40), .ZN(n95) );
  NAND2_X1 U71 ( .A1(n37), .A2(n109), .ZN(n34) );
  INV_X1 U72 ( .A(n90), .ZN(n71) );
  NAND3_X1 U73 ( .A1(n57), .A2(n12), .A3(n110), .ZN(n90) );
  AND3_X1 U74 ( .A1(n60), .A2(n111), .A3(n112), .ZN(n110) );
  NAND3_X1 U75 ( .A1(FUNC[3]), .A2(FUNC[0]), .A3(n88), .ZN(n60) );
  INV_X1 U76 ( .A(n99), .ZN(n12) );
  OAI22_X1 U77 ( .A1(n264), .A2(n9), .B1(n99), .B2(n113), .ZN(n291) );
  OAI21_X1 U78 ( .B1(n114), .B2(n115), .A(INSTR_HIT_MISS), .ZN(n113) );
  NOR4_X1 U79 ( .A1(n116), .A2(n117), .A3(n52), .A4(n118), .ZN(n115) );
  MUX2_X1 U80 ( .A(n26), .B(n119), .S(OPCODE[0]), .Z(n118) );
  OAI21_X1 U81 ( .B1(OPCODE[4]), .B2(n120), .A(n17), .ZN(n119) );
  NAND2_X1 U82 ( .A1(n121), .A2(n122), .ZN(n52) );
  OR3_X1 U83 ( .A1(n123), .A2(OPCODE[0]), .A3(n87), .ZN(n121) );
  MUX2_X1 U84 ( .A(n22), .B(n124), .S(n125), .Z(n117) );
  NOR2_X1 U85 ( .A1(n51), .A2(n25), .ZN(n124) );
  OAI211_X1 U86 ( .C1(n23), .C2(n126), .A(n127), .B(n128), .ZN(n116) );
  INV_X1 U87 ( .A(n129), .ZN(n128) );
  NOR4_X1 U88 ( .A1(n130), .A2(n131), .A3(n38), .A4(n132), .ZN(n114) );
  INV_X1 U89 ( .A(n92), .ZN(n132) );
  NAND3_X1 U90 ( .A1(FUNC[3]), .A2(n133), .A3(n37), .ZN(n92) );
  NOR2_X1 U91 ( .A1(n112), .A2(n134), .ZN(n38) );
  NAND2_X1 U92 ( .A1(n88), .A2(n135), .ZN(n112) );
  NOR3_X1 U93 ( .A1(n136), .A2(FUNC[1]), .A3(n137), .ZN(n88) );
  NAND2_X1 U94 ( .A1(n108), .A2(n57), .ZN(n131) );
  AND2_X1 U95 ( .A1(n24), .A2(n138), .ZN(n57) );
  INV_X1 U96 ( .A(n89), .ZN(n108) );
  OAI21_X1 U97 ( .B1(n139), .B2(n33), .A(n43), .ZN(n89) );
  NAND3_X1 U98 ( .A1(FUNC[0]), .A2(n140), .A3(FUNC[1]), .ZN(n43) );
  NAND4_X1 U99 ( .A1(n40), .A2(n44), .A3(n72), .A4(n111), .ZN(n130) );
  NAND2_X1 U100 ( .A1(n37), .A2(n141), .ZN(n111) );
  NOR3_X1 U101 ( .A1(FUNC[2]), .A2(FUNC[4]), .A3(n137), .ZN(n37) );
  INV_X1 U102 ( .A(n94), .ZN(n137) );
  NAND3_X1 U103 ( .A1(n94), .A2(n136), .A3(n36), .ZN(n72) );
  NOR3_X1 U104 ( .A1(n45), .A2(n134), .A3(n109), .ZN(n36) );
  INV_X1 U105 ( .A(FUNC[3]), .ZN(n109) );
  INV_X1 U106 ( .A(FUNC[1]), .ZN(n45) );
  INV_X1 U107 ( .A(FUNC[2]), .ZN(n136) );
  NAND2_X1 U108 ( .A1(n141), .A2(n140), .ZN(n44) );
  INV_X1 U109 ( .A(n139), .ZN(n140) );
  NAND4_X1 U110 ( .A1(FUNC[2]), .A2(n135), .A3(n142), .A4(n143), .ZN(n139) );
  NOR4_X1 U111 ( .A1(FUNC[9]), .A2(FUNC[8]), .A3(FUNC[7]), .A4(FUNC[6]), .ZN(
        n143) );
  NOR2_X1 U112 ( .A1(FUNC[5]), .A2(FUNC[10]), .ZN(n142) );
  NOR2_X1 U113 ( .A1(FUNC[0]), .A2(FUNC[1]), .ZN(n141) );
  NAND4_X1 U114 ( .A1(n94), .A2(n133), .A3(FUNC[2]), .A4(n135), .ZN(n40) );
  NOR2_X1 U115 ( .A1(FUNC[3]), .A2(FUNC[4]), .ZN(n135) );
  INV_X1 U116 ( .A(n33), .ZN(n133) );
  NAND2_X1 U117 ( .A1(FUNC[1]), .A2(n134), .ZN(n33) );
  INV_X1 U118 ( .A(FUNC[0]), .ZN(n134) );
  NOR4_X1 U119 ( .A1(FUNC[10]), .A2(FUNC[6]), .A3(n144), .A4(n145), .ZN(n94)
         );
  OR3_X1 U120 ( .A1(FUNC[7]), .A2(FUNC[9]), .A3(FUNC[8]), .ZN(n145) );
  INV_X1 U121 ( .A(FUNC[5]), .ZN(n144) );
  NAND2_X1 U122 ( .A1(n146), .A2(n9), .ZN(n99) );
  OAI22_X1 U123 ( .A1(STALL_BRANCH), .A2(n146), .B1(n147), .B2(n4), .ZN(n9) );
  NOR4_X1 U124 ( .A1(n148), .A2(n149), .A3(n104), .A4(n63), .ZN(n147) );
  NAND3_X1 U125 ( .A1(n107), .A2(n81), .A3(n150), .ZN(n63) );
  INV_X1 U126 ( .A(n151), .ZN(n150) );
  OAI21_X1 U127 ( .B1(n102), .B2(OPCODE[4]), .A(n79), .ZN(n151) );
  AOI22_X1 U128 ( .A1(n152), .A2(n24), .B1(n153), .B2(n22), .ZN(n79) );
  OR2_X1 U129 ( .A1(n125), .A2(n23), .ZN(n153) );
  AOI221_X1 U130 ( .B1(n152), .B2(n27), .C1(n154), .C2(n48), .A(n49), .ZN(n102) );
  AOI21_X1 U131 ( .B1(n49), .B2(n123), .A(n29), .ZN(n81) );
  INV_X1 U132 ( .A(n127), .ZN(n29) );
  NAND2_X1 U133 ( .A1(n155), .A2(OPCODE[2]), .ZN(n127) );
  AOI21_X1 U134 ( .B1(OPCODE[0]), .B2(n156), .A(n26), .ZN(n107) );
  AND3_X1 U135 ( .A1(n157), .A2(n23), .A3(n158), .ZN(n26) );
  OR2_X1 U136 ( .A1(n156), .A2(n155), .ZN(n104) );
  NOR3_X1 U137 ( .A1(n25), .A2(n51), .A3(n23), .ZN(n155) );
  INV_X1 U138 ( .A(n17), .ZN(n156) );
  NAND2_X1 U139 ( .A1(n159), .A2(n25), .ZN(n17) );
  OAI21_X1 U140 ( .B1(n160), .B2(n105), .A(n161), .ZN(n149) );
  INV_X1 U141 ( .A(n77), .ZN(n161) );
  NAND2_X1 U142 ( .A1(n122), .A2(n162), .ZN(n77) );
  NAND3_X1 U143 ( .A1(n46), .A2(n23), .A3(OPCODE[0]), .ZN(n162) );
  NAND3_X1 U144 ( .A1(n46), .A2(n23), .A3(n138), .ZN(n122) );
  OR4_X1 U145 ( .A1(n163), .A2(n78), .A3(n75), .A4(n129), .ZN(n148) );
  OAI211_X1 U146 ( .C1(OPCODE[1]), .C2(n106), .A(n164), .B(n80), .ZN(n129) );
  NAND3_X1 U147 ( .A1(n154), .A2(n152), .A3(n123), .ZN(n80) );
  NOR2_X1 U148 ( .A1(n25), .A2(OPCODE[4]), .ZN(n123) );
  OAI21_X1 U149 ( .B1(n24), .B2(n159), .A(n48), .ZN(n164) );
  NOR4_X1 U150 ( .A1(n165), .A2(OPCODE[2]), .A3(OPCODE[3]), .A4(OPCODE[4]), 
        .ZN(n159) );
  INV_X1 U151 ( .A(n24), .ZN(n106) );
  NOR3_X1 U152 ( .A1(OPCODE[2]), .A2(OPCODE[4]), .A3(n51), .ZN(n24) );
  NAND3_X1 U153 ( .A1(n166), .A2(n120), .A3(n167), .ZN(n75) );
  AOI22_X1 U154 ( .A1(n168), .A2(n125), .B1(n138), .B2(n49), .ZN(n167) );
  NOR2_X1 U155 ( .A1(OPCODE[1]), .A2(OPCODE[0]), .ZN(n138) );
  INV_X1 U156 ( .A(n62), .ZN(n166) );
  AOI21_X1 U157 ( .B1(n126), .B2(n169), .A(n23), .ZN(n62) );
  OAI21_X1 U158 ( .B1(n168), .B2(n27), .A(n152), .ZN(n169) );
  INV_X1 U159 ( .A(n120), .ZN(n27) );
  NAND2_X1 U160 ( .A1(n154), .A2(n25), .ZN(n120) );
  INV_X1 U161 ( .A(n160), .ZN(n154) );
  NAND3_X1 U162 ( .A1(OPCODE[3]), .A2(n165), .A3(OPCODE[2]), .ZN(n160) );
  INV_X1 U163 ( .A(n19), .ZN(n168) );
  NAND2_X1 U164 ( .A1(n158), .A2(OPCODE[3]), .ZN(n19) );
  NOR3_X1 U165 ( .A1(n170), .A2(OPCODE[1]), .A3(n165), .ZN(n158) );
  OAI21_X1 U166 ( .B1(n49), .B2(n46), .A(n48), .ZN(n126) );
  INV_X1 U167 ( .A(n105), .ZN(n48) );
  NAND2_X1 U168 ( .A1(OPCODE[0]), .A2(OPCODE[1]), .ZN(n105) );
  NAND2_X1 U169 ( .A1(n18), .A2(n171), .ZN(n78) );
  OR3_X1 U170 ( .A1(n172), .A2(OPCODE[0]), .A3(n23), .ZN(n171) );
  AOI211_X1 U171 ( .C1(n46), .C2(OPCODE[1]), .A(n22), .B(n49), .ZN(n172) );
  NOR3_X1 U172 ( .A1(n51), .A2(OPCODE[1]), .A3(n170), .ZN(n22) );
  NAND2_X1 U173 ( .A1(n157), .A2(n165), .ZN(n51) );
  NOR3_X1 U174 ( .A1(n157), .A2(OPCODE[2]), .A3(n165), .ZN(n46) );
  INV_X1 U175 ( .A(OPCODE[3]), .ZN(n157) );
  NAND3_X1 U176 ( .A1(n125), .A2(n25), .A3(n49), .ZN(n18) );
  INV_X1 U177 ( .A(n87), .ZN(n49) );
  NAND3_X1 U178 ( .A1(n170), .A2(n165), .A3(OPCODE[3]), .ZN(n87) );
  INV_X1 U179 ( .A(OPCODE[5]), .ZN(n165) );
  INV_X1 U180 ( .A(OPCODE[2]), .ZN(n170) );
  INV_X1 U181 ( .A(OPCODE[1]), .ZN(n25) );
  NOR2_X1 U182 ( .A1(n152), .A2(n23), .ZN(n125) );
  INV_X1 U183 ( .A(OPCODE[0]), .ZN(n152) );
  AND2_X1 U184 ( .A1(n100), .A2(n173), .ZN(n146) );
  NAND3_X1 U185 ( .A1(n174), .A2(n175), .A3(n176), .ZN(n173) );
  NOR2_X1 U186 ( .A1(DISABLE_WR_2), .A2(n177), .ZN(WR) );
  INV_X1 U187 ( .A(\CW3[2] ), .ZN(n177) );
  OR2_X1 U188 ( .A1(EXE_CW[6]), .A2(SEL_DEST[0]), .ZN(WB_CW[2]) );
  OR4_X1 U189 ( .A1(n178), .A2(n179), .A3(n180), .A4(n181), .ZN(SEL_DEST[1])
         );
  NAND2_X1 U190 ( .A1(n182), .A2(n183), .ZN(SEL_DEST[0]) );
  INV_X1 U191 ( .A(WB_CW[0]), .ZN(n183) );
  OAI21_X1 U192 ( .B1(n184), .B2(n185), .A(n186), .ZN(WB_CW[0]) );
  NAND2_X1 U193 ( .A1(n187), .A2(n188), .ZN(RD2) );
  NAND3_X1 U194 ( .A1(n189), .A2(n190), .A3(n191), .ZN(RD1) );
  OAI21_X1 U195 ( .B1(n192), .B2(n185), .A(n193), .ZN(MEM_CW[6]) );
  OAI21_X1 U196 ( .B1(n194), .B2(n195), .A(n196), .ZN(n193) );
  INV_X1 U197 ( .A(n197), .ZN(MEM_CW[5]) );
  INV_X1 U198 ( .A(n186), .ZN(MEM_CW[3]) );
  NOR2_X1 U199 ( .A1(n192), .A2(n198), .ZN(MEM_CW[1]) );
  NAND3_X1 U200 ( .A1(n199), .A2(n200), .A3(n201), .ZN(EXE_CW[5]) );
  NAND3_X1 U201 ( .A1(n202), .A2(n201), .A3(n203), .ZN(EXE_CW[4]) );
  AOI221_X1 U202 ( .B1(n204), .B2(n205), .C1(n206), .C2(n174), .A(n207), .ZN(
        n203) );
  OAI21_X1 U203 ( .B1(n184), .B2(n208), .A(n209), .ZN(n207) );
  INV_X1 U204 ( .A(n210), .ZN(n184) );
  INV_X1 U205 ( .A(n211), .ZN(n204) );
  INV_X1 U206 ( .A(n212), .ZN(n202) );
  OAI21_X1 U207 ( .B1(n213), .B2(n298), .A(n214), .ZN(n212) );
  NAND3_X1 U208 ( .A1(n201), .A2(n214), .A3(n215), .ZN(EXE_CW[3]) );
  AOI221_X1 U209 ( .B1(n206), .B2(n216), .C1(n217), .C2(n210), .A(n218), .ZN(
        n215) );
  AOI21_X1 U210 ( .B1(n213), .B2(n209), .A(n219), .ZN(n218) );
  OAI211_X1 U211 ( .C1(n220), .C2(n221), .A(n222), .B(n223), .ZN(EXE_CW[2]) );
  AOI221_X1 U212 ( .B1(n224), .B2(n210), .C1(n196), .C2(n225), .A(n226), .ZN(
        n223) );
  NAND2_X1 U213 ( .A1(n220), .A2(n175), .ZN(n210) );
  OAI211_X1 U214 ( .C1(n175), .C2(n198), .A(n222), .B(n227), .ZN(EXE_CW[1]) );
  AOI221_X1 U215 ( .B1(n228), .B2(n224), .C1(n229), .C2(n230), .A(n231), .ZN(
        n227) );
  AOI21_X1 U216 ( .B1(n232), .B2(n233), .A(n192), .ZN(n231) );
  OAI21_X1 U217 ( .B1(n234), .B2(n235), .A(n213), .ZN(n224) );
  INV_X1 U218 ( .A(n236), .ZN(n222) );
  OAI211_X1 U219 ( .C1(n221), .C2(n237), .A(n201), .B(n238), .ZN(n236) );
  AOI21_X1 U220 ( .B1(n228), .B2(n225), .A(n239), .ZN(n238) );
  NAND2_X1 U221 ( .A1(n240), .A2(n209), .ZN(n225) );
  INV_X1 U222 ( .A(n217), .ZN(n240) );
  OAI211_X1 U223 ( .C1(n241), .C2(n235), .A(n211), .B(n208), .ZN(n217) );
  NOR3_X1 U224 ( .A1(n180), .A2(CONFIRM_JMP), .A3(n179), .ZN(n201) );
  OAI221_X1 U225 ( .B1(n241), .B2(n242), .C1(n192), .C2(n221), .A(n100), .ZN(
        n179) );
  NAND3_X1 U226 ( .A1(n196), .A2(n243), .A3(n244), .ZN(n100) );
  NOR3_X1 U227 ( .A1(n4), .A2(n245), .A3(n163), .ZN(EN_IF) );
  INV_X1 U228 ( .A(INSTR_HIT_MISS), .ZN(n163) );
  AOI21_X1 U229 ( .B1(n196), .B2(n174), .A(MEM_CW[0]), .ZN(n245) );
  INV_X1 U230 ( .A(n246), .ZN(MEM_CW[0]) );
  NOR3_X1 U231 ( .A1(n4), .A2(DIS_DEC), .A3(n246), .ZN(n265) );
  NAND3_X1 U232 ( .A1(n187), .A2(n186), .A3(n182), .ZN(WB_CW[1]) );
  AND4_X1 U233 ( .A1(n200), .A2(n247), .A3(n232), .A4(n248), .ZN(n182) );
  AOI211_X1 U234 ( .C1(n229), .C2(n228), .A(n249), .B(LHI_SEL), .ZN(n248) );
  NOR2_X1 U235 ( .A1(n237), .A2(n250), .ZN(n266) );
  AND2_X1 U236 ( .A1(n209), .A2(n251), .ZN(n232) );
  OAI21_X1 U237 ( .B1(n216), .B2(n174), .A(n252), .ZN(n251) );
  NAND2_X1 U238 ( .A1(n253), .A2(n243), .ZN(n209) );
  NAND2_X1 U239 ( .A1(n206), .A2(n254), .ZN(n247) );
  AOI22_X1 U240 ( .A1(n196), .A2(n255), .B1(n205), .B2(n249), .ZN(n200) );
  INV_X1 U241 ( .A(n208), .ZN(n249) );
  NAND2_X1 U242 ( .A1(n253), .A2(n254), .ZN(n208) );
  AOI21_X1 U243 ( .B1(n196), .B2(n195), .A(MEM_CW[7]), .ZN(n186) );
  OAI221_X1 U244 ( .B1(n250), .B2(n220), .C1(n192), .C2(n185), .A(n197), .ZN(
        MEM_CW[7]) );
  NAND2_X1 U245 ( .A1(n194), .A2(n230), .ZN(n197) );
  NAND2_X1 U246 ( .A1(n175), .A2(n192), .ZN(n230) );
  INV_X1 U247 ( .A(n250), .ZN(n194) );
  INV_X1 U248 ( .A(n256), .ZN(n192) );
  NAND2_X1 U249 ( .A1(n254), .A2(n176), .ZN(n250) );
  INV_X1 U250 ( .A(n221), .ZN(n195) );
  INV_X1 U251 ( .A(EXE_CW[6]), .ZN(n187) );
  AOI21_X1 U252 ( .B1(n237), .B2(n220), .A(n221), .ZN(n259) );
  NAND2_X1 U253 ( .A1(n216), .A2(n176), .ZN(n221) );
  NOR2_X1 U254 ( .A1(n235), .A2(n219), .ZN(n206) );
  AND2_X1 U255 ( .A1(n252), .A2(n254), .ZN(n229) );
  NOR2_X1 U256 ( .A1(n98), .A2(n299), .ZN(n254) );
  INV_X1 U257 ( .A(n235), .ZN(n252) );
  NOR2_X1 U258 ( .A1(n226), .A2(n239), .ZN(n214) );
  NOR3_X1 U259 ( .A1(n220), .A2(n260), .A3(n235), .ZN(n239) );
  NOR3_X1 U260 ( .A1(n175), .A2(n260), .A3(n235), .ZN(n226) );
  NAND2_X1 U261 ( .A1(n263), .A2(n69), .ZN(n235) );
  NAND2_X1 U262 ( .A1(n216), .A2(n244), .ZN(n211) );
  NAND2_X1 U263 ( .A1(n244), .A2(n1), .ZN(n213) );
  OAI21_X1 U264 ( .B1(n228), .B2(n205), .A(n244), .ZN(n257) );
  INV_X1 U265 ( .A(n233), .ZN(n244) );
  NAND2_X1 U266 ( .A1(n263), .A2(n300), .ZN(n233) );
  INV_X1 U267 ( .A(n219), .ZN(n205) );
  INV_X1 U268 ( .A(n188), .ZN(MEM_CW[4]) );
  AOI21_X1 U269 ( .B1(n228), .B2(n255), .A(MEM_CW[2]), .ZN(n188) );
  NOR2_X1 U270 ( .A1(n198), .A2(n219), .ZN(MEM_CW[2]) );
  INV_X1 U271 ( .A(n198), .ZN(n255) );
  NAND2_X1 U272 ( .A1(n253), .A2(n216), .ZN(n198) );
  NAND2_X1 U273 ( .A1(n299), .A2(n98), .ZN(n234) );
  INV_X1 U274 ( .A(n220), .ZN(n228) );
  NOR2_X1 U275 ( .A1(STALL_BRANCH), .A2(STALL), .ZN(REG_EN) );
  NOR2_X1 U276 ( .A1(DIS_EXE), .A2(n261), .ZN(EN_EXE) );
  INV_X1 U277 ( .A(CW1_0), .ZN(n261) );
  OAI21_X1 U278 ( .B1(n175), .B2(n185), .A(n191), .ZN(CONFIRM_JMP) );
  AOI21_X1 U279 ( .B1(n256), .B2(n180), .A(JMP_SEL), .ZN(n191) );
  AOI21_X1 U280 ( .B1(n220), .B2(n237), .A(n185), .ZN(n267) );
  NOR2_X1 U281 ( .A1(n264), .A2(n301), .ZN(n256) );
  NAND2_X1 U282 ( .A1(n243), .A2(n176), .ZN(n185) );
  INV_X1 U283 ( .A(n242), .ZN(n176) );
  NAND2_X1 U284 ( .A1(n69), .A2(n2), .ZN(n242) );
  INV_X1 U285 ( .A(n260), .ZN(n243) );
  NAND2_X1 U286 ( .A1(n299), .A2(n298), .ZN(n260) );
  INV_X1 U287 ( .A(n190), .ZN(CONFIRM_BRANCH) );
  AOI21_X1 U288 ( .B1(n196), .B2(n180), .A(BRANCH_TYPE), .ZN(n190) );
  INV_X1 U289 ( .A(n262), .ZN(n180) );
  INV_X1 U290 ( .A(n175), .ZN(n196) );
  NAND2_X1 U291 ( .A1(n264), .A2(n301), .ZN(n175) );
  NOR2_X1 U292 ( .A1(n262), .A2(n220), .ZN(BRANCH_TYPE) );
  NAND2_X1 U293 ( .A1(n253), .A2(n174), .ZN(n262) );
  INV_X1 U294 ( .A(n241), .ZN(n174) );
  NAND2_X1 U295 ( .A1(n1), .A2(n98), .ZN(n241) );
  INV_X1 U296 ( .A(n298), .ZN(n98) );
  NOR2_X1 U297 ( .A1(n69), .A2(n263), .ZN(n253) );
  INV_X1 U298 ( .A(n300), .ZN(n69) );
endmodule


module DLX ( CLK, RST, DATA_IN_INSTR, DATA_IN_MEM, RM, WM, ADDR_MEM, 
        DATA_OUT_MEM, ADDR_INSTR );
  input [7:0] DATA_IN_INSTR;
  input [31:0] DATA_IN_MEM;
  output [31:0] ADDR_MEM;
  output [31:0] DATA_OUT_MEM;
  output [31:0] ADDR_INSTR;
  input CLK, RST;
  output RM, WM;
  wire   STALL_BRANCH, STALL, INSTR_CACHE_H_M, WRONG_FETCH, INSTR_SIG_31,
         INSTR_SIG_30, INSTR_SIG_29, INSTR_SIG_28, INSTR_SIG_27, INSTR_SIG_26,
         EN_IF_SIG, EN_2_SIG, CONFIRM_JMP_SIG, CONFIRM_BRANCH_SIG,
         BRANCH_TYPE_SIG, RD1_SIG, RD2_SIG, LHI_SEL_SIG, JMP_SEL_SIG, EN_3_SIG,
         OP_SEL_SIG, EN_4_SIG, WR_SIG;
  wire   [10:0] INSTR_SIG;
  wire   [1:0] SEL_DEST_SIG;
  wire   [4:0] ALU_CODE_SIG;
  wire   [1:0] STORE_MASK;
  wire   [2:0] LOAD_TYPE;
  wire   [1:0] SEL_SIG;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14;

  FSM_CU_CW_SIZE29_FETCH_SIGs1_DECODE_SIGs10_EXECUTE_SIGs7_MEM_SIGs8_WB_SIG3_ALU_CODE_SIZE5_IR_SIZE32_OPCODE_SIZE6_FUNC_SIZE11 INST_CU ( 
        .CLK(CLK), .RST(RST), .STALL_BRANCH(STALL_BRANCH), .STALL(STALL), 
        .INSTR_HIT_MISS(INSTR_CACHE_H_M), .WRONG_FETCH(WRONG_FETCH), .OPCODE({
        INSTR_SIG_31, INSTR_SIG_30, INSTR_SIG_29, INSTR_SIG_28, INSTR_SIG_27, 
        INSTR_SIG_26}), .FUNC(INSTR_SIG), .EN_IF(EN_IF_SIG), .EN_ID(EN_2_SIG), 
        .CONFIRM_JMP(CONFIRM_JMP_SIG), .CONFIRM_BRANCH(CONFIRM_BRANCH_SIG), 
        .BRANCH_TYPE(BRANCH_TYPE_SIG), .RD1(RD1_SIG), .RD2(RD2_SIG), 
        .SEL_DEST(SEL_DEST_SIG), .LHI_SEL(LHI_SEL_SIG), .JMP_SEL(JMP_SEL_SIG), 
        .EN_EXE(EN_3_SIG), .ALU_CODE(ALU_CODE_SIG), .OP_SEL(OP_SEL_SIG), 
        .EN_MEM(EN_4_SIG), .STORE_MASK(STORE_MASK), .RM(RM), .WM(WM), 
        .LOAD_TYPE(LOAD_TYPE), .WB_SEL(SEL_SIG), .WR(WR_SIG) );
  DATAPATH_N32_N_ADDR5_IMM_SIZE16_OP_CODE_SIZE6_M5_ALUSIZE5 DATAPATH_INST ( 
        .CLK(CLK), .RST(RST), .EN_PC(EN_IF_SIG), .EN_1(EN_IF_SIG), .EN_2(
        EN_2_SIG), .CONFIRM_JMP(CONFIRM_JMP_SIG), .CONFIRM_BRANCH(
        CONFIRM_BRANCH_SIG), .BRANCH_TYPE(BRANCH_TYPE_SIG), .RD1(RD1_SIG), 
        .RD2(RD2_SIG), .WR(WR_SIG), .SEL_DEST(SEL_DEST_SIG), .LHI_SEL(
        LHI_SEL_SIG), .JMP_SEL(JMP_SEL_SIG), .EN_3(EN_3_SIG), .ALU_CODE(
        ALU_CODE_SIG), .OP_SEL(OP_SEL_SIG), .EN_4(EN_4_SIG), .STORE_MASK(
        STORE_MASK), .LOAD_TYPE(LOAD_TYPE), .SEL(SEL_SIG), .DATA_IN_IRAM(
        DATA_IN_INSTR), .DATA_IN_MEM(DATA_IN_MEM), .DATA_OUT_MEM(DATA_OUT_MEM), 
        .ADDR_MEM(ADDR_MEM), .INSTR_CACHE_H_M(INSTR_CACHE_H_M), .ADDR_IRAM(
        ADDR_INSTR), .INSTR({INSTR_SIG_31, INSTR_SIG_30, INSTR_SIG_29, 
        INSTR_SIG_28, INSTR_SIG_27, INSTR_SIG_26, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, INSTR_SIG}), 
        .STALL(STALL), .STALL_BRANCH(STALL_BRANCH), .WRONG_FETCH(WRONG_FETCH)
         );
endmodule

