library IEEE;
use IEEE.std_logic_1164.all;
use work.myTypes.all;

entity EXECUTE is
	generic (	N:		integer;
			N_ADDR:		integer;
			ALUSIZE:	integer);
	port	(	REG_A:		in	std_logic_vector(N-1 downto 0);
			REG_B:		in	std_logic_vector(N-1 downto 0);
			IMMEDIATE:	in	std_logic_vector(N-1 downto 0);
			FORW_ALU_MEM:	in	std_logic_vector(N-1 downto 0);
			FORW_ALU_WB:	in	std_logic_vector(N-1 downto 0);
			FORW_MEM_WB:	in	std_logic_vector(N-1 downto 0);
			DEST_REG_IN:	in	std_logic_vector(N_ADDR-1 downto 0);
			ALU_CODE:	in 	std_logic_vector(ALUSIZE-1 downto 0);
			OP_SEL_A:	in	std_logic_vector(1 downto 0);
			OP_SEL_B:	in	std_logic_vector(2 downto 0);
			CLK:		in	std_logic;
			RST:		in	std_logic;
			DEST_REG_OUT:	out	std_logic_vector(N_ADDR-1 downto 0);
			OUTPUT_ALU:	out	std_logic_vector(N-1 downto 0);
			RST_DIV: 	in 	std_logic;
			REG_B_OUT:	out	std_logic_vector(N-1 downto 0));
end EXECUTE;

architecture STRUCTURAL of EXECUTE is

-- Component Declaration

	component MUX41_GEN
		generic (	N:	integer);
		port (		A:	in	std_logic_vector(N-1 downto 0);
				B:	in	std_logic_vector(N-1 downto 0);
				C:	in	std_logic_vector(N-1 downto 0);
				D:	in	std_logic_vector(N-1 downto 0);
				SEL:	in	std_logic_vector(1 downto 0);
				Y:	out	std_logic_vector(N-1 downto 0));
	end component;
	
	component MUX51_GEN
		generic (	N:	integer);
		port (		A:	in	std_logic_vector(N-1 downto 0);
				B:	in	std_logic_vector(N-1 downto 0);
				C:	in	std_logic_vector(N-1 downto 0);
				D:	in	std_logic_vector(N-1 downto 0);
				E:	in	std_logic_vector(N-1 downto 0);
				SEL:	in	std_logic_vector(2 downto 0);
				Y:	out	std_logic_vector(N-1 downto 0));
	end component;

	component ALU
		generic (	N:		integer;
				ALU_SIZE:	integer);
		port	(	IN_A:		in	std_logic_vector(N-1 downto 0);
				IN_B:		in	std_logic_vector(N-1 downto 0);
				ALU_OP_CODE:	in 	std_logic_vector(ALU_SIZE-1 downto 0);
				CLK:		in	std_logic;
				RST:		in	std_logic;
				RST_DIV:	in 	std_logic;
				OUT_ALU:	out	std_logic_vector(N-1 downto 0));
	end component;


-- Signal declaration

	signal IN_A_MUX_A_SIG:	std_logic_vector(N-1 downto 0);
	signal IN_B_MUX_A_SIG:	std_logic_vector(N-1 downto 0);
	signal IN_C_MUX_A_SIG:	std_logic_vector(N-1 downto 0);
	signal IN_D_MUX_A_SIG:	std_logic_vector(N-1 downto 0);
	signal IN_A_MUX_B_SIG:	std_logic_vector(N-1 downto 0);
	signal IN_B_MUX_B_SIG:	std_logic_vector(N-1 downto 0);
	signal IN_C_MUX_B_SIG:	std_logic_vector(N-1 downto 0);
	signal IN_D_MUX_B_SIG:	std_logic_vector(N-1 downto 0);
	signal IN_E_MUX_B_SIG:	std_logic_vector(N-1 downto 0);
	signal DEST_REG_SIG:	std_logic_vector(N_ADDR-1 downto 0);
	signal IN_A_ALU_SIG:	std_logic_vector(N-1 downto 0);
	signal IN_B_ALU_SIG:	std_logic_vector(N-1 downto 0);
	signal RST_DIV_SIG: 	std_logic;

	begin

		-- Signal mapping
	
		IN_A_MUX_A_SIG <= REG_A;
		IN_B_MUX_A_SIG <= FORW_ALU_MEM;
		IN_C_MUX_A_SIG <= FORW_ALU_WB;
		IN_D_MUX_A_SIG <= FORW_MEM_WB;
		IN_A_MUX_B_SIG <= REG_B;
		IN_B_MUX_B_SIG <= FORW_ALU_MEM;
		IN_C_MUX_B_SIG <= FORW_ALU_WB;
		IN_D_MUX_B_SIG <= FORW_MEM_WB;
		IN_E_MUX_B_SIG <= IMMEDIATE;
		DEST_REG_SIG <= DEST_REG_IN;	-- Dest Reg buffer
		DEST_REG_OUT <= DEST_REG_SIG;	-- Dest Reg buffer
		REG_B_OUT <= REG_B; 		-- FOR STORE INS
		RST_DIV_SIG <= RST_DIV;

		-- Port Mapping
		
		OP_A_SEL_MUX: MUX41_GEN	generic map(	N => N)
					port map(	A => IN_A_MUX_A_SIG,
							B => IN_B_MUX_A_SIG,
							C => IN_C_MUX_A_SIG,
							D => IN_D_MUX_A_SIG,
							SEL => OP_SEL_A,
							Y => IN_A_ALU_SIG);

		OP_B_SEL_MUX: MUX51_GEN	generic map(	N => N)
					port map(	A => IN_A_MUX_B_SIG,
							B => IN_B_MUX_B_SIG,
							C => IN_C_MUX_B_SIG,
							D => IN_D_MUX_B_SIG,
							E => IN_E_MUX_B_SIG,
							SEL => OP_SEL_B,
							Y => IN_B_ALU_SIG);
		
		ALUCOMP: ALU	generic map(	N => N,
						ALU_SIZE => ALUSIZE)
				port map(	IN_A => IN_A_ALU_SIG,
						IN_B => IN_B_ALU_SIG,
						ALU_OP_CODE => ALU_CODE,
						CLK => CLK,
						RST => RST,
						RST_DIV => RST_DIV_SIG,
						OUT_ALU => OUTPUT_ALU);

end STRUCTURAL;

configuration CFG_EXECUTE_STRUCTURAL of EXECUTE is
	for STRUCTURAL
		for all: MUX41_GEN
			use configuration WORK.CFG_MUX41_GEN_BEHAVIORAL;
		end for;
		for all: MUX51_GEN
			use configuration WORK.CFG_MUX51_GEN_BEHAVIORAL;
		end for;
		for all: ALU
			 use configuration WORK.CFG_ALU_STRUCTURAL;
		end for;
	end for;
end CFG_EXECUTE_STRUCTURAL;
