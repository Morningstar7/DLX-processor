library IEEE;
use IEEE.std_logic_1164.all;

entity MUX41 is
	port (		A:	in	std_logic;
			B:	in	std_logic;
			C:	in	std_logic;
			D:	in	std_logic;
			SEL:	in	std_logic_vector(1 downto 0);
			Y:	out	std_logic);
end MUX41;

architecture BEHAVIORAL of MUX41 is

	begin

		Y <=	A when SEL = "11" else
			B when SEL = "10" else
			C when SEL = "01" else
			D;

end BEHAVIORAL;

configuration CFG_MUX41_BEHAVIORAL of MUX41 is
	for BEHAVIORAL
	end for;
end CFG_MUX41_BEHAVIORAL;